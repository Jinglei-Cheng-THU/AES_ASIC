
module TOP_PAD ( CLK, RSTB, START, WR, DIN, ADDR, OK, DOUT );
  input [7:0] DIN;
  input [6:0] ADDR;
  output [7:0] DOUT;
  input CLK, RSTB, START, WR;
  output OK;
  wire   n_CLK, n_RSTB, n_WR, n_START, n_OK, top_core_clk_slow,
         top_core_k_ready, top_core_op, top_core_t_ready, top_core_c_ready,
         top_core_Core_Full, top_core_io_n1343, top_core_io_n1342,
         top_core_io_n1341, top_core_io_n1340, top_core_io_n1339,
         top_core_io_n1338, top_core_io_n1337, top_core_io_n1336,
         top_core_io_n1335, top_core_io_n1334, top_core_io_n1333,
         top_core_io_n1332, top_core_io_n1331, top_core_io_n1330,
         top_core_io_n1329, top_core_io_n1328, top_core_io_n1327,
         top_core_io_n1326, top_core_io_n1325, top_core_io_n1324,
         top_core_io_n1323, top_core_io_n1322, top_core_io_n1321,
         top_core_io_n1320, top_core_io_n1319, top_core_io_n1318,
         top_core_io_n1317, top_core_io_n1316, top_core_io_n1315,
         top_core_io_n1314, top_core_io_n1313, top_core_io_n1312,
         top_core_io_n1311, top_core_io_n1310, top_core_io_n1309,
         top_core_io_n1308, top_core_io_n1307, top_core_io_n1306,
         top_core_io_n1305, top_core_io_n1304, top_core_io_n1303,
         top_core_io_n1302, top_core_io_n1301, top_core_io_n1300,
         top_core_io_n1299, top_core_io_n1298, top_core_io_n1297,
         top_core_io_n1296, top_core_io_n1295, top_core_io_n1294,
         top_core_io_n1293, top_core_io_n1292, top_core_io_n1291,
         top_core_io_n1290, top_core_io_n1289, top_core_io_n1288,
         top_core_io_n1287, top_core_io_n1286, top_core_io_n1285,
         top_core_io_n1284, top_core_io_n1283, top_core_io_n1282,
         top_core_io_n1281, top_core_io_n1280, top_core_io_n1279,
         top_core_io_n1278, top_core_io_n1277, top_core_io_n1276,
         top_core_io_n1275, top_core_io_n1274, top_core_io_n1273,
         top_core_io_n1272, top_core_io_n1271, top_core_io_n1270,
         top_core_io_n1269, top_core_io_n1268, top_core_io_n1267,
         top_core_io_n1266, top_core_io_n1265, top_core_io_n1264,
         top_core_io_n1263, top_core_io_n1262, top_core_io_n1261,
         top_core_io_n1260, top_core_io_n1259, top_core_io_n1258,
         top_core_io_n1257, top_core_io_n1256, top_core_io_n1255,
         top_core_io_n1254, top_core_io_n1253, top_core_io_n1252,
         top_core_io_n1251, top_core_io_n1250, top_core_io_n1249,
         top_core_io_n1248, top_core_io_n1247, top_core_io_n1246,
         top_core_io_n1245, top_core_io_n1244, top_core_io_n1243,
         top_core_io_n1242, top_core_io_n1241, top_core_io_n1240,
         top_core_io_n1239, top_core_io_n1238, top_core_io_n1237,
         top_core_io_n1236, top_core_io_n1235, top_core_io_n1234,
         top_core_io_n1233, top_core_io_n1232, top_core_io_n1231,
         top_core_io_n1230, top_core_io_n1229, top_core_io_n1228,
         top_core_io_n1227, top_core_io_n1226, top_core_io_n1225,
         top_core_io_n1224, top_core_io_n1223, top_core_io_n1222,
         top_core_io_n1221, top_core_io_n1220, top_core_io_n1219,
         top_core_io_n1218, top_core_io_n1217, top_core_io_n1216,
         top_core_io_n1215, top_core_io_n1214, top_core_io_n1213,
         top_core_io_n1212, top_core_io_n1211, top_core_io_n1210,
         top_core_io_n1209, top_core_io_n1208, top_core_io_n1207,
         top_core_io_n1206, top_core_io_n1205, top_core_io_n1204,
         top_core_io_n1203, top_core_io_n1202, top_core_io_n1201,
         top_core_io_n1200, top_core_io_n1199, top_core_io_n1198,
         top_core_io_n1197, top_core_io_n1196, top_core_io_n1195,
         top_core_io_n1194, top_core_io_n1193, top_core_io_n1192,
         top_core_io_n1191, top_core_io_n1190, top_core_io_n1189,
         top_core_io_n1188, top_core_io_n1187, top_core_io_n1186,
         top_core_io_n1185, top_core_io_n1184, top_core_io_n1183,
         top_core_io_n1182, top_core_io_n1180, top_core_io_n1179,
         top_core_io_n1178, top_core_io_n1177, top_core_io_n1176,
         top_core_io_n1175, top_core_io_n1174, top_core_io_n1173,
         top_core_io_n1172, top_core_io_n1171, top_core_io_n1170,
         top_core_io_n1169, top_core_io_n1168, top_core_io_n1167,
         top_core_io_n1166, top_core_io_n1165, top_core_io_n1164,
         top_core_io_n1163, top_core_io_n1162, top_core_io_n1161,
         top_core_io_n1160, top_core_io_n1159, top_core_io_n1158,
         top_core_io_n1157, top_core_io_n1156, top_core_io_n1155,
         top_core_io_n1154, top_core_io_n1153, top_core_io_n1152,
         top_core_io_n1151, top_core_io_n1150, top_core_io_n1149,
         top_core_io_n1148, top_core_io_n1147, top_core_io_n1146,
         top_core_io_n1145, top_core_io_n1144, top_core_io_n1143,
         top_core_io_n1142, top_core_io_n1141, top_core_io_n1140,
         top_core_io_n1139, top_core_io_n1138, top_core_io_n1137,
         top_core_io_n1136, top_core_io_n1135, top_core_io_n1134,
         top_core_io_n1133, top_core_io_n1132, top_core_io_n1131,
         top_core_io_n1130, top_core_io_n1129, top_core_io_n1128,
         top_core_io_n1127, top_core_io_n1126, top_core_io_n1125,
         top_core_io_n1124, top_core_io_n1123, top_core_io_n1122,
         top_core_io_n1121, top_core_io_n1120, top_core_io_n1119,
         top_core_io_n1118, top_core_io_n1117, top_core_io_n1116,
         top_core_io_n1115, top_core_io_n1114, top_core_io_n1113,
         top_core_io_n1112, top_core_io_n1111, top_core_io_n1110,
         top_core_io_n1109, top_core_io_n1108, top_core_io_n1107,
         top_core_io_n1106, top_core_io_n1105, top_core_io_n1104,
         top_core_io_n1103, top_core_io_n1102, top_core_io_n1101,
         top_core_io_n1100, top_core_io_n1099, top_core_io_n1098,
         top_core_io_n1097, top_core_io_n1096, top_core_io_n1095,
         top_core_io_n1094, top_core_io_n1093, top_core_io_n1092,
         top_core_io_n1091, top_core_io_n1090, top_core_io_n1089,
         top_core_io_n1088, top_core_io_n1087, top_core_io_n1086,
         top_core_io_n1085, top_core_io_n1084, top_core_io_n1083,
         top_core_io_n1082, top_core_io_n1081, top_core_io_n1080,
         top_core_io_n1079, top_core_io_n1078, top_core_io_n1077,
         top_core_io_n1076, top_core_io_n1075, top_core_io_n1074,
         top_core_io_n1073, top_core_io_n1072, top_core_io_n1071,
         top_core_io_n1070, top_core_io_n1069, top_core_io_n1068,
         top_core_io_n1067, top_core_io_n1066, top_core_io_n1065,
         top_core_io_n1064, top_core_io_n1063, top_core_io_n1062,
         top_core_io_n1061, top_core_io_n1060, top_core_io_n1059,
         top_core_io_n1058, top_core_io_n1057, top_core_io_n1056,
         top_core_io_n1055, top_core_io_n1054, top_core_io_n1053,
         top_core_io_n1052, top_core_io_n1051, top_core_io_n922,
         top_core_io_n921, top_core_io_n920, top_core_io_n919,
         top_core_io_n918, top_core_io_n917, top_core_io_n916,
         top_core_io_n915, top_core_io_n914, top_core_io_n913,
         top_core_io_n912, top_core_io_n911, top_core_io_n910,
         top_core_io_n909, top_core_io_n908, top_core_io_n907,
         top_core_io_n906, top_core_io_n905, top_core_io_n904,
         top_core_io_n903, top_core_io_n902, top_core_io_n901,
         top_core_io_n900, top_core_io_n899, top_core_io_n898,
         top_core_io_n897, top_core_io_n896, top_core_io_n895,
         top_core_io_n894, top_core_io_n893, top_core_io_n892,
         top_core_io_n891, top_core_io_n890, top_core_io_n889,
         top_core_io_n888, top_core_io_n887, top_core_io_n886,
         top_core_io_n885, top_core_io_n884, top_core_io_n883,
         top_core_io_n882, top_core_io_n881, top_core_io_n880,
         top_core_io_n879, top_core_io_n878, top_core_io_n877,
         top_core_io_n876, top_core_io_n875, top_core_io_n874,
         top_core_io_n873, top_core_io_n872, top_core_io_n871,
         top_core_io_n870, top_core_io_n869, top_core_io_n868,
         top_core_io_n867, top_core_io_n866, top_core_io_n865,
         top_core_io_n864, top_core_io_n863, top_core_io_n862,
         top_core_io_n861, top_core_io_n860, top_core_io_n859,
         top_core_io_n858, top_core_io_n857, top_core_io_n856,
         top_core_io_n855, top_core_io_n854, top_core_io_n853,
         top_core_io_n852, top_core_io_n851, top_core_io_n850,
         top_core_io_n849, top_core_io_n848, top_core_io_n847,
         top_core_io_n846, top_core_io_n845, top_core_io_n844,
         top_core_io_n843, top_core_io_n842, top_core_io_n841,
         top_core_io_n840, top_core_io_n839, top_core_io_n838,
         top_core_io_n837, top_core_io_n836, top_core_io_n835,
         top_core_io_n834, top_core_io_n833, top_core_io_n832,
         top_core_io_n831, top_core_io_n830, top_core_io_n829,
         top_core_io_n828, top_core_io_n827, top_core_io_n826,
         top_core_io_n825, top_core_io_n824, top_core_io_n823,
         top_core_io_n822, top_core_io_n821, top_core_io_n820,
         top_core_io_n819, top_core_io_n818, top_core_io_n817,
         top_core_io_n816, top_core_io_n815, top_core_io_n814,
         top_core_io_n813, top_core_io_n812, top_core_io_n811,
         top_core_io_n810, top_core_io_n809, top_core_io_n808,
         top_core_io_n807, top_core_io_n806, top_core_io_n805,
         top_core_io_n804, top_core_io_n803, top_core_io_n802,
         top_core_io_n801, top_core_io_n800, top_core_io_n799,
         top_core_io_n798, top_core_io_n797, top_core_io_n796,
         top_core_io_n795, top_core_io_n794, top_core_io_n793,
         top_core_io_n792, top_core_io_n791, top_core_io_n790,
         top_core_io_n789, top_core_io_n788, top_core_io_n787,
         top_core_io_n786, top_core_io_n785, top_core_io_n784,
         top_core_io_n783, top_core_io_n782, top_core_io_n781,
         top_core_io_n780, top_core_io_n779, top_core_io_n778,
         top_core_io_n777, top_core_io_n776, top_core_io_n775,
         top_core_io_n774, top_core_io_n773, top_core_io_n772,
         top_core_io_n771, top_core_io_n770, top_core_io_n769,
         top_core_io_n768, top_core_io_n767, top_core_io_n766,
         top_core_io_n765, top_core_io_n764, top_core_io_n763,
         top_core_io_n762, top_core_io_n761, top_core_io_n760,
         top_core_io_n759, top_core_io_n758, top_core_io_n757,
         top_core_io_n756, top_core_io_n755, top_core_io_n754,
         top_core_io_n753, top_core_io_n752, top_core_io_n751,
         top_core_io_n750, top_core_io_n749, top_core_io_n748,
         top_core_io_n747, top_core_io_n746, top_core_io_n745,
         top_core_io_n744, top_core_io_n743, top_core_io_n742,
         top_core_io_n741, top_core_io_n740, top_core_io_n739,
         top_core_io_n738, top_core_io_n737, top_core_io_n736,
         top_core_io_n735, top_core_io_n734, top_core_io_n733,
         top_core_io_n732, top_core_io_n731, top_core_io_n730,
         top_core_io_n729, top_core_io_n728, top_core_io_n727,
         top_core_io_n726, top_core_io_n725, top_core_io_n724,
         top_core_io_n723, top_core_io_n722, top_core_io_n721,
         top_core_io_n720, top_core_io_n719, top_core_io_n718,
         top_core_io_n717, top_core_io_n716, top_core_io_n715,
         top_core_io_n714, top_core_io_n713, top_core_io_n712,
         top_core_io_n711, top_core_io_n710, top_core_io_n709,
         top_core_io_n708, top_core_io_n707, top_core_io_n706,
         top_core_io_n705, top_core_io_n704, top_core_io_n703,
         top_core_io_n702, top_core_io_n701, top_core_io_n700,
         top_core_io_n699, top_core_io_n698, top_core_io_n697,
         top_core_io_n696, top_core_io_n695, top_core_io_n694,
         top_core_io_n693, top_core_io_n692, top_core_io_n691,
         top_core_io_n690, top_core_io_n689, top_core_io_n688,
         top_core_io_n687, top_core_io_n686, top_core_io_n685,
         top_core_io_n684, top_core_io_n683, top_core_io_n682,
         top_core_io_n681, top_core_io_n680, top_core_io_n679,
         top_core_io_n678, top_core_io_n677, top_core_io_n676,
         top_core_io_n675, top_core_io_n674, top_core_io_n673,
         top_core_io_n672, top_core_io_n671, top_core_io_n670,
         top_core_io_n669, top_core_io_n668, top_core_io_n667,
         top_core_io_n666, top_core_io_n665, top_core_io_n664,
         top_core_io_n663, top_core_io_n661, top_core_io_n660,
         top_core_io_n659, top_core_io_n657, top_core_io_n656,
         top_core_io_n655, top_core_io_n653, top_core_io_n621,
         top_core_io_n528, top_core_io_n517, top_core_io_n506,
         top_core_io_n495, top_core_io_n484, top_core_io_n483,
         top_core_io_n482, top_core_io_n481, top_core_io_n480,
         top_core_io_n479, top_core_io_n478, top_core_io_n477,
         top_core_io_n476, top_core_io_n475, top_core_io_n474,
         top_core_io_n473, top_core_io_n472, top_core_io_n471,
         top_core_io_n470, top_core_io_n469, top_core_io_n468,
         top_core_io_n467, top_core_io_n466, top_core_io_n465,
         top_core_io_n464, top_core_io_n463, top_core_io_n462,
         top_core_io_n461, top_core_io_n460, top_core_io_n459,
         top_core_io_n458, top_core_io_n457, top_core_io_n456,
         top_core_io_n455, top_core_io_n454, top_core_io_n453,
         top_core_io_n452, top_core_io_n451, top_core_io_n450,
         top_core_io_n449, top_core_io_n448, top_core_io_n447,
         top_core_io_n446, top_core_io_n445, top_core_io_n444,
         top_core_io_n443, top_core_io_n442, top_core_io_n441,
         top_core_io_n440, top_core_io_n439, top_core_io_n438,
         top_core_io_n437, top_core_io_n436, top_core_io_n435,
         top_core_io_n434, top_core_io_n433, top_core_io_n432,
         top_core_io_n431, top_core_io_n430, top_core_io_n429,
         top_core_io_n428, top_core_io_n427, top_core_io_n426,
         top_core_io_n425, top_core_io_n424, top_core_io_n423,
         top_core_io_n422, top_core_io_n421, top_core_io_n420,
         top_core_io_n419, top_core_io_n418, top_core_io_n417,
         top_core_io_n416, top_core_io_n415, top_core_io_n414,
         top_core_io_n413, top_core_io_n412, top_core_io_n411,
         top_core_io_n410, top_core_io_n409, top_core_io_n408,
         top_core_io_n407, top_core_io_n406, top_core_io_n405,
         top_core_io_n404, top_core_io_n403, top_core_io_n402,
         top_core_io_n401, top_core_io_n400, top_core_io_n399,
         top_core_io_n398, top_core_io_n397, top_core_io_n396,
         top_core_io_n395, top_core_io_n394, top_core_io_n393,
         top_core_io_n392, top_core_io_n391, top_core_io_n390,
         top_core_io_n389, top_core_io_n388, top_core_io_n387,
         top_core_io_n386, top_core_io_n385, top_core_io_n384,
         top_core_io_n383, top_core_io_n382, top_core_io_n381,
         top_core_io_n380, top_core_io_n379, top_core_io_n378,
         top_core_io_n377, top_core_io_n376, top_core_io_n375,
         top_core_io_n374, top_core_io_n373, top_core_io_n372,
         top_core_io_n371, top_core_io_n370, top_core_io_n369,
         top_core_io_n368, top_core_io_n367, top_core_io_n366,
         top_core_io_n365, top_core_io_n364, top_core_io_n363,
         top_core_io_n362, top_core_io_n361, top_core_io_n360,
         top_core_io_n359, top_core_io_n358, top_core_io_n356,
         top_core_io_n324, top_core_io_n233, top_core_io_n222,
         top_core_io_n211, top_core_io_n200, top_core_io_n189,
         top_core_io_n188, top_core_io_n177, top_core_io_n166,
         top_core_io_n155, top_core_io_n154, top_core_io_n60, top_core_io_n49,
         top_core_io_n38, top_core_io_n27, top_core_io_n5, top_core_io_n1,
         top_core_io_N515, top_core_io_N514, top_core_io_N513,
         top_core_io_N512, top_core_io_N511, top_core_io_N510,
         top_core_io_N509, top_core_io_N508, top_core_io_N507,
         top_core_io_N506, top_core_io_N505, top_core_io_N504,
         top_core_io_N503, top_core_io_N502, top_core_io_N501,
         top_core_io_N500, top_core_io_N499, top_core_io_N498,
         top_core_io_N497, top_core_io_N496, top_core_io_N495,
         top_core_io_N494, top_core_io_N493, top_core_io_N492,
         top_core_io_N491, top_core_io_N490, top_core_io_N489,
         top_core_io_N488, top_core_io_N487, top_core_io_N486,
         top_core_io_N485, top_core_io_N484, top_core_io_N483,
         top_core_io_N482, top_core_io_N481, top_core_io_N480,
         top_core_io_N479, top_core_io_N478, top_core_io_N477,
         top_core_io_N476, top_core_io_N475, top_core_io_N474,
         top_core_io_N473, top_core_io_N472, top_core_io_N471,
         top_core_io_N470, top_core_io_N469, top_core_io_N468,
         top_core_io_N467, top_core_io_N466, top_core_io_N465,
         top_core_io_N464, top_core_io_N463, top_core_io_N462,
         top_core_io_N461, top_core_io_N460, top_core_io_N459,
         top_core_io_N458, top_core_io_N457, top_core_io_N456,
         top_core_io_N455, top_core_io_N454, top_core_io_N453,
         top_core_io_N452, top_core_io_N451, top_core_io_N450,
         top_core_io_N449, top_core_io_N448, top_core_io_N447,
         top_core_io_N446, top_core_io_N445, top_core_io_N444,
         top_core_io_N443, top_core_io_N442, top_core_io_N441,
         top_core_io_N440, top_core_io_N439, top_core_io_N438,
         top_core_io_N437, top_core_io_N436, top_core_io_N435,
         top_core_io_N434, top_core_io_N433, top_core_io_N432,
         top_core_io_N431, top_core_io_N430, top_core_io_N429,
         top_core_io_N428, top_core_io_N427, top_core_io_N426,
         top_core_io_N425, top_core_io_N424, top_core_io_N423,
         top_core_io_N422, top_core_io_N421, top_core_io_N420,
         top_core_io_N419, top_core_io_N418, top_core_io_N417,
         top_core_io_N416, top_core_io_N415, top_core_io_N414,
         top_core_io_N413, top_core_io_N412, top_core_io_N411,
         top_core_io_N410, top_core_io_N409, top_core_io_N408,
         top_core_io_N407, top_core_io_N406, top_core_io_N405,
         top_core_io_N404, top_core_io_N403, top_core_io_N402,
         top_core_io_N401, top_core_io_N400, top_core_io_N399,
         top_core_io_N398, top_core_io_N397, top_core_io_N396,
         top_core_io_N395, top_core_io_N394, top_core_io_N393,
         top_core_io_N392, top_core_io_N391, top_core_io_N390,
         top_core_io_N389, top_core_io_N388, top_core_io_N387,
         top_core_io_N386, top_core_io_N385, top_core_io_N384,
         top_core_io_N383, top_core_io_N382, top_core_io_N381,
         top_core_io_N380, top_core_io_N379, top_core_io_N378,
         top_core_io_N377, top_core_io_N376, top_core_io_N375,
         top_core_io_N374, top_core_io_N373, top_core_io_N372,
         top_core_io_N371, top_core_io_N370, top_core_io_N369,
         top_core_io_N368, top_core_io_N367, top_core_io_N366,
         top_core_io_N365, top_core_io_N364, top_core_io_N363,
         top_core_io_N362, top_core_io_N361, top_core_io_N360,
         top_core_io_N359, top_core_io_N358, top_core_io_N357,
         top_core_io_N356, top_core_io_N355, top_core_io_N354,
         top_core_io_N353, top_core_io_N352, top_core_io_N351,
         top_core_io_N350, top_core_io_N349, top_core_io_N348,
         top_core_io_N347, top_core_io_N346, top_core_io_N345,
         top_core_io_N344, top_core_io_N343, top_core_io_N342,
         top_core_io_N341, top_core_io_N340, top_core_io_N339,
         top_core_io_N338, top_core_io_N337, top_core_io_N336,
         top_core_io_N335, top_core_io_N334, top_core_io_N333,
         top_core_io_N332, top_core_io_N331, top_core_io_N330,
         top_core_io_N329, top_core_io_N328, top_core_io_N327,
         top_core_io_N326, top_core_io_N325, top_core_io_N324,
         top_core_io_N323, top_core_io_N322, top_core_io_N321,
         top_core_io_N320, top_core_io_N319, top_core_io_N318,
         top_core_io_N317, top_core_io_N316, top_core_io_N315,
         top_core_io_N314, top_core_io_N313, top_core_io_N312,
         top_core_io_N311, top_core_io_N310, top_core_io_N309,
         top_core_io_N308, top_core_io_N307, top_core_io_N306,
         top_core_io_N305, top_core_io_N304, top_core_io_N303,
         top_core_io_N302, top_core_io_N301, top_core_io_N300,
         top_core_io_N299, top_core_io_N298, top_core_io_N297,
         top_core_io_N296, top_core_io_N295, top_core_io_N294,
         top_core_io_N293, top_core_io_N292, top_core_io_N291,
         top_core_io_N290, top_core_io_N289, top_core_io_N288,
         top_core_io_N287, top_core_io_N286, top_core_io_N285,
         top_core_io_N284, top_core_io_N283, top_core_io_N282,
         top_core_io_N281, top_core_io_N280, top_core_io_N279,
         top_core_io_N278, top_core_io_N277, top_core_io_N276,
         top_core_io_N275, top_core_io_N274, top_core_io_N273,
         top_core_io_N272, top_core_io_N271, top_core_io_N270,
         top_core_io_N269, top_core_io_N268, top_core_io_N267,
         top_core_io_N266, top_core_io_N265, top_core_io_N264,
         top_core_io_N263, top_core_io_N262, top_core_io_N261,
         top_core_io_N260, top_core_io_N259, top_core_io_N258,
         top_core_io_N257, top_core_io_N256, top_core_io_N255,
         top_core_io_N254, top_core_io_N253, top_core_io_N252,
         top_core_io_N251, top_core_io_N250, top_core_io_N249,
         top_core_io_N248, top_core_io_N247, top_core_io_N246,
         top_core_io_N245, top_core_io_N244, top_core_io_N243,
         top_core_io_N242, top_core_io_N241, top_core_io_N240,
         top_core_io_N239, top_core_io_N238, top_core_io_N237,
         top_core_io_N236, top_core_io_N235, top_core_io_N234,
         top_core_io_N233, top_core_io_N232, top_core_io_N231,
         top_core_io_N230, top_core_io_N229, top_core_io_N228,
         top_core_io_N227, top_core_io_N226, top_core_io_N225,
         top_core_io_N224, top_core_io_N223, top_core_io_N222,
         top_core_io_N221, top_core_io_N220, top_core_io_N219,
         top_core_io_N218, top_core_io_N217, top_core_io_N216,
         top_core_io_N215, top_core_io_N214, top_core_io_N213,
         top_core_io_N212, top_core_io_N211, top_core_io_N210,
         top_core_io_N209, top_core_io_N208, top_core_io_N207,
         top_core_io_N206, top_core_io_N205, top_core_io_N204,
         top_core_io_N203, top_core_io_N202, top_core_io_N201,
         top_core_io_N200, top_core_io_N199, top_core_io_N198,
         top_core_io_N197, top_core_io_N196, top_core_io_N195,
         top_core_io_N194, top_core_io_N193, top_core_io_N192,
         top_core_io_N191, top_core_io_N190, top_core_io_N189,
         top_core_io_N188, top_core_io_N187, top_core_io_N186,
         top_core_io_N185, top_core_io_N184, top_core_io_N183,
         top_core_io_N182, top_core_io_N181, top_core_io_N180,
         top_core_io_N179, top_core_io_N178, top_core_io_N177,
         top_core_io_N176, top_core_io_N175, top_core_io_N174,
         top_core_io_N173, top_core_io_N172, top_core_io_N171,
         top_core_io_N170, top_core_io_N169, top_core_io_N168,
         top_core_io_N167, top_core_io_N166, top_core_io_N165,
         top_core_io_N164, top_core_io_N163, top_core_io_N162,
         top_core_io_N161, top_core_io_N160, top_core_io_N159,
         top_core_io_N158, top_core_io_N157, top_core_io_N156,
         top_core_io_N155, top_core_io_N154, top_core_io_N153,
         top_core_io_N152, top_core_io_N151, top_core_io_N150,
         top_core_io_N149, top_core_io_N148, top_core_io_N147,
         top_core_io_N146, top_core_io_N145, top_core_io_N144,
         top_core_io_N143, top_core_io_N142, top_core_io_N141,
         top_core_io_N140, top_core_io_N139, top_core_io_N138,
         top_core_io_N137, top_core_io_N136, top_core_io_N135,
         top_core_io_N134, top_core_io_N133, top_core_io_N132,
         top_core_io_N131, top_core_io_N127, top_core_io_N126,
         top_core_io_N125, top_core_io_inter_ok, top_core_io_N97,
         top_core_io_N96, top_core_io_N95, top_core_io_N94, top_core_io_N93,
         top_core_io_N92, top_core_io_N91, top_core_io_N90, top_core_io_N81,
         top_core_io_N80, top_core_io_N79, top_core_io_N78, top_core_io_N77,
         top_core_io_N76, top_core_io_N75, top_core_io_N74,
         top_core_io_CORE_FULL, top_core_io_NK_0_, top_core_io_NK_1_,
         top_core_io_NK_2_, top_core_io_operation, top_core_io_CipherKey_w_0_,
         top_core_io_CipherKey_w_1_, top_core_io_CipherKey_w_2_,
         top_core_io_CipherKey_w_3_, top_core_io_CipherKey_w_4_,
         top_core_io_CipherKey_w_5_, top_core_io_CipherKey_w_6_,
         top_core_io_CipherKey_w_7_, top_core_io_CipherKey_w_8_,
         top_core_io_CipherKey_w_9_, top_core_io_CipherKey_w_10_,
         top_core_io_CipherKey_w_11_, top_core_io_CipherKey_w_12_,
         top_core_io_CipherKey_w_13_, top_core_io_CipherKey_w_14_,
         top_core_io_CipherKey_w_15_, top_core_io_CipherKey_w_16_,
         top_core_io_CipherKey_w_17_, top_core_io_CipherKey_w_18_,
         top_core_io_CipherKey_w_19_, top_core_io_CipherKey_w_20_,
         top_core_io_CipherKey_w_21_, top_core_io_CipherKey_w_22_,
         top_core_io_CipherKey_w_23_, top_core_io_CipherKey_w_24_,
         top_core_io_CipherKey_w_25_, top_core_io_CipherKey_w_26_,
         top_core_io_CipherKey_w_27_, top_core_io_CipherKey_w_28_,
         top_core_io_CipherKey_w_29_, top_core_io_CipherKey_w_30_,
         top_core_io_CipherKey_w_31_, top_core_io_CipherKey_w_32_,
         top_core_io_CipherKey_w_33_, top_core_io_CipherKey_w_34_,
         top_core_io_CipherKey_w_35_, top_core_io_CipherKey_w_36_,
         top_core_io_CipherKey_w_37_, top_core_io_CipherKey_w_38_,
         top_core_io_CipherKey_w_39_, top_core_io_CipherKey_w_40_,
         top_core_io_CipherKey_w_41_, top_core_io_CipherKey_w_42_,
         top_core_io_CipherKey_w_43_, top_core_io_CipherKey_w_44_,
         top_core_io_CipherKey_w_45_, top_core_io_CipherKey_w_46_,
         top_core_io_CipherKey_w_47_, top_core_io_CipherKey_w_48_,
         top_core_io_CipherKey_w_49_, top_core_io_CipherKey_w_50_,
         top_core_io_CipherKey_w_51_, top_core_io_CipherKey_w_52_,
         top_core_io_CipherKey_w_53_, top_core_io_CipherKey_w_54_,
         top_core_io_CipherKey_w_55_, top_core_io_CipherKey_w_56_,
         top_core_io_CipherKey_w_57_, top_core_io_CipherKey_w_58_,
         top_core_io_CipherKey_w_59_, top_core_io_CipherKey_w_60_,
         top_core_io_CipherKey_w_61_, top_core_io_CipherKey_w_62_,
         top_core_io_CipherKey_w_63_, top_core_io_CipherKey_w_64_,
         top_core_io_CipherKey_w_65_, top_core_io_CipherKey_w_66_,
         top_core_io_CipherKey_w_67_, top_core_io_CipherKey_w_68_,
         top_core_io_CipherKey_w_69_, top_core_io_CipherKey_w_70_,
         top_core_io_CipherKey_w_71_, top_core_io_CipherKey_w_72_,
         top_core_io_CipherKey_w_73_, top_core_io_CipherKey_w_74_,
         top_core_io_CipherKey_w_75_, top_core_io_CipherKey_w_76_,
         top_core_io_CipherKey_w_77_, top_core_io_CipherKey_w_78_,
         top_core_io_CipherKey_w_79_, top_core_io_CipherKey_w_80_,
         top_core_io_CipherKey_w_81_, top_core_io_CipherKey_w_82_,
         top_core_io_CipherKey_w_83_, top_core_io_CipherKey_w_84_,
         top_core_io_CipherKey_w_85_, top_core_io_CipherKey_w_86_,
         top_core_io_CipherKey_w_87_, top_core_io_CipherKey_w_88_,
         top_core_io_CipherKey_w_89_, top_core_io_CipherKey_w_90_,
         top_core_io_CipherKey_w_91_, top_core_io_CipherKey_w_92_,
         top_core_io_CipherKey_w_93_, top_core_io_CipherKey_w_94_,
         top_core_io_CipherKey_w_95_, top_core_io_CipherKey_w_96_,
         top_core_io_CipherKey_w_97_, top_core_io_CipherKey_w_98_,
         top_core_io_CipherKey_w_99_, top_core_io_CipherKey_w_100_,
         top_core_io_CipherKey_w_101_, top_core_io_CipherKey_w_102_,
         top_core_io_CipherKey_w_103_, top_core_io_CipherKey_w_104_,
         top_core_io_CipherKey_w_105_, top_core_io_CipherKey_w_106_,
         top_core_io_CipherKey_w_107_, top_core_io_CipherKey_w_108_,
         top_core_io_CipherKey_w_109_, top_core_io_CipherKey_w_110_,
         top_core_io_CipherKey_w_111_, top_core_io_CipherKey_w_112_,
         top_core_io_CipherKey_w_113_, top_core_io_CipherKey_w_114_,
         top_core_io_CipherKey_w_115_, top_core_io_CipherKey_w_116_,
         top_core_io_CipherKey_w_117_, top_core_io_CipherKey_w_118_,
         top_core_io_CipherKey_w_119_, top_core_io_CipherKey_w_120_,
         top_core_io_CipherKey_w_121_, top_core_io_CipherKey_w_122_,
         top_core_io_CipherKey_w_123_, top_core_io_CipherKey_w_124_,
         top_core_io_CipherKey_w_125_, top_core_io_CipherKey_w_126_,
         top_core_io_CipherKey_w_127_, top_core_io_CipherKey_w_128_,
         top_core_io_CipherKey_w_129_, top_core_io_CipherKey_w_130_,
         top_core_io_CipherKey_w_131_, top_core_io_CipherKey_w_132_,
         top_core_io_CipherKey_w_133_, top_core_io_CipherKey_w_134_,
         top_core_io_CipherKey_w_135_, top_core_io_CipherKey_w_136_,
         top_core_io_CipherKey_w_137_, top_core_io_CipherKey_w_138_,
         top_core_io_CipherKey_w_139_, top_core_io_CipherKey_w_140_,
         top_core_io_CipherKey_w_141_, top_core_io_CipherKey_w_142_,
         top_core_io_CipherKey_w_143_, top_core_io_CipherKey_w_144_,
         top_core_io_CipherKey_w_145_, top_core_io_CipherKey_w_146_,
         top_core_io_CipherKey_w_147_, top_core_io_CipherKey_w_148_,
         top_core_io_CipherKey_w_149_, top_core_io_CipherKey_w_150_,
         top_core_io_CipherKey_w_151_, top_core_io_CipherKey_w_152_,
         top_core_io_CipherKey_w_153_, top_core_io_CipherKey_w_154_,
         top_core_io_CipherKey_w_155_, top_core_io_CipherKey_w_156_,
         top_core_io_CipherKey_w_157_, top_core_io_CipherKey_w_158_,
         top_core_io_CipherKey_w_159_, top_core_io_CipherKey_w_160_,
         top_core_io_CipherKey_w_161_, top_core_io_CipherKey_w_162_,
         top_core_io_CipherKey_w_163_, top_core_io_CipherKey_w_164_,
         top_core_io_CipherKey_w_165_, top_core_io_CipherKey_w_166_,
         top_core_io_CipherKey_w_167_, top_core_io_CipherKey_w_168_,
         top_core_io_CipherKey_w_169_, top_core_io_CipherKey_w_170_,
         top_core_io_CipherKey_w_171_, top_core_io_CipherKey_w_172_,
         top_core_io_CipherKey_w_173_, top_core_io_CipherKey_w_174_,
         top_core_io_CipherKey_w_175_, top_core_io_CipherKey_w_176_,
         top_core_io_CipherKey_w_177_, top_core_io_CipherKey_w_178_,
         top_core_io_CipherKey_w_179_, top_core_io_CipherKey_w_180_,
         top_core_io_CipherKey_w_181_, top_core_io_CipherKey_w_182_,
         top_core_io_CipherKey_w_183_, top_core_io_CipherKey_w_184_,
         top_core_io_CipherKey_w_185_, top_core_io_CipherKey_w_186_,
         top_core_io_CipherKey_w_187_, top_core_io_CipherKey_w_188_,
         top_core_io_CipherKey_w_189_, top_core_io_CipherKey_w_190_,
         top_core_io_CipherKey_w_191_, top_core_io_CipherKey_w_192_,
         top_core_io_CipherKey_w_193_, top_core_io_CipherKey_w_194_,
         top_core_io_CipherKey_w_195_, top_core_io_CipherKey_w_196_,
         top_core_io_CipherKey_w_197_, top_core_io_CipherKey_w_198_,
         top_core_io_CipherKey_w_199_, top_core_io_CipherKey_w_200_,
         top_core_io_CipherKey_w_201_, top_core_io_CipherKey_w_202_,
         top_core_io_CipherKey_w_203_, top_core_io_CipherKey_w_204_,
         top_core_io_CipherKey_w_205_, top_core_io_CipherKey_w_206_,
         top_core_io_CipherKey_w_207_, top_core_io_CipherKey_w_208_,
         top_core_io_CipherKey_w_209_, top_core_io_CipherKey_w_210_,
         top_core_io_CipherKey_w_211_, top_core_io_CipherKey_w_212_,
         top_core_io_CipherKey_w_213_, top_core_io_CipherKey_w_214_,
         top_core_io_CipherKey_w_215_, top_core_io_CipherKey_w_216_,
         top_core_io_CipherKey_w_217_, top_core_io_CipherKey_w_218_,
         top_core_io_CipherKey_w_219_, top_core_io_CipherKey_w_220_,
         top_core_io_CipherKey_w_221_, top_core_io_CipherKey_w_222_,
         top_core_io_CipherKey_w_223_, top_core_io_CipherKey_w_224_,
         top_core_io_CipherKey_w_225_, top_core_io_CipherKey_w_226_,
         top_core_io_CipherKey_w_227_, top_core_io_CipherKey_w_228_,
         top_core_io_CipherKey_w_229_, top_core_io_CipherKey_w_230_,
         top_core_io_CipherKey_w_231_, top_core_io_CipherKey_w_232_,
         top_core_io_CipherKey_w_233_, top_core_io_CipherKey_w_234_,
         top_core_io_CipherKey_w_235_, top_core_io_CipherKey_w_236_,
         top_core_io_CipherKey_w_237_, top_core_io_CipherKey_w_238_,
         top_core_io_CipherKey_w_239_, top_core_io_CipherKey_w_240_,
         top_core_io_CipherKey_w_241_, top_core_io_CipherKey_w_242_,
         top_core_io_CipherKey_w_243_, top_core_io_CipherKey_w_244_,
         top_core_io_CipherKey_w_245_, top_core_io_CipherKey_w_246_,
         top_core_io_CipherKey_w_247_, top_core_io_CipherKey_w_248_,
         top_core_io_CipherKey_w_249_, top_core_io_CipherKey_w_250_,
         top_core_io_CipherKey_w_251_, top_core_io_CipherKey_w_252_,
         top_core_io_CipherKey_w_253_, top_core_io_CipherKey_w_254_,
         top_core_io_CipherKey_w_255_, top_core_io_Plain_text_w_0_,
         top_core_io_Plain_text_w_1_, top_core_io_Plain_text_w_2_,
         top_core_io_Plain_text_w_3_, top_core_io_Plain_text_w_4_,
         top_core_io_Plain_text_w_5_, top_core_io_Plain_text_w_6_,
         top_core_io_Plain_text_w_7_, top_core_io_Plain_text_w_8_,
         top_core_io_Plain_text_w_9_, top_core_io_Plain_text_w_10_,
         top_core_io_Plain_text_w_11_, top_core_io_Plain_text_w_12_,
         top_core_io_Plain_text_w_13_, top_core_io_Plain_text_w_14_,
         top_core_io_Plain_text_w_15_, top_core_io_Plain_text_w_16_,
         top_core_io_Plain_text_w_17_, top_core_io_Plain_text_w_18_,
         top_core_io_Plain_text_w_19_, top_core_io_Plain_text_w_20_,
         top_core_io_Plain_text_w_21_, top_core_io_Plain_text_w_22_,
         top_core_io_Plain_text_w_23_, top_core_io_Plain_text_w_24_,
         top_core_io_Plain_text_w_25_, top_core_io_Plain_text_w_26_,
         top_core_io_Plain_text_w_27_, top_core_io_Plain_text_w_28_,
         top_core_io_Plain_text_w_29_, top_core_io_Plain_text_w_30_,
         top_core_io_Plain_text_w_31_, top_core_io_Plain_text_w_32_,
         top_core_io_Plain_text_w_33_, top_core_io_Plain_text_w_34_,
         top_core_io_Plain_text_w_35_, top_core_io_Plain_text_w_36_,
         top_core_io_Plain_text_w_37_, top_core_io_Plain_text_w_38_,
         top_core_io_Plain_text_w_39_, top_core_io_Plain_text_w_40_,
         top_core_io_Plain_text_w_41_, top_core_io_Plain_text_w_42_,
         top_core_io_Plain_text_w_43_, top_core_io_Plain_text_w_44_,
         top_core_io_Plain_text_w_45_, top_core_io_Plain_text_w_46_,
         top_core_io_Plain_text_w_47_, top_core_io_Plain_text_w_48_,
         top_core_io_Plain_text_w_49_, top_core_io_Plain_text_w_50_,
         top_core_io_Plain_text_w_51_, top_core_io_Plain_text_w_52_,
         top_core_io_Plain_text_w_53_, top_core_io_Plain_text_w_54_,
         top_core_io_Plain_text_w_55_, top_core_io_Plain_text_w_56_,
         top_core_io_Plain_text_w_57_, top_core_io_Plain_text_w_58_,
         top_core_io_Plain_text_w_59_, top_core_io_Plain_text_w_60_,
         top_core_io_Plain_text_w_61_, top_core_io_Plain_text_w_62_,
         top_core_io_Plain_text_w_63_, top_core_io_Plain_text_w_64_,
         top_core_io_Plain_text_w_65_, top_core_io_Plain_text_w_66_,
         top_core_io_Plain_text_w_67_, top_core_io_Plain_text_w_68_,
         top_core_io_Plain_text_w_69_, top_core_io_Plain_text_w_70_,
         top_core_io_Plain_text_w_71_, top_core_io_Plain_text_w_72_,
         top_core_io_Plain_text_w_73_, top_core_io_Plain_text_w_74_,
         top_core_io_Plain_text_w_75_, top_core_io_Plain_text_w_76_,
         top_core_io_Plain_text_w_77_, top_core_io_Plain_text_w_78_,
         top_core_io_Plain_text_w_79_, top_core_io_Plain_text_w_80_,
         top_core_io_Plain_text_w_81_, top_core_io_Plain_text_w_82_,
         top_core_io_Plain_text_w_83_, top_core_io_Plain_text_w_84_,
         top_core_io_Plain_text_w_85_, top_core_io_Plain_text_w_86_,
         top_core_io_Plain_text_w_87_, top_core_io_Plain_text_w_88_,
         top_core_io_Plain_text_w_89_, top_core_io_Plain_text_w_90_,
         top_core_io_Plain_text_w_91_, top_core_io_Plain_text_w_92_,
         top_core_io_Plain_text_w_93_, top_core_io_Plain_text_w_94_,
         top_core_io_Plain_text_w_95_, top_core_io_Plain_text_w_96_,
         top_core_io_Plain_text_w_97_, top_core_io_Plain_text_w_98_,
         top_core_io_Plain_text_w_99_, top_core_io_Plain_text_w_100_,
         top_core_io_Plain_text_w_101_, top_core_io_Plain_text_w_102_,
         top_core_io_Plain_text_w_103_, top_core_io_Plain_text_w_104_,
         top_core_io_Plain_text_w_105_, top_core_io_Plain_text_w_106_,
         top_core_io_Plain_text_w_107_, top_core_io_Plain_text_w_108_,
         top_core_io_Plain_text_w_109_, top_core_io_Plain_text_w_110_,
         top_core_io_Plain_text_w_111_, top_core_io_Plain_text_w_112_,
         top_core_io_Plain_text_w_113_, top_core_io_Plain_text_w_114_,
         top_core_io_Plain_text_w_115_, top_core_io_Plain_text_w_116_,
         top_core_io_Plain_text_w_117_, top_core_io_Plain_text_w_118_,
         top_core_io_Plain_text_w_119_, top_core_io_Plain_text_w_120_,
         top_core_io_Plain_text_w_121_, top_core_io_Plain_text_w_122_,
         top_core_io_Plain_text_w_123_, top_core_io_Plain_text_w_124_,
         top_core_io_Plain_text_w_125_, top_core_io_Plain_text_w_126_,
         top_core_io_Plain_text_w_127_, top_core_io_Data_reg_16__0_,
         top_core_io_Data_reg_16__1_, top_core_io_Data_reg_16__2_,
         top_core_io_Data_reg_16__3_, top_core_io_Data_reg_16__4_,
         top_core_io_Data_reg_16__5_, top_core_io_Data_reg_16__6_,
         top_core_io_Data_reg_16__7_, top_core_io_Data_reg_17__0_,
         top_core_io_Data_reg_17__1_, top_core_io_Data_reg_17__2_,
         top_core_io_Data_reg_17__3_, top_core_io_Data_reg_17__4_,
         top_core_io_Data_reg_17__5_, top_core_io_Data_reg_17__6_,
         top_core_io_Data_reg_17__7_, top_core_io_Data_reg_18__0_,
         top_core_io_Data_reg_18__1_, top_core_io_Data_reg_18__2_,
         top_core_io_Data_reg_18__3_, top_core_io_Data_reg_18__4_,
         top_core_io_Data_reg_18__5_, top_core_io_Data_reg_18__6_,
         top_core_io_Data_reg_18__7_, top_core_io_Data_reg_19__0_,
         top_core_io_Data_reg_19__1_, top_core_io_Data_reg_19__2_,
         top_core_io_Data_reg_19__3_, top_core_io_Data_reg_19__4_,
         top_core_io_Data_reg_19__5_, top_core_io_Data_reg_19__6_,
         top_core_io_Data_reg_19__7_, top_core_io_Data_reg_20__0_,
         top_core_io_Data_reg_20__1_, top_core_io_Data_reg_20__2_,
         top_core_io_Data_reg_20__3_, top_core_io_Data_reg_20__4_,
         top_core_io_Data_reg_20__5_, top_core_io_Data_reg_20__6_,
         top_core_io_Data_reg_20__7_, top_core_io_Data_reg_21__0_,
         top_core_io_Data_reg_21__1_, top_core_io_Data_reg_21__2_,
         top_core_io_Data_reg_21__3_, top_core_io_Data_reg_21__4_,
         top_core_io_Data_reg_21__5_, top_core_io_Data_reg_21__6_,
         top_core_io_Data_reg_21__7_, top_core_io_Data_reg_22__0_,
         top_core_io_Data_reg_22__1_, top_core_io_Data_reg_22__2_,
         top_core_io_Data_reg_22__3_, top_core_io_Data_reg_22__4_,
         top_core_io_Data_reg_22__5_, top_core_io_Data_reg_22__6_,
         top_core_io_Data_reg_22__7_, top_core_io_Data_reg_23__0_,
         top_core_io_Data_reg_23__1_, top_core_io_Data_reg_23__2_,
         top_core_io_Data_reg_23__3_, top_core_io_Data_reg_23__4_,
         top_core_io_Data_reg_23__5_, top_core_io_Data_reg_23__6_,
         top_core_io_Data_reg_23__7_, top_core_io_Data_reg_24__0_,
         top_core_io_Data_reg_24__1_, top_core_io_Data_reg_24__2_,
         top_core_io_Data_reg_24__3_, top_core_io_Data_reg_24__4_,
         top_core_io_Data_reg_24__5_, top_core_io_Data_reg_24__6_,
         top_core_io_Data_reg_24__7_, top_core_io_Data_reg_25__0_,
         top_core_io_Data_reg_25__1_, top_core_io_Data_reg_25__2_,
         top_core_io_Data_reg_25__3_, top_core_io_Data_reg_25__4_,
         top_core_io_Data_reg_25__5_, top_core_io_Data_reg_25__6_,
         top_core_io_Data_reg_25__7_, top_core_io_Data_reg_26__0_,
         top_core_io_Data_reg_26__1_, top_core_io_Data_reg_26__2_,
         top_core_io_Data_reg_26__3_, top_core_io_Data_reg_26__4_,
         top_core_io_Data_reg_26__5_, top_core_io_Data_reg_26__6_,
         top_core_io_Data_reg_26__7_, top_core_io_Data_reg_27__0_,
         top_core_io_Data_reg_27__1_, top_core_io_Data_reg_27__2_,
         top_core_io_Data_reg_27__3_, top_core_io_Data_reg_27__4_,
         top_core_io_Data_reg_27__5_, top_core_io_Data_reg_27__6_,
         top_core_io_Data_reg_27__7_, top_core_io_Data_reg_28__0_,
         top_core_io_Data_reg_28__1_, top_core_io_Data_reg_28__2_,
         top_core_io_Data_reg_28__3_, top_core_io_Data_reg_28__4_,
         top_core_io_Data_reg_28__5_, top_core_io_Data_reg_28__6_,
         top_core_io_Data_reg_28__7_, top_core_io_Data_reg_29__0_,
         top_core_io_Data_reg_29__1_, top_core_io_Data_reg_29__2_,
         top_core_io_Data_reg_29__3_, top_core_io_Data_reg_29__4_,
         top_core_io_Data_reg_29__5_, top_core_io_Data_reg_29__6_,
         top_core_io_Data_reg_29__7_, top_core_io_Data_reg_30__0_,
         top_core_io_Data_reg_30__1_, top_core_io_Data_reg_30__2_,
         top_core_io_Data_reg_30__3_, top_core_io_Data_reg_30__4_,
         top_core_io_Data_reg_30__5_, top_core_io_Data_reg_30__6_,
         top_core_io_Data_reg_30__7_, top_core_io_Data_reg_31__0_,
         top_core_io_Data_reg_31__1_, top_core_io_Data_reg_31__2_,
         top_core_io_Data_reg_31__3_, top_core_io_Data_reg_31__4_,
         top_core_io_Data_reg_31__5_, top_core_io_Data_reg_31__6_,
         top_core_io_Data_reg_31__7_, top_core_EC_n1299, top_core_EC_n1298,
         top_core_EC_n1297, top_core_EC_n1296, top_core_EC_n1295,
         top_core_EC_n1294, top_core_EC_n1293, top_core_EC_n1292,
         top_core_EC_n1291, top_core_EC_n1290, top_core_EC_n1289,
         top_core_EC_n1288, top_core_EC_n1287, top_core_EC_n1286,
         top_core_EC_n1285, top_core_EC_n1284, top_core_EC_n1283,
         top_core_EC_n1282, top_core_EC_n1281, top_core_EC_n1280,
         top_core_EC_n1279, top_core_EC_n1278, top_core_EC_n1277,
         top_core_EC_n1276, top_core_EC_n1275, top_core_EC_n1274,
         top_core_EC_n1273, top_core_EC_n1272, top_core_EC_n1271,
         top_core_EC_n1270, top_core_EC_n1269, top_core_EC_n1268,
         top_core_EC_n1267, top_core_EC_n1266, top_core_EC_n1265,
         top_core_EC_n1264, top_core_EC_n1263, top_core_EC_n1262,
         top_core_EC_n1261, top_core_EC_n1260, top_core_EC_n1259,
         top_core_EC_n1258, top_core_EC_n1257, top_core_EC_n1256,
         top_core_EC_n1255, top_core_EC_n1254, top_core_EC_n1253,
         top_core_EC_n1252, top_core_EC_n1251, top_core_EC_n1250,
         top_core_EC_n1249, top_core_EC_n1248, top_core_EC_n1247,
         top_core_EC_n1246, top_core_EC_n1245, top_core_EC_n1244,
         top_core_EC_n1243, top_core_EC_n1242, top_core_EC_n1241,
         top_core_EC_n1240, top_core_EC_n1239, top_core_EC_n1238,
         top_core_EC_n1237, top_core_EC_n1236, top_core_EC_n1235,
         top_core_EC_n1234, top_core_EC_n1233, top_core_EC_n1232,
         top_core_EC_n1231, top_core_EC_n1230, top_core_EC_n1229,
         top_core_EC_n1228, top_core_EC_n1227, top_core_EC_n1226,
         top_core_EC_n1225, top_core_EC_n1224, top_core_EC_n1223,
         top_core_EC_n1222, top_core_EC_n1221, top_core_EC_n1220,
         top_core_EC_n1219, top_core_EC_n1218, top_core_EC_n1217,
         top_core_EC_n1216, top_core_EC_n1215, top_core_EC_n1214,
         top_core_EC_n1213, top_core_EC_n1212, top_core_EC_n1211,
         top_core_EC_n1210, top_core_EC_n1209, top_core_EC_n1208,
         top_core_EC_n1207, top_core_EC_n1206, top_core_EC_n1205,
         top_core_EC_n1204, top_core_EC_n1203, top_core_EC_n1202,
         top_core_EC_n1201, top_core_EC_n1200, top_core_EC_n1199,
         top_core_EC_n1198, top_core_EC_n1197, top_core_EC_n1196,
         top_core_EC_n1195, top_core_EC_n1194, top_core_EC_n1193,
         top_core_EC_n1192, top_core_EC_n1191, top_core_EC_n1190,
         top_core_EC_n1189, top_core_EC_n1188, top_core_EC_n1187,
         top_core_EC_n1186, top_core_EC_n1185, top_core_EC_n1184,
         top_core_EC_n1183, top_core_EC_n1182, top_core_EC_n1181,
         top_core_EC_n1180, top_core_EC_n1179, top_core_EC_n1178,
         top_core_EC_n1177, top_core_EC_n1176, top_core_EC_n1175,
         top_core_EC_n1174, top_core_EC_n1173, top_core_EC_n1172,
         top_core_EC_n1171, top_core_EC_n1170, top_core_EC_n1169,
         top_core_EC_n1168, top_core_EC_n1167, top_core_EC_n1166,
         top_core_EC_n1165, top_core_EC_n1164, top_core_EC_n1163,
         top_core_EC_n1162, top_core_EC_n1161, top_core_EC_n1160,
         top_core_EC_n1159, top_core_EC_n1158, top_core_EC_n1157,
         top_core_EC_n1156, top_core_EC_n1155, top_core_EC_n1154,
         top_core_EC_n1153, top_core_EC_n1152, top_core_EC_n1151,
         top_core_EC_n1150, top_core_EC_n1149, top_core_EC_n1148,
         top_core_EC_n1147, top_core_EC_n1146, top_core_EC_n1145,
         top_core_EC_n1144, top_core_EC_n1143, top_core_EC_n1142,
         top_core_EC_n1141, top_core_EC_n1140, top_core_EC_n1139,
         top_core_EC_n1138, top_core_EC_n1137, top_core_EC_n1136,
         top_core_EC_n1135, top_core_EC_n1134, top_core_EC_n1133,
         top_core_EC_n1132, top_core_EC_n1131, top_core_EC_n1130,
         top_core_EC_n1129, top_core_EC_n1128, top_core_EC_n1127,
         top_core_EC_n1126, top_core_EC_n1125, top_core_EC_n1124,
         top_core_EC_n1123, top_core_EC_n1122, top_core_EC_n1121,
         top_core_EC_n1120, top_core_EC_n1119, top_core_EC_n1118,
         top_core_EC_n1117, top_core_EC_n1116, top_core_EC_n1115,
         top_core_EC_n1114, top_core_EC_n1113, top_core_EC_n1112,
         top_core_EC_n1111, top_core_EC_n1110, top_core_EC_n1109,
         top_core_EC_n1108, top_core_EC_n1107, top_core_EC_n1106,
         top_core_EC_n1105, top_core_EC_n1104, top_core_EC_n1103,
         top_core_EC_n1102, top_core_EC_n1101, top_core_EC_n1100,
         top_core_EC_n1099, top_core_EC_n1098, top_core_EC_n1097,
         top_core_EC_n1096, top_core_EC_n1095, top_core_EC_n1094,
         top_core_EC_n1093, top_core_EC_n1092, top_core_EC_n1091,
         top_core_EC_n1090, top_core_EC_n1089, top_core_EC_n1088,
         top_core_EC_n1087, top_core_EC_n1086, top_core_EC_n1085,
         top_core_EC_n1084, top_core_EC_n1083, top_core_EC_n1082,
         top_core_EC_n1081, top_core_EC_n1080, top_core_EC_n1079,
         top_core_EC_n1078, top_core_EC_n1077, top_core_EC_n1076,
         top_core_EC_n1075, top_core_EC_n1074, top_core_EC_n1073,
         top_core_EC_n1072, top_core_EC_n1071, top_core_EC_n1070,
         top_core_EC_n1069, top_core_EC_n1068, top_core_EC_n1067,
         top_core_EC_n1066, top_core_EC_n1065, top_core_EC_n1064,
         top_core_EC_n1063, top_core_EC_n1062, top_core_EC_n1061,
         top_core_EC_n1060, top_core_EC_n1059, top_core_EC_n1058,
         top_core_EC_n1057, top_core_EC_n1056, top_core_EC_n1055,
         top_core_EC_n1054, top_core_EC_n1053, top_core_EC_n1052,
         top_core_EC_n1051, top_core_EC_n1050, top_core_EC_n1049,
         top_core_EC_n1048, top_core_EC_n1047, top_core_EC_n1046,
         top_core_EC_n1045, top_core_EC_n1044, top_core_EC_n1043,
         top_core_EC_n1042, top_core_EC_n1041, top_core_EC_n1040,
         top_core_EC_n1039, top_core_EC_n1038, top_core_EC_n1037,
         top_core_EC_n1036, top_core_EC_n1035, top_core_EC_n1034,
         top_core_EC_n1033, top_core_EC_n1027, top_core_EC_n1026,
         top_core_EC_n1025, top_core_EC_n1024, top_core_EC_n1023,
         top_core_EC_n1022, top_core_EC_n1021, top_core_EC_n1020,
         top_core_EC_n1019, top_core_EC_n1018, top_core_EC_n1017,
         top_core_EC_n1016, top_core_EC_n1015, top_core_EC_n1014,
         top_core_EC_n1013, top_core_EC_n1012, top_core_EC_n1011,
         top_core_EC_n1009, top_core_EC_n1008, top_core_EC_n1007,
         top_core_EC_n1006, top_core_EC_n1005, top_core_EC_n1004,
         top_core_EC_n1003, top_core_EC_n1002, top_core_EC_n1001,
         top_core_EC_n1000, top_core_EC_n999, top_core_EC_n998,
         top_core_EC_n997, top_core_EC_n996, top_core_EC_n995,
         top_core_EC_n994, top_core_EC_n993, top_core_EC_n992,
         top_core_EC_n991, top_core_EC_n990, top_core_EC_n989,
         top_core_EC_n988, top_core_EC_n987, top_core_EC_n986,
         top_core_EC_n985, top_core_EC_n984, top_core_EC_n983,
         top_core_EC_n982, top_core_EC_n981, top_core_EC_n980,
         top_core_EC_n979, top_core_EC_n978, top_core_EC_n977,
         top_core_EC_n976, top_core_EC_n975, top_core_EC_n974,
         top_core_EC_n973, top_core_EC_n972, top_core_EC_n971,
         top_core_EC_n970, top_core_EC_n969, top_core_EC_n968,
         top_core_EC_n967, top_core_EC_n966, top_core_EC_n965,
         top_core_EC_n964, top_core_EC_n963, top_core_EC_n962,
         top_core_EC_n961, top_core_EC_n960, top_core_EC_n959,
         top_core_EC_n958, top_core_EC_n957, top_core_EC_n956,
         top_core_EC_n955, top_core_EC_n954, top_core_EC_n953,
         top_core_EC_n952, top_core_EC_n951, top_core_EC_n950,
         top_core_EC_n949, top_core_EC_n948, top_core_EC_n947,
         top_core_EC_n946, top_core_EC_n944, top_core_EC_n943,
         top_core_EC_n942, top_core_EC_n941, top_core_EC_n940,
         top_core_EC_n939, top_core_EC_n938, top_core_EC_n937,
         top_core_EC_n936, top_core_EC_n935, top_core_EC_n934,
         top_core_EC_n933, top_core_EC_n932, top_core_EC_n931,
         top_core_EC_n930, top_core_EC_n929, top_core_EC_n928,
         top_core_EC_n927, top_core_EC_n926, top_core_EC_n925,
         top_core_EC_n924, top_core_EC_n923, top_core_EC_n922,
         top_core_EC_n921, top_core_EC_n920, top_core_EC_n919,
         top_core_EC_n918, top_core_EC_n917, top_core_EC_n916,
         top_core_EC_n915, top_core_EC_n914, top_core_EC_n913,
         top_core_EC_n912, top_core_EC_n911, top_core_EC_n910,
         top_core_EC_n909, top_core_EC_n908, top_core_EC_n907,
         top_core_EC_n906, top_core_EC_n905, top_core_EC_n904,
         top_core_EC_n903, top_core_EC_n902, top_core_EC_n901,
         top_core_EC_n900, top_core_EC_n899, top_core_EC_n898,
         top_core_EC_n897, top_core_EC_n896, top_core_EC_n895,
         top_core_EC_n894, top_core_EC_n893, top_core_EC_n892,
         top_core_EC_n891, top_core_EC_n890, top_core_EC_n889,
         top_core_EC_n888, top_core_EC_n887, top_core_EC_n886,
         top_core_EC_n885, top_core_EC_n884, top_core_EC_n883,
         top_core_EC_n882, top_core_EC_n881, top_core_EC_n880,
         top_core_EC_n879, top_core_EC_n878, top_core_EC_n877,
         top_core_EC_n876, top_core_EC_n875, top_core_EC_n874,
         top_core_EC_n872, top_core_EC_n871, top_core_EC_n870,
         top_core_EC_n869, top_core_EC_n868, top_core_EC_n867,
         top_core_EC_n866, top_core_EC_n865, top_core_EC_n864,
         top_core_EC_n863, top_core_EC_n862, top_core_EC_n861,
         top_core_EC_n860, top_core_EC_n859, top_core_EC_n858,
         top_core_EC_n857, top_core_EC_n856, top_core_EC_n855,
         top_core_EC_n854, top_core_EC_n853, top_core_EC_n852,
         top_core_EC_n851, top_core_EC_n850, top_core_EC_n849,
         top_core_EC_n848, top_core_EC_n847, top_core_EC_n846,
         top_core_EC_n845, top_core_EC_n844, top_core_EC_n843,
         top_core_EC_n842, top_core_EC_n841, top_core_EC_n840,
         top_core_EC_n839, top_core_EC_n838, top_core_EC_n837,
         top_core_EC_n836, top_core_EC_n835, top_core_EC_n834,
         top_core_EC_n833, top_core_EC_n832, top_core_EC_n831,
         top_core_EC_n830, top_core_EC_n829, top_core_EC_n828,
         top_core_EC_n827, top_core_EC_n826, top_core_EC_n825,
         top_core_EC_n824, top_core_EC_n823, top_core_EC_n822,
         top_core_EC_n821, top_core_EC_n820, top_core_EC_n819,
         top_core_EC_n818, top_core_EC_n817, top_core_EC_n816,
         top_core_EC_n815, top_core_EC_n814, top_core_EC_n813,
         top_core_EC_n812, top_core_EC_n811, top_core_EC_n810,
         top_core_EC_n809, top_core_EC_n808, top_core_EC_n807,
         top_core_EC_n806, top_core_EC_n805, top_core_EC_n804,
         top_core_EC_n803, top_core_EC_n802, top_core_EC_n801,
         top_core_EC_n800, top_core_EC_n799, top_core_EC_n798,
         top_core_EC_n797, top_core_EC_n796, top_core_EC_n795,
         top_core_EC_n794, top_core_EC_n793, top_core_EC_n792,
         top_core_EC_n791, top_core_EC_n790, top_core_EC_n789,
         top_core_EC_n788, top_core_EC_n787, top_core_EC_n786,
         top_core_EC_n785, top_core_EC_n784, top_core_EC_n783,
         top_core_EC_n782, top_core_EC_n781, top_core_EC_n780,
         top_core_EC_n779, top_core_EC_n778, top_core_EC_n777,
         top_core_EC_n776, top_core_EC_n775, top_core_EC_n774,
         top_core_EC_n773, top_core_EC_n772, top_core_EC_n771,
         top_core_EC_n770, top_core_EC_n769, top_core_EC_n768,
         top_core_EC_n767, top_core_EC_n766, top_core_EC_n765,
         top_core_EC_n764, top_core_EC_n763, top_core_EC_n762,
         top_core_EC_n761, top_core_EC_n760, top_core_EC_n759,
         top_core_EC_n758, top_core_EC_n757, top_core_EC_n756,
         top_core_EC_n755, top_core_EC_n754, top_core_EC_n753,
         top_core_EC_n752, top_core_EC_n751, top_core_EC_n750,
         top_core_EC_n749, top_core_EC_n748, top_core_EC_n747,
         top_core_EC_n746, top_core_EC_n745, top_core_EC_n744,
         top_core_EC_n743, top_core_EC_n742, top_core_EC_n741,
         top_core_EC_n740, top_core_EC_n739, top_core_EC_n738,
         top_core_EC_n737, top_core_EC_n736, top_core_EC_n735,
         top_core_EC_n734, top_core_EC_n733, top_core_EC_n731,
         top_core_EC_n730, top_core_EC_n25, top_core_EC_N577, top_core_EC_N575,
         top_core_EC_mix_out_0_, top_core_EC_mix_out_1_,
         top_core_EC_mix_out_2_, top_core_EC_mix_out_3_,
         top_core_EC_mix_out_4_, top_core_EC_mix_out_5_,
         top_core_EC_mix_out_6_, top_core_EC_mix_out_7_,
         top_core_EC_mix_out_8_, top_core_EC_mix_out_9_,
         top_core_EC_mix_out_10_, top_core_EC_mix_out_11_,
         top_core_EC_mix_out_12_, top_core_EC_mix_out_13_,
         top_core_EC_mix_out_14_, top_core_EC_mix_out_15_,
         top_core_EC_mix_out_16_, top_core_EC_mix_out_17_,
         top_core_EC_mix_out_18_, top_core_EC_mix_out_19_,
         top_core_EC_mix_out_20_, top_core_EC_mix_out_21_,
         top_core_EC_mix_out_22_, top_core_EC_mix_out_23_,
         top_core_EC_mix_out_24_, top_core_EC_mix_out_25_,
         top_core_EC_mix_out_26_, top_core_EC_mix_out_27_,
         top_core_EC_mix_out_28_, top_core_EC_mix_out_29_,
         top_core_EC_mix_out_30_, top_core_EC_mix_out_31_,
         top_core_EC_mix_out_32_, top_core_EC_mix_out_33_,
         top_core_EC_mix_out_34_, top_core_EC_mix_out_35_,
         top_core_EC_mix_out_36_, top_core_EC_mix_out_37_,
         top_core_EC_mix_out_38_, top_core_EC_mix_out_39_,
         top_core_EC_mix_out_40_, top_core_EC_mix_out_41_,
         top_core_EC_mix_out_42_, top_core_EC_mix_out_43_,
         top_core_EC_mix_out_44_, top_core_EC_mix_out_45_,
         top_core_EC_mix_out_46_, top_core_EC_mix_out_47_,
         top_core_EC_mix_out_48_, top_core_EC_mix_out_49_,
         top_core_EC_mix_out_50_, top_core_EC_mix_out_51_,
         top_core_EC_mix_out_52_, top_core_EC_mix_out_53_,
         top_core_EC_mix_out_54_, top_core_EC_mix_out_55_,
         top_core_EC_mix_out_56_, top_core_EC_mix_out_57_,
         top_core_EC_mix_out_58_, top_core_EC_mix_out_59_,
         top_core_EC_mix_out_60_, top_core_EC_mix_out_61_,
         top_core_EC_mix_out_62_, top_core_EC_mix_out_63_,
         top_core_EC_mix_out_64_, top_core_EC_mix_out_65_,
         top_core_EC_mix_out_66_, top_core_EC_mix_out_67_,
         top_core_EC_mix_out_68_, top_core_EC_mix_out_69_,
         top_core_EC_mix_out_70_, top_core_EC_mix_out_71_,
         top_core_EC_mix_out_72_, top_core_EC_mix_out_73_,
         top_core_EC_mix_out_74_, top_core_EC_mix_out_75_,
         top_core_EC_mix_out_76_, top_core_EC_mix_out_77_,
         top_core_EC_mix_out_78_, top_core_EC_mix_out_79_,
         top_core_EC_mix_out_80_, top_core_EC_mix_out_81_,
         top_core_EC_mix_out_82_, top_core_EC_mix_out_83_,
         top_core_EC_mix_out_84_, top_core_EC_mix_out_85_,
         top_core_EC_mix_out_86_, top_core_EC_mix_out_87_,
         top_core_EC_mix_out_88_, top_core_EC_mix_out_89_,
         top_core_EC_mix_out_90_, top_core_EC_mix_out_91_,
         top_core_EC_mix_out_92_, top_core_EC_mix_out_93_,
         top_core_EC_mix_out_94_, top_core_EC_mix_out_95_,
         top_core_EC_mix_out_96_, top_core_EC_mix_out_97_,
         top_core_EC_mix_out_98_, top_core_EC_mix_out_99_,
         top_core_EC_mix_out_100_, top_core_EC_mix_out_101_,
         top_core_EC_mix_out_102_, top_core_EC_mix_out_103_,
         top_core_EC_mix_out_104_, top_core_EC_mix_out_105_,
         top_core_EC_mix_out_106_, top_core_EC_mix_out_107_,
         top_core_EC_mix_out_108_, top_core_EC_mix_out_109_,
         top_core_EC_mix_out_110_, top_core_EC_mix_out_111_,
         top_core_EC_mix_out_112_, top_core_EC_mix_out_113_,
         top_core_EC_mix_out_114_, top_core_EC_mix_out_115_,
         top_core_EC_mix_out_116_, top_core_EC_mix_out_117_,
         top_core_EC_mix_out_118_, top_core_EC_mix_out_119_,
         top_core_EC_mix_out_120_, top_core_EC_mix_out_121_,
         top_core_EC_mix_out_122_, top_core_EC_mix_out_123_,
         top_core_EC_mix_out_124_, top_core_EC_mix_out_125_,
         top_core_EC_mix_out_126_, top_core_EC_mix_out_127_,
         top_core_EC_round_result_r_0_, top_core_EC_round_result_r_1_,
         top_core_EC_round_result_r_2_, top_core_EC_round_result_r_3_,
         top_core_EC_round_result_r_4_, top_core_EC_round_result_r_5_,
         top_core_EC_round_result_r_6_, top_core_EC_round_result_r_7_,
         top_core_EC_round_result_r_8_, top_core_EC_round_result_r_9_,
         top_core_EC_round_result_r_10_, top_core_EC_round_result_r_11_,
         top_core_EC_round_result_r_12_, top_core_EC_round_result_r_13_,
         top_core_EC_round_result_r_14_, top_core_EC_round_result_r_15_,
         top_core_EC_round_result_r_16_, top_core_EC_round_result_r_17_,
         top_core_EC_round_result_r_18_, top_core_EC_round_result_r_19_,
         top_core_EC_round_result_r_20_, top_core_EC_round_result_r_21_,
         top_core_EC_round_result_r_22_, top_core_EC_round_result_r_23_,
         top_core_EC_round_result_r_24_, top_core_EC_round_result_r_25_,
         top_core_EC_round_result_r_26_, top_core_EC_round_result_r_27_,
         top_core_EC_round_result_r_28_, top_core_EC_round_result_r_29_,
         top_core_EC_round_result_r_30_, top_core_EC_round_result_r_31_,
         top_core_EC_round_result_r_32_, top_core_EC_round_result_r_33_,
         top_core_EC_round_result_r_34_, top_core_EC_round_result_r_35_,
         top_core_EC_round_result_r_36_, top_core_EC_round_result_r_37_,
         top_core_EC_round_result_r_38_, top_core_EC_round_result_r_39_,
         top_core_EC_round_result_r_40_, top_core_EC_round_result_r_41_,
         top_core_EC_round_result_r_42_, top_core_EC_round_result_r_43_,
         top_core_EC_round_result_r_44_, top_core_EC_round_result_r_45_,
         top_core_EC_round_result_r_46_, top_core_EC_round_result_r_47_,
         top_core_EC_round_result_r_48_, top_core_EC_round_result_r_49_,
         top_core_EC_round_result_r_50_, top_core_EC_round_result_r_51_,
         top_core_EC_round_result_r_52_, top_core_EC_round_result_r_53_,
         top_core_EC_round_result_r_54_, top_core_EC_round_result_r_55_,
         top_core_EC_round_result_r_56_, top_core_EC_round_result_r_57_,
         top_core_EC_round_result_r_58_, top_core_EC_round_result_r_59_,
         top_core_EC_round_result_r_60_, top_core_EC_round_result_r_61_,
         top_core_EC_round_result_r_62_, top_core_EC_round_result_r_63_,
         top_core_EC_round_result_r_64_, top_core_EC_round_result_r_65_,
         top_core_EC_round_result_r_66_, top_core_EC_round_result_r_67_,
         top_core_EC_round_result_r_68_, top_core_EC_round_result_r_69_,
         top_core_EC_round_result_r_70_, top_core_EC_round_result_r_71_,
         top_core_EC_round_result_r_72_, top_core_EC_round_result_r_73_,
         top_core_EC_round_result_r_74_, top_core_EC_round_result_r_75_,
         top_core_EC_round_result_r_76_, top_core_EC_round_result_r_77_,
         top_core_EC_round_result_r_78_, top_core_EC_round_result_r_79_,
         top_core_EC_round_result_r_80_, top_core_EC_round_result_r_81_,
         top_core_EC_round_result_r_82_, top_core_EC_round_result_r_83_,
         top_core_EC_round_result_r_84_, top_core_EC_round_result_r_85_,
         top_core_EC_round_result_r_86_, top_core_EC_round_result_r_87_,
         top_core_EC_round_result_r_88_, top_core_EC_round_result_r_89_,
         top_core_EC_round_result_r_90_, top_core_EC_round_result_r_91_,
         top_core_EC_round_result_r_92_, top_core_EC_round_result_r_93_,
         top_core_EC_round_result_r_94_, top_core_EC_round_result_r_95_,
         top_core_EC_round_result_r_96_, top_core_EC_round_result_r_97_,
         top_core_EC_round_result_r_98_, top_core_EC_round_result_r_99_,
         top_core_EC_round_result_r_100_, top_core_EC_round_result_r_101_,
         top_core_EC_round_result_r_102_, top_core_EC_round_result_r_103_,
         top_core_EC_round_result_r_104_, top_core_EC_round_result_r_105_,
         top_core_EC_round_result_r_106_, top_core_EC_round_result_r_107_,
         top_core_EC_round_result_r_108_, top_core_EC_round_result_r_109_,
         top_core_EC_round_result_r_110_, top_core_EC_round_result_r_111_,
         top_core_EC_round_result_r_112_, top_core_EC_round_result_r_113_,
         top_core_EC_round_result_r_114_, top_core_EC_round_result_r_115_,
         top_core_EC_round_result_r_116_, top_core_EC_round_result_r_117_,
         top_core_EC_round_result_r_118_, top_core_EC_round_result_r_119_,
         top_core_EC_round_result_r_120_, top_core_EC_round_result_r_121_,
         top_core_EC_round_result_r_122_, top_core_EC_round_result_r_123_,
         top_core_EC_round_result_r_124_, top_core_EC_round_result_r_125_,
         top_core_EC_round_result_r_126_, top_core_EC_round_result_r_127_,
         top_core_EC_round_result_0_, top_core_EC_round_result_1_,
         top_core_EC_round_result_2_, top_core_EC_round_result_3_,
         top_core_EC_round_result_4_, top_core_EC_round_result_5_,
         top_core_EC_round_result_6_, top_core_EC_round_result_7_,
         top_core_EC_round_result_8_, top_core_EC_round_result_9_,
         top_core_EC_round_result_10_, top_core_EC_round_result_11_,
         top_core_EC_round_result_12_, top_core_EC_round_result_13_,
         top_core_EC_round_result_14_, top_core_EC_round_result_15_,
         top_core_EC_round_result_16_, top_core_EC_round_result_17_,
         top_core_EC_round_result_18_, top_core_EC_round_result_19_,
         top_core_EC_round_result_20_, top_core_EC_round_result_21_,
         top_core_EC_round_result_22_, top_core_EC_round_result_23_,
         top_core_EC_round_result_24_, top_core_EC_round_result_25_,
         top_core_EC_round_result_26_, top_core_EC_round_result_27_,
         top_core_EC_round_result_28_, top_core_EC_round_result_29_,
         top_core_EC_round_result_30_, top_core_EC_round_result_31_,
         top_core_EC_round_result_32_, top_core_EC_round_result_33_,
         top_core_EC_round_result_34_, top_core_EC_round_result_35_,
         top_core_EC_round_result_36_, top_core_EC_round_result_37_,
         top_core_EC_round_result_38_, top_core_EC_round_result_39_,
         top_core_EC_round_result_40_, top_core_EC_round_result_41_,
         top_core_EC_round_result_42_, top_core_EC_round_result_43_,
         top_core_EC_round_result_44_, top_core_EC_round_result_45_,
         top_core_EC_round_result_46_, top_core_EC_round_result_47_,
         top_core_EC_round_result_48_, top_core_EC_round_result_49_,
         top_core_EC_round_result_50_, top_core_EC_round_result_51_,
         top_core_EC_round_result_52_, top_core_EC_round_result_53_,
         top_core_EC_round_result_54_, top_core_EC_round_result_55_,
         top_core_EC_round_result_56_, top_core_EC_round_result_57_,
         top_core_EC_round_result_58_, top_core_EC_round_result_59_,
         top_core_EC_round_result_60_, top_core_EC_round_result_61_,
         top_core_EC_round_result_62_, top_core_EC_round_result_63_,
         top_core_EC_round_result_64_, top_core_EC_round_result_65_,
         top_core_EC_round_result_66_, top_core_EC_round_result_67_,
         top_core_EC_round_result_68_, top_core_EC_round_result_69_,
         top_core_EC_round_result_70_, top_core_EC_round_result_71_,
         top_core_EC_round_result_72_, top_core_EC_round_result_73_,
         top_core_EC_round_result_74_, top_core_EC_round_result_75_,
         top_core_EC_round_result_76_, top_core_EC_round_result_77_,
         top_core_EC_round_result_78_, top_core_EC_round_result_79_,
         top_core_EC_round_result_80_, top_core_EC_round_result_81_,
         top_core_EC_round_result_82_, top_core_EC_round_result_83_,
         top_core_EC_round_result_84_, top_core_EC_round_result_85_,
         top_core_EC_round_result_86_, top_core_EC_round_result_87_,
         top_core_EC_round_result_88_, top_core_EC_round_result_89_,
         top_core_EC_round_result_90_, top_core_EC_round_result_91_,
         top_core_EC_round_result_92_, top_core_EC_round_result_93_,
         top_core_EC_round_result_94_, top_core_EC_round_result_95_,
         top_core_EC_round_result_96_, top_core_EC_round_result_97_,
         top_core_EC_round_result_98_, top_core_EC_round_result_99_,
         top_core_EC_round_result_100_, top_core_EC_round_result_101_,
         top_core_EC_round_result_102_, top_core_EC_round_result_103_,
         top_core_EC_round_result_104_, top_core_EC_round_result_105_,
         top_core_EC_round_result_106_, top_core_EC_round_result_107_,
         top_core_EC_round_result_108_, top_core_EC_round_result_109_,
         top_core_EC_round_result_110_, top_core_EC_round_result_111_,
         top_core_EC_round_result_112_, top_core_EC_round_result_113_,
         top_core_EC_round_result_114_, top_core_EC_round_result_115_,
         top_core_EC_round_result_116_, top_core_EC_round_result_117_,
         top_core_EC_round_result_118_, top_core_EC_round_result_119_,
         top_core_EC_round_result_120_, top_core_EC_round_result_121_,
         top_core_EC_round_result_122_, top_core_EC_round_result_123_,
         top_core_EC_round_result_124_, top_core_EC_round_result_125_,
         top_core_EC_round_result_126_, top_core_EC_round_result_127_,
         top_core_EC_N276, top_core_EC_N275, top_core_EC_N274,
         top_core_EC_N273, top_core_EC_N272, top_core_EC_N271,
         top_core_EC_N270, top_core_EC_N269, top_core_EC_N268,
         top_core_EC_N267, top_core_EC_N266, top_core_EC_N265,
         top_core_EC_N264, top_core_EC_N263, top_core_EC_N262,
         top_core_EC_N261, top_core_EC_N260, top_core_EC_N259,
         top_core_EC_N258, top_core_EC_N257, top_core_EC_N256,
         top_core_EC_N255, top_core_EC_N254, top_core_EC_N253,
         top_core_EC_N252, top_core_EC_N251, top_core_EC_N250,
         top_core_EC_N249, top_core_EC_N248, top_core_EC_N247,
         top_core_EC_N246, top_core_EC_N245, top_core_EC_N244,
         top_core_EC_N243, top_core_EC_N242, top_core_EC_N241,
         top_core_EC_N240, top_core_EC_N239, top_core_EC_N238,
         top_core_EC_N237, top_core_EC_N236, top_core_EC_N235,
         top_core_EC_N234, top_core_EC_N233, top_core_EC_N232,
         top_core_EC_N231, top_core_EC_N230, top_core_EC_N229,
         top_core_EC_N228, top_core_EC_N227, top_core_EC_N226,
         top_core_EC_N225, top_core_EC_N224, top_core_EC_N223,
         top_core_EC_N222, top_core_EC_N221, top_core_EC_N220,
         top_core_EC_N219, top_core_EC_N218, top_core_EC_N217,
         top_core_EC_N216, top_core_EC_N215, top_core_EC_N214,
         top_core_EC_N213, top_core_EC_N212, top_core_EC_N211,
         top_core_EC_N210, top_core_EC_N209, top_core_EC_N208,
         top_core_EC_N207, top_core_EC_N206, top_core_EC_N205,
         top_core_EC_N204, top_core_EC_N203, top_core_EC_N202,
         top_core_EC_N201, top_core_EC_N200, top_core_EC_N199,
         top_core_EC_N198, top_core_EC_N197, top_core_EC_N196,
         top_core_EC_N195, top_core_EC_N194, top_core_EC_N193,
         top_core_EC_N192, top_core_EC_N191, top_core_EC_N190,
         top_core_EC_N189, top_core_EC_N188, top_core_EC_N187,
         top_core_EC_N186, top_core_EC_N185, top_core_EC_N184,
         top_core_EC_N183, top_core_EC_N182, top_core_EC_N181,
         top_core_EC_N180, top_core_EC_N179, top_core_EC_N178,
         top_core_EC_N177, top_core_EC_N176, top_core_EC_N175,
         top_core_EC_N174, top_core_EC_N173, top_core_EC_N172,
         top_core_EC_N171, top_core_EC_N170, top_core_EC_N169,
         top_core_EC_N168, top_core_EC_N167, top_core_EC_N166,
         top_core_EC_N165, top_core_EC_N164, top_core_EC_N163,
         top_core_EC_N162, top_core_EC_N161, top_core_EC_N160,
         top_core_EC_N159, top_core_EC_N158, top_core_EC_N157,
         top_core_EC_N156, top_core_EC_N155, top_core_EC_N154,
         top_core_EC_N153, top_core_EC_N152, top_core_EC_N151,
         top_core_EC_N150, top_core_EC_N149, top_core_EC_add_out_r_0_,
         top_core_EC_add_out_r_1_, top_core_EC_add_out_r_2_,
         top_core_EC_add_out_r_3_, top_core_EC_add_out_r_4_,
         top_core_EC_add_out_r_5_, top_core_EC_add_out_r_6_,
         top_core_EC_add_out_r_7_, top_core_EC_add_out_r_8_,
         top_core_EC_add_out_r_9_, top_core_EC_add_out_r_10_,
         top_core_EC_add_out_r_11_, top_core_EC_add_out_r_12_,
         top_core_EC_add_out_r_13_, top_core_EC_add_out_r_14_,
         top_core_EC_add_out_r_15_, top_core_EC_add_out_r_16_,
         top_core_EC_add_out_r_17_, top_core_EC_add_out_r_18_,
         top_core_EC_add_out_r_19_, top_core_EC_add_out_r_20_,
         top_core_EC_add_out_r_21_, top_core_EC_add_out_r_22_,
         top_core_EC_add_out_r_23_, top_core_EC_add_out_r_24_,
         top_core_EC_add_out_r_25_, top_core_EC_add_out_r_26_,
         top_core_EC_add_out_r_27_, top_core_EC_add_out_r_28_,
         top_core_EC_add_out_r_29_, top_core_EC_add_out_r_30_,
         top_core_EC_add_out_r_31_, top_core_EC_add_out_r_32_,
         top_core_EC_add_out_r_33_, top_core_EC_add_out_r_34_,
         top_core_EC_add_out_r_35_, top_core_EC_add_out_r_36_,
         top_core_EC_add_out_r_37_, top_core_EC_add_out_r_38_,
         top_core_EC_add_out_r_39_, top_core_EC_add_out_r_40_,
         top_core_EC_add_out_r_41_, top_core_EC_add_out_r_42_,
         top_core_EC_add_out_r_43_, top_core_EC_add_out_r_44_,
         top_core_EC_add_out_r_45_, top_core_EC_add_out_r_46_,
         top_core_EC_add_out_r_47_, top_core_EC_add_out_r_48_,
         top_core_EC_add_out_r_49_, top_core_EC_add_out_r_50_,
         top_core_EC_add_out_r_51_, top_core_EC_add_out_r_52_,
         top_core_EC_add_out_r_53_, top_core_EC_add_out_r_54_,
         top_core_EC_add_out_r_55_, top_core_EC_add_out_r_56_,
         top_core_EC_add_out_r_57_, top_core_EC_rounds_2_,
         top_core_EC_rounds_3_, top_core_EC_operation, top_core_KE_n5707,
         top_core_KE_n5706, top_core_KE_n5705, top_core_KE_n5704,
         top_core_KE_n5703, top_core_KE_n5702, top_core_KE_n5701,
         top_core_KE_n5700, top_core_KE_n5699, top_core_KE_n5698,
         top_core_KE_n5697, top_core_KE_n5696, top_core_KE_n5695,
         top_core_KE_n5694, top_core_KE_n5693, top_core_KE_n5692,
         top_core_KE_n5691, top_core_KE_n5690, top_core_KE_n5689,
         top_core_KE_n5688, top_core_KE_n5687, top_core_KE_n5686,
         top_core_KE_n5685, top_core_KE_n5684, top_core_KE_n5683,
         top_core_KE_n5682, top_core_KE_n5681, top_core_KE_n5680,
         top_core_KE_n5679, top_core_KE_n5678, top_core_KE_n5677,
         top_core_KE_n5676, top_core_KE_n5675, top_core_KE_n5674,
         top_core_KE_n5673, top_core_KE_n5672, top_core_KE_n5671,
         top_core_KE_n5670, top_core_KE_n5669, top_core_KE_n5668,
         top_core_KE_n5667, top_core_KE_n5666, top_core_KE_n5665,
         top_core_KE_n5664, top_core_KE_n5663, top_core_KE_n5662,
         top_core_KE_n5661, top_core_KE_n5660, top_core_KE_n5659,
         top_core_KE_n5658, top_core_KE_n5657, top_core_KE_n5656,
         top_core_KE_n5655, top_core_KE_n5654, top_core_KE_n5653,
         top_core_KE_n5652, top_core_KE_n5651, top_core_KE_n5650,
         top_core_KE_n5649, top_core_KE_n5648, top_core_KE_n5647,
         top_core_KE_n5646, top_core_KE_n5645, top_core_KE_n5644,
         top_core_KE_n5643, top_core_KE_n5642, top_core_KE_n5641,
         top_core_KE_n5640, top_core_KE_n5639, top_core_KE_n5638,
         top_core_KE_n5637, top_core_KE_n5636, top_core_KE_n5635,
         top_core_KE_n5634, top_core_KE_n5633, top_core_KE_n5632,
         top_core_KE_n5631, top_core_KE_n5630, top_core_KE_n5629,
         top_core_KE_n5628, top_core_KE_n5627, top_core_KE_n5626,
         top_core_KE_n5625, top_core_KE_n5624, top_core_KE_n5623,
         top_core_KE_n5622, top_core_KE_n5621, top_core_KE_n5620,
         top_core_KE_n5619, top_core_KE_n5618, top_core_KE_n5617,
         top_core_KE_n5616, top_core_KE_n5615, top_core_KE_n5614,
         top_core_KE_n5613, top_core_KE_n5612, top_core_KE_n5611,
         top_core_KE_n5610, top_core_KE_n5609, top_core_KE_n5608,
         top_core_KE_n5607, top_core_KE_n5606, top_core_KE_n5605,
         top_core_KE_n5604, top_core_KE_n5603, top_core_KE_n5602,
         top_core_KE_n5601, top_core_KE_n5600, top_core_KE_n5599,
         top_core_KE_n5598, top_core_KE_n5597, top_core_KE_n5596,
         top_core_KE_n5595, top_core_KE_n5594, top_core_KE_n5593,
         top_core_KE_n5592, top_core_KE_n5591, top_core_KE_n5590,
         top_core_KE_n5589, top_core_KE_n5588, top_core_KE_n5587,
         top_core_KE_n5586, top_core_KE_n5585, top_core_KE_n5584,
         top_core_KE_n5583, top_core_KE_n5582, top_core_KE_n5581,
         top_core_KE_n5580, top_core_KE_n5579, top_core_KE_n5578,
         top_core_KE_n5577, top_core_KE_n5576, top_core_KE_n5575,
         top_core_KE_n5574, top_core_KE_n5573, top_core_KE_n5572,
         top_core_KE_n5571, top_core_KE_n5570, top_core_KE_n5569,
         top_core_KE_n5568, top_core_KE_n5567, top_core_KE_n5566,
         top_core_KE_n5565, top_core_KE_n5564, top_core_KE_n5563,
         top_core_KE_n5562, top_core_KE_n5561, top_core_KE_n5560,
         top_core_KE_n5559, top_core_KE_n5558, top_core_KE_n5557,
         top_core_KE_n5556, top_core_KE_n5555, top_core_KE_n5554,
         top_core_KE_n5553, top_core_KE_n5552, top_core_KE_n5551,
         top_core_KE_n5550, top_core_KE_n5549, top_core_KE_n5548,
         top_core_KE_n5547, top_core_KE_n5546, top_core_KE_n5545,
         top_core_KE_n5544, top_core_KE_n5543, top_core_KE_n5542,
         top_core_KE_n5541, top_core_KE_n5540, top_core_KE_n5539,
         top_core_KE_n5538, top_core_KE_n5537, top_core_KE_n5536,
         top_core_KE_n5535, top_core_KE_n5534, top_core_KE_n5533,
         top_core_KE_n5532, top_core_KE_n5531, top_core_KE_n5530,
         top_core_KE_n5529, top_core_KE_n5528, top_core_KE_n5527,
         top_core_KE_n5526, top_core_KE_n5525, top_core_KE_n5524,
         top_core_KE_n5523, top_core_KE_n5522, top_core_KE_n5521,
         top_core_KE_n5520, top_core_KE_n5519, top_core_KE_n5518,
         top_core_KE_n5517, top_core_KE_n5516, top_core_KE_n5515,
         top_core_KE_n5514, top_core_KE_n5513, top_core_KE_n5512,
         top_core_KE_n5511, top_core_KE_n5510, top_core_KE_n5509,
         top_core_KE_n5508, top_core_KE_n5507, top_core_KE_n5506,
         top_core_KE_n5505, top_core_KE_n5504, top_core_KE_n5503,
         top_core_KE_n5502, top_core_KE_n5501, top_core_KE_n5500,
         top_core_KE_n5499, top_core_KE_n5498, top_core_KE_n5497,
         top_core_KE_n5496, top_core_KE_n5495, top_core_KE_n5494,
         top_core_KE_n5493, top_core_KE_n5492, top_core_KE_n5491,
         top_core_KE_n5490, top_core_KE_n5489, top_core_KE_n5488,
         top_core_KE_n5487, top_core_KE_n5486, top_core_KE_n5485,
         top_core_KE_n5484, top_core_KE_n5483, top_core_KE_n5482,
         top_core_KE_n5481, top_core_KE_n5480, top_core_KE_n5479,
         top_core_KE_n5478, top_core_KE_n5477, top_core_KE_n5476,
         top_core_KE_n5475, top_core_KE_n5474, top_core_KE_n5473,
         top_core_KE_n5472, top_core_KE_n5471, top_core_KE_n5470,
         top_core_KE_n5469, top_core_KE_n5468, top_core_KE_n5467,
         top_core_KE_n5466, top_core_KE_n5465, top_core_KE_n5464,
         top_core_KE_n5463, top_core_KE_n5462, top_core_KE_n5461,
         top_core_KE_n5460, top_core_KE_n5459, top_core_KE_n5458,
         top_core_KE_n5457, top_core_KE_n5456, top_core_KE_n5455,
         top_core_KE_n5454, top_core_KE_n5453, top_core_KE_n5452,
         top_core_KE_n5451, top_core_KE_n5450, top_core_KE_n5449,
         top_core_KE_n5448, top_core_KE_n5447, top_core_KE_n5446,
         top_core_KE_n5445, top_core_KE_n5444, top_core_KE_n5443,
         top_core_KE_n5442, top_core_KE_n5441, top_core_KE_n5440,
         top_core_KE_n5439, top_core_KE_n5438, top_core_KE_n5437,
         top_core_KE_n5436, top_core_KE_n5435, top_core_KE_n5434,
         top_core_KE_n5433, top_core_KE_n5432, top_core_KE_n5431,
         top_core_KE_n5430, top_core_KE_n5429, top_core_KE_n5428,
         top_core_KE_n5427, top_core_KE_n5426, top_core_KE_n5425,
         top_core_KE_n5424, top_core_KE_n5423, top_core_KE_n5422,
         top_core_KE_n5421, top_core_KE_n5420, top_core_KE_n5419,
         top_core_KE_n5418, top_core_KE_n5417, top_core_KE_n5416,
         top_core_KE_n5415, top_core_KE_n5414, top_core_KE_n5413,
         top_core_KE_n5412, top_core_KE_n5411, top_core_KE_n5410,
         top_core_KE_n5409, top_core_KE_n5408, top_core_KE_n5407,
         top_core_KE_n5406, top_core_KE_n5405, top_core_KE_n5404,
         top_core_KE_n5403, top_core_KE_n5402, top_core_KE_n5401,
         top_core_KE_n5400, top_core_KE_n5399, top_core_KE_n5398,
         top_core_KE_n5397, top_core_KE_n5396, top_core_KE_n5395,
         top_core_KE_n5394, top_core_KE_n5393, top_core_KE_n5392,
         top_core_KE_n5391, top_core_KE_n5390, top_core_KE_n5389,
         top_core_KE_n5388, top_core_KE_n5387, top_core_KE_n5386,
         top_core_KE_n5385, top_core_KE_n5384, top_core_KE_n5383,
         top_core_KE_n5382, top_core_KE_n5381, top_core_KE_n5380,
         top_core_KE_n5379, top_core_KE_n5378, top_core_KE_n5377,
         top_core_KE_n5376, top_core_KE_n5375, top_core_KE_n5374,
         top_core_KE_n5373, top_core_KE_n5372, top_core_KE_n5371,
         top_core_KE_n5370, top_core_KE_n5369, top_core_KE_n5368,
         top_core_KE_n5367, top_core_KE_n5366, top_core_KE_n5365,
         top_core_KE_n5364, top_core_KE_n5363, top_core_KE_n5362,
         top_core_KE_n5361, top_core_KE_n5360, top_core_KE_n5359,
         top_core_KE_n5358, top_core_KE_n5357, top_core_KE_n5356,
         top_core_KE_n5355, top_core_KE_n5354, top_core_KE_n5353,
         top_core_KE_n5352, top_core_KE_n5351, top_core_KE_n5350,
         top_core_KE_n5349, top_core_KE_n5348, top_core_KE_n5347,
         top_core_KE_n5346, top_core_KE_n5345, top_core_KE_n5344,
         top_core_KE_n5343, top_core_KE_n5342, top_core_KE_n5341,
         top_core_KE_n5340, top_core_KE_n5339, top_core_KE_n5338,
         top_core_KE_n5337, top_core_KE_n5336, top_core_KE_n5335,
         top_core_KE_n5334, top_core_KE_n5333, top_core_KE_n5332,
         top_core_KE_n5331, top_core_KE_n5330, top_core_KE_n5329,
         top_core_KE_n5328, top_core_KE_n5327, top_core_KE_n5326,
         top_core_KE_n5325, top_core_KE_n5324, top_core_KE_n5323,
         top_core_KE_n5322, top_core_KE_n5321, top_core_KE_n5320,
         top_core_KE_n5319, top_core_KE_n5318, top_core_KE_n5317,
         top_core_KE_n5316, top_core_KE_n5315, top_core_KE_n5314,
         top_core_KE_n5313, top_core_KE_n5312, top_core_KE_n5311,
         top_core_KE_n5310, top_core_KE_n5309, top_core_KE_n5308,
         top_core_KE_n5307, top_core_KE_n5306, top_core_KE_n5305,
         top_core_KE_n5304, top_core_KE_n5303, top_core_KE_n5302,
         top_core_KE_n5301, top_core_KE_n5300, top_core_KE_n5299,
         top_core_KE_n5298, top_core_KE_n5297, top_core_KE_n5296,
         top_core_KE_n5295, top_core_KE_n5294, top_core_KE_n5293,
         top_core_KE_n5292, top_core_KE_n5291, top_core_KE_n5290,
         top_core_KE_n5289, top_core_KE_n5288, top_core_KE_n5287,
         top_core_KE_n5286, top_core_KE_n5285, top_core_KE_n5284,
         top_core_KE_n5283, top_core_KE_n5282, top_core_KE_n5281,
         top_core_KE_n5280, top_core_KE_n5279, top_core_KE_n5278,
         top_core_KE_n5277, top_core_KE_n5276, top_core_KE_n5275,
         top_core_KE_n5274, top_core_KE_n5273, top_core_KE_n5272,
         top_core_KE_n5271, top_core_KE_n5270, top_core_KE_n5269,
         top_core_KE_n5268, top_core_KE_n5267, top_core_KE_n5266,
         top_core_KE_n5265, top_core_KE_n5264, top_core_KE_n5263,
         top_core_KE_n5262, top_core_KE_n5261, top_core_KE_n5260,
         top_core_KE_n5259, top_core_KE_n5258, top_core_KE_n5257,
         top_core_KE_n5256, top_core_KE_n5255, top_core_KE_n5254,
         top_core_KE_n5253, top_core_KE_n5252, top_core_KE_n5251,
         top_core_KE_n5250, top_core_KE_n5249, top_core_KE_n5248,
         top_core_KE_n5247, top_core_KE_n5246, top_core_KE_n5245,
         top_core_KE_n5244, top_core_KE_n5243, top_core_KE_n5242,
         top_core_KE_n5241, top_core_KE_n5240, top_core_KE_n5239,
         top_core_KE_n5238, top_core_KE_n5237, top_core_KE_n5236,
         top_core_KE_n5235, top_core_KE_n5234, top_core_KE_n5233,
         top_core_KE_n5232, top_core_KE_n5231, top_core_KE_n5230,
         top_core_KE_n5229, top_core_KE_n5228, top_core_KE_n5227,
         top_core_KE_n5226, top_core_KE_n5225, top_core_KE_n5224,
         top_core_KE_n5223, top_core_KE_n5222, top_core_KE_n5221,
         top_core_KE_n5220, top_core_KE_n5219, top_core_KE_n5218,
         top_core_KE_n5217, top_core_KE_n5216, top_core_KE_n5215,
         top_core_KE_n5214, top_core_KE_n5213, top_core_KE_n5212,
         top_core_KE_n5211, top_core_KE_n5210, top_core_KE_n5209,
         top_core_KE_n5208, top_core_KE_n5207, top_core_KE_n5206,
         top_core_KE_n5205, top_core_KE_n5204, top_core_KE_n5203,
         top_core_KE_n5202, top_core_KE_n5201, top_core_KE_n5200,
         top_core_KE_n5199, top_core_KE_n5198, top_core_KE_n5197,
         top_core_KE_n5196, top_core_KE_n5195, top_core_KE_n5194,
         top_core_KE_n5193, top_core_KE_n5192, top_core_KE_n5191,
         top_core_KE_n5190, top_core_KE_n5189, top_core_KE_n5188,
         top_core_KE_n5187, top_core_KE_n5186, top_core_KE_n5185,
         top_core_KE_n5184, top_core_KE_n5183, top_core_KE_n5182,
         top_core_KE_n5181, top_core_KE_n5180, top_core_KE_n5179,
         top_core_KE_n5178, top_core_KE_n5177, top_core_KE_n5176,
         top_core_KE_n5175, top_core_KE_n5174, top_core_KE_n5173,
         top_core_KE_n5172, top_core_KE_n5171, top_core_KE_n5170,
         top_core_KE_n5169, top_core_KE_n5168, top_core_KE_n5167,
         top_core_KE_n5166, top_core_KE_n5165, top_core_KE_n5164,
         top_core_KE_n5163, top_core_KE_n5162, top_core_KE_n5161,
         top_core_KE_n5160, top_core_KE_n5159, top_core_KE_n5158,
         top_core_KE_n5157, top_core_KE_n5156, top_core_KE_n5155,
         top_core_KE_n5154, top_core_KE_n5153, top_core_KE_n5152,
         top_core_KE_n5151, top_core_KE_n5150, top_core_KE_n5149,
         top_core_KE_n5148, top_core_KE_n5147, top_core_KE_n5146,
         top_core_KE_n5145, top_core_KE_n5144, top_core_KE_n5143,
         top_core_KE_n5142, top_core_KE_n5141, top_core_KE_n5140,
         top_core_KE_n5139, top_core_KE_n5138, top_core_KE_n5137,
         top_core_KE_n5136, top_core_KE_n5135, top_core_KE_n5134,
         top_core_KE_n5133, top_core_KE_n5132, top_core_KE_n5131,
         top_core_KE_n5130, top_core_KE_n5129, top_core_KE_n5128,
         top_core_KE_n5127, top_core_KE_n5126, top_core_KE_n5125,
         top_core_KE_n5124, top_core_KE_n5123, top_core_KE_n5122,
         top_core_KE_n5121, top_core_KE_n5120, top_core_KE_n5119,
         top_core_KE_n5118, top_core_KE_n5117, top_core_KE_n5116,
         top_core_KE_n5115, top_core_KE_n5114, top_core_KE_n5113,
         top_core_KE_n5112, top_core_KE_n5111, top_core_KE_n5110,
         top_core_KE_n5109, top_core_KE_n5108, top_core_KE_n5107,
         top_core_KE_n5106, top_core_KE_n5105, top_core_KE_n5104,
         top_core_KE_n5103, top_core_KE_n5102, top_core_KE_n5101,
         top_core_KE_n5100, top_core_KE_n5099, top_core_KE_n5098,
         top_core_KE_n5097, top_core_KE_n5096, top_core_KE_n5095,
         top_core_KE_n5094, top_core_KE_n5093, top_core_KE_n5092,
         top_core_KE_n5091, top_core_KE_n5090, top_core_KE_n5089,
         top_core_KE_n5088, top_core_KE_n5087, top_core_KE_n5086,
         top_core_KE_n5085, top_core_KE_n5084, top_core_KE_n5083,
         top_core_KE_n5082, top_core_KE_n5081, top_core_KE_n5080,
         top_core_KE_n5079, top_core_KE_n5078, top_core_KE_n5077,
         top_core_KE_n5076, top_core_KE_n5075, top_core_KE_n5074,
         top_core_KE_n5073, top_core_KE_n5072, top_core_KE_n5071,
         top_core_KE_n5070, top_core_KE_n5069, top_core_KE_n5068,
         top_core_KE_n5067, top_core_KE_n5066, top_core_KE_n5065,
         top_core_KE_n5064, top_core_KE_n5063, top_core_KE_n5062,
         top_core_KE_n5061, top_core_KE_n5060, top_core_KE_n5059,
         top_core_KE_n5058, top_core_KE_n5057, top_core_KE_n5056,
         top_core_KE_n5055, top_core_KE_n5054, top_core_KE_n5053,
         top_core_KE_n5052, top_core_KE_n5051, top_core_KE_n5050,
         top_core_KE_n5049, top_core_KE_n5048, top_core_KE_n5047,
         top_core_KE_n5046, top_core_KE_n5045, top_core_KE_n5044,
         top_core_KE_n5043, top_core_KE_n5042, top_core_KE_n5041,
         top_core_KE_n5040, top_core_KE_n5039, top_core_KE_n5038,
         top_core_KE_n5037, top_core_KE_n5036, top_core_KE_n5035,
         top_core_KE_n5034, top_core_KE_n5033, top_core_KE_n5032,
         top_core_KE_n5031, top_core_KE_n5030, top_core_KE_n5029,
         top_core_KE_n5028, top_core_KE_n5027, top_core_KE_n5026,
         top_core_KE_n5025, top_core_KE_n5024, top_core_KE_n5023,
         top_core_KE_n5022, top_core_KE_n5021, top_core_KE_n5020,
         top_core_KE_n5019, top_core_KE_n5018, top_core_KE_n5017,
         top_core_KE_n5016, top_core_KE_n5015, top_core_KE_n5014,
         top_core_KE_n5013, top_core_KE_n5012, top_core_KE_n5011,
         top_core_KE_n5010, top_core_KE_n5009, top_core_KE_n5008,
         top_core_KE_n5007, top_core_KE_n5006, top_core_KE_n5005,
         top_core_KE_n5004, top_core_KE_n5003, top_core_KE_n5002,
         top_core_KE_n5001, top_core_KE_n5000, top_core_KE_n4999,
         top_core_KE_n4998, top_core_KE_n4997, top_core_KE_n4996,
         top_core_KE_n4995, top_core_KE_n4994, top_core_KE_n4993,
         top_core_KE_n4992, top_core_KE_n4991, top_core_KE_n4990,
         top_core_KE_n4989, top_core_KE_n4988, top_core_KE_n4987,
         top_core_KE_n4986, top_core_KE_n4985, top_core_KE_n4984,
         top_core_KE_n4983, top_core_KE_n4982, top_core_KE_n4981,
         top_core_KE_n4980, top_core_KE_n4979, top_core_KE_n4978,
         top_core_KE_n4977, top_core_KE_n4976, top_core_KE_n4975,
         top_core_KE_n4974, top_core_KE_n4973, top_core_KE_n4972,
         top_core_KE_n4971, top_core_KE_n4970, top_core_KE_n4969,
         top_core_KE_n4968, top_core_KE_n4967, top_core_KE_n4966,
         top_core_KE_n4965, top_core_KE_n4964, top_core_KE_n4963,
         top_core_KE_n4962, top_core_KE_n4961, top_core_KE_n4960,
         top_core_KE_n4959, top_core_KE_n4958, top_core_KE_n4957,
         top_core_KE_n4956, top_core_KE_n4955, top_core_KE_n4954,
         top_core_KE_n4953, top_core_KE_n4952, top_core_KE_n4951,
         top_core_KE_n4950, top_core_KE_n4949, top_core_KE_n4948,
         top_core_KE_n4947, top_core_KE_n4946, top_core_KE_n4945,
         top_core_KE_n4944, top_core_KE_n4943, top_core_KE_n4942,
         top_core_KE_n4941, top_core_KE_n4940, top_core_KE_n4939,
         top_core_KE_n4938, top_core_KE_n4937, top_core_KE_n4936,
         top_core_KE_n4935, top_core_KE_n4934, top_core_KE_n4933,
         top_core_KE_n4932, top_core_KE_n4931, top_core_KE_n4930,
         top_core_KE_n4929, top_core_KE_n4928, top_core_KE_n4927,
         top_core_KE_n4926, top_core_KE_n4925, top_core_KE_n4924,
         top_core_KE_n4923, top_core_KE_n4922, top_core_KE_n4921,
         top_core_KE_n4920, top_core_KE_n4919, top_core_KE_n4918,
         top_core_KE_n4917, top_core_KE_n4916, top_core_KE_n4915,
         top_core_KE_n4914, top_core_KE_n4913, top_core_KE_n4912,
         top_core_KE_n4911, top_core_KE_n4910, top_core_KE_n4909,
         top_core_KE_n4908, top_core_KE_n4907, top_core_KE_n4906,
         top_core_KE_n4905, top_core_KE_n4904, top_core_KE_n4903,
         top_core_KE_n4902, top_core_KE_n4901, top_core_KE_n4900,
         top_core_KE_n4899, top_core_KE_n4898, top_core_KE_n4897,
         top_core_KE_n4896, top_core_KE_n4895, top_core_KE_n4894,
         top_core_KE_n4893, top_core_KE_n4892, top_core_KE_n4891,
         top_core_KE_n4890, top_core_KE_n4889, top_core_KE_n4888,
         top_core_KE_n4887, top_core_KE_n4886, top_core_KE_n4885,
         top_core_KE_n4884, top_core_KE_n4883, top_core_KE_n4882,
         top_core_KE_n4881, top_core_KE_n4880, top_core_KE_n4879,
         top_core_KE_n4878, top_core_KE_n4877, top_core_KE_n4876,
         top_core_KE_n4875, top_core_KE_n4874, top_core_KE_n4873,
         top_core_KE_n4872, top_core_KE_n4871, top_core_KE_n4870,
         top_core_KE_n4869, top_core_KE_n4868, top_core_KE_n4867,
         top_core_KE_n4866, top_core_KE_n4865, top_core_KE_n4864,
         top_core_KE_n4863, top_core_KE_n4862, top_core_KE_n4861,
         top_core_KE_n4860, top_core_KE_n4859, top_core_KE_n4858,
         top_core_KE_n4857, top_core_KE_n4856, top_core_KE_n4855,
         top_core_KE_n4854, top_core_KE_n4853, top_core_KE_n4852,
         top_core_KE_n4851, top_core_KE_n4850, top_core_KE_n4849,
         top_core_KE_n4848, top_core_KE_n4847, top_core_KE_n4846,
         top_core_KE_n4845, top_core_KE_n4844, top_core_KE_n4843,
         top_core_KE_n4842, top_core_KE_n4841, top_core_KE_n4840,
         top_core_KE_n4839, top_core_KE_n4838, top_core_KE_n4837,
         top_core_KE_n4836, top_core_KE_n4835, top_core_KE_n4834,
         top_core_KE_n4833, top_core_KE_n4832, top_core_KE_n4831,
         top_core_KE_n4830, top_core_KE_n4829, top_core_KE_n4828,
         top_core_KE_n4827, top_core_KE_n4826, top_core_KE_n4825,
         top_core_KE_n4824, top_core_KE_n4823, top_core_KE_n4822,
         top_core_KE_n4821, top_core_KE_n4820, top_core_KE_n4819,
         top_core_KE_n4818, top_core_KE_n4817, top_core_KE_n4816,
         top_core_KE_n4815, top_core_KE_n4814, top_core_KE_n4813,
         top_core_KE_n4812, top_core_KE_n4811, top_core_KE_n4810,
         top_core_KE_n4809, top_core_KE_n4808, top_core_KE_n4807,
         top_core_KE_n4806, top_core_KE_n4805, top_core_KE_n4804,
         top_core_KE_n4803, top_core_KE_n4802, top_core_KE_n4801,
         top_core_KE_n4800, top_core_KE_n4799, top_core_KE_n4798,
         top_core_KE_n4797, top_core_KE_n4796, top_core_KE_n4795,
         top_core_KE_n4794, top_core_KE_n4793, top_core_KE_n4792,
         top_core_KE_n4791, top_core_KE_n4790, top_core_KE_n4789,
         top_core_KE_n4788, top_core_KE_n4787, top_core_KE_n4786,
         top_core_KE_n4785, top_core_KE_n4784, top_core_KE_n4783,
         top_core_KE_n4782, top_core_KE_n4781, top_core_KE_n4780,
         top_core_KE_n4779, top_core_KE_n4778, top_core_KE_n4777,
         top_core_KE_n4776, top_core_KE_n4775, top_core_KE_n4774,
         top_core_KE_n4773, top_core_KE_n4772, top_core_KE_n4771,
         top_core_KE_n4770, top_core_KE_n4769, top_core_KE_n4768,
         top_core_KE_n4767, top_core_KE_n4766, top_core_KE_n4765,
         top_core_KE_n4764, top_core_KE_n4763, top_core_KE_n4762,
         top_core_KE_n4761, top_core_KE_n4760, top_core_KE_n4759,
         top_core_KE_n4758, top_core_KE_n4757, top_core_KE_n4756,
         top_core_KE_n4755, top_core_KE_n4754, top_core_KE_n4753,
         top_core_KE_n4752, top_core_KE_n4751, top_core_KE_n4750,
         top_core_KE_n4749, top_core_KE_n4748, top_core_KE_n4747,
         top_core_KE_n4746, top_core_KE_n4745, top_core_KE_n4744,
         top_core_KE_n4743, top_core_KE_n4742, top_core_KE_n4741,
         top_core_KE_n4740, top_core_KE_n4739, top_core_KE_n4738,
         top_core_KE_n4737, top_core_KE_n4736, top_core_KE_n4735,
         top_core_KE_n4734, top_core_KE_n4733, top_core_KE_n4732,
         top_core_KE_n4731, top_core_KE_n4730, top_core_KE_n4729,
         top_core_KE_n4728, top_core_KE_n4727, top_core_KE_n4726,
         top_core_KE_n4725, top_core_KE_n4724, top_core_KE_n4723,
         top_core_KE_n4722, top_core_KE_n4721, top_core_KE_n4720,
         top_core_KE_n4719, top_core_KE_n4718, top_core_KE_n4717,
         top_core_KE_n4716, top_core_KE_n4715, top_core_KE_n4714,
         top_core_KE_n4713, top_core_KE_n4712, top_core_KE_n4711,
         top_core_KE_n4710, top_core_KE_n4709, top_core_KE_n4708,
         top_core_KE_n4707, top_core_KE_n4706, top_core_KE_n4705,
         top_core_KE_n4704, top_core_KE_n4703, top_core_KE_n4702,
         top_core_KE_n4701, top_core_KE_n4700, top_core_KE_n4699,
         top_core_KE_n4698, top_core_KE_n4697, top_core_KE_n4696,
         top_core_KE_n4695, top_core_KE_n4694, top_core_KE_n4693,
         top_core_KE_n4692, top_core_KE_n4691, top_core_KE_n4690,
         top_core_KE_n4689, top_core_KE_n4688, top_core_KE_n4687,
         top_core_KE_n4686, top_core_KE_n4685, top_core_KE_n4684,
         top_core_KE_n4683, top_core_KE_n4682, top_core_KE_n4681,
         top_core_KE_n4680, top_core_KE_n4679, top_core_KE_n4678,
         top_core_KE_n4677, top_core_KE_n4676, top_core_KE_n4675,
         top_core_KE_n4674, top_core_KE_n4673, top_core_KE_n4672,
         top_core_KE_n4671, top_core_KE_n4670, top_core_KE_n4669,
         top_core_KE_n4668, top_core_KE_n4667, top_core_KE_n4666,
         top_core_KE_n4665, top_core_KE_n4664, top_core_KE_n4663,
         top_core_KE_n4662, top_core_KE_n4661, top_core_KE_n4660,
         top_core_KE_n4659, top_core_KE_n4658, top_core_KE_n4657,
         top_core_KE_n4656, top_core_KE_n4655, top_core_KE_n4654,
         top_core_KE_n4653, top_core_KE_n4652, top_core_KE_n4651,
         top_core_KE_n4650, top_core_KE_n4649, top_core_KE_n4648,
         top_core_KE_n4647, top_core_KE_n4646, top_core_KE_n4645,
         top_core_KE_n4644, top_core_KE_n4643, top_core_KE_n4642,
         top_core_KE_n4641, top_core_KE_n4640, top_core_KE_n4639,
         top_core_KE_n4638, top_core_KE_n4637, top_core_KE_n4636,
         top_core_KE_n4635, top_core_KE_n4634, top_core_KE_n4633,
         top_core_KE_n4632, top_core_KE_n4631, top_core_KE_n4630,
         top_core_KE_n4629, top_core_KE_n4628, top_core_KE_n4627,
         top_core_KE_n4626, top_core_KE_n4625, top_core_KE_n4624,
         top_core_KE_n4623, top_core_KE_n4622, top_core_KE_n4621,
         top_core_KE_n4620, top_core_KE_n4619, top_core_KE_n4618,
         top_core_KE_n4617, top_core_KE_n4616, top_core_KE_n4615,
         top_core_KE_n4614, top_core_KE_n4613, top_core_KE_n4612,
         top_core_KE_n4611, top_core_KE_n4610, top_core_KE_n4609,
         top_core_KE_n4608, top_core_KE_n4607, top_core_KE_n4606,
         top_core_KE_n4605, top_core_KE_n4604, top_core_KE_n4603,
         top_core_KE_n4602, top_core_KE_n4601, top_core_KE_n4600,
         top_core_KE_n4599, top_core_KE_n4598, top_core_KE_n4597,
         top_core_KE_n4596, top_core_KE_n4595, top_core_KE_n4594,
         top_core_KE_n4593, top_core_KE_n4592, top_core_KE_n4591,
         top_core_KE_n4590, top_core_KE_n4589, top_core_KE_n4588,
         top_core_KE_n4587, top_core_KE_n4586, top_core_KE_n4585,
         top_core_KE_n4584, top_core_KE_n4583, top_core_KE_n4582,
         top_core_KE_n4581, top_core_KE_n4580, top_core_KE_n4579,
         top_core_KE_n4578, top_core_KE_n4577, top_core_KE_n4576,
         top_core_KE_n4575, top_core_KE_n4574, top_core_KE_n4573,
         top_core_KE_n4572, top_core_KE_n4571, top_core_KE_n4570,
         top_core_KE_n4569, top_core_KE_n4568, top_core_KE_n4567,
         top_core_KE_n4566, top_core_KE_n4565, top_core_KE_n4564,
         top_core_KE_n4563, top_core_KE_n4562, top_core_KE_n4561,
         top_core_KE_n4560, top_core_KE_n4559, top_core_KE_n4558,
         top_core_KE_n4557, top_core_KE_n4556, top_core_KE_n4555,
         top_core_KE_n4554, top_core_KE_n4553, top_core_KE_n4552,
         top_core_KE_n4551, top_core_KE_n4550, top_core_KE_n4549,
         top_core_KE_n4548, top_core_KE_n4547, top_core_KE_n4546,
         top_core_KE_n4545, top_core_KE_n4544, top_core_KE_n4543,
         top_core_KE_n4542, top_core_KE_n4541, top_core_KE_n4540,
         top_core_KE_n4539, top_core_KE_n4538, top_core_KE_n4537,
         top_core_KE_n4536, top_core_KE_n4535, top_core_KE_n4534,
         top_core_KE_n4533, top_core_KE_n4532, top_core_KE_n4531,
         top_core_KE_n4530, top_core_KE_n4529, top_core_KE_n4528,
         top_core_KE_n4527, top_core_KE_n4526, top_core_KE_n4525,
         top_core_KE_n4524, top_core_KE_n4523, top_core_KE_n4522,
         top_core_KE_n4521, top_core_KE_n4520, top_core_KE_n4519,
         top_core_KE_n4518, top_core_KE_n4517, top_core_KE_n4516,
         top_core_KE_n4515, top_core_KE_n4514, top_core_KE_n4513,
         top_core_KE_n4512, top_core_KE_n4511, top_core_KE_n4510,
         top_core_KE_n4509, top_core_KE_n4508, top_core_KE_n4507,
         top_core_KE_n4506, top_core_KE_n4505, top_core_KE_n4504,
         top_core_KE_n4503, top_core_KE_n4502, top_core_KE_n4501,
         top_core_KE_n4500, top_core_KE_n4499, top_core_KE_n4498,
         top_core_KE_n4497, top_core_KE_n4496, top_core_KE_n4495,
         top_core_KE_n4494, top_core_KE_n4493, top_core_KE_n4492,
         top_core_KE_n4491, top_core_KE_n4490, top_core_KE_n4489,
         top_core_KE_n4488, top_core_KE_n4487, top_core_KE_n4486,
         top_core_KE_n4485, top_core_KE_n4484, top_core_KE_n4483,
         top_core_KE_n4482, top_core_KE_n4481, top_core_KE_n4480,
         top_core_KE_n4479, top_core_KE_n4478, top_core_KE_n4477,
         top_core_KE_n4476, top_core_KE_n4475, top_core_KE_n4474,
         top_core_KE_n4473, top_core_KE_n4472, top_core_KE_n4471,
         top_core_KE_n4470, top_core_KE_n4469, top_core_KE_n4468,
         top_core_KE_n4467, top_core_KE_n4466, top_core_KE_n4465,
         top_core_KE_n4464, top_core_KE_n4463, top_core_KE_n4462,
         top_core_KE_n4461, top_core_KE_n4460, top_core_KE_n4459,
         top_core_KE_n4458, top_core_KE_n4457, top_core_KE_n4456,
         top_core_KE_n4455, top_core_KE_n4454, top_core_KE_n4453,
         top_core_KE_n4452, top_core_KE_n4451, top_core_KE_n4450,
         top_core_KE_n4449, top_core_KE_n4448, top_core_KE_n4447,
         top_core_KE_n4446, top_core_KE_n4445, top_core_KE_n4444,
         top_core_KE_n4443, top_core_KE_n4442, top_core_KE_n4441,
         top_core_KE_n4440, top_core_KE_n4439, top_core_KE_n4438,
         top_core_KE_n4437, top_core_KE_n4436, top_core_KE_n4435,
         top_core_KE_n4434, top_core_KE_n4433, top_core_KE_n4432,
         top_core_KE_n4431, top_core_KE_n4430, top_core_KE_n4429,
         top_core_KE_n4428, top_core_KE_n4427, top_core_KE_n4426,
         top_core_KE_n4425, top_core_KE_n4424, top_core_KE_n4423,
         top_core_KE_n4422, top_core_KE_n4421, top_core_KE_n4420,
         top_core_KE_n4419, top_core_KE_n4418, top_core_KE_n4417,
         top_core_KE_n4416, top_core_KE_n4415, top_core_KE_n4414,
         top_core_KE_n4413, top_core_KE_n4412, top_core_KE_n4411,
         top_core_KE_n4410, top_core_KE_n4409, top_core_KE_n4408,
         top_core_KE_n4407, top_core_KE_n4406, top_core_KE_n4405,
         top_core_KE_n4404, top_core_KE_n4403, top_core_KE_n4402,
         top_core_KE_n4401, top_core_KE_n4400, top_core_KE_n4399,
         top_core_KE_n4398, top_core_KE_n4397, top_core_KE_n4396,
         top_core_KE_n4395, top_core_KE_n4394, top_core_KE_n4393,
         top_core_KE_n4392, top_core_KE_n4391, top_core_KE_n4390,
         top_core_KE_n4389, top_core_KE_n4388, top_core_KE_n4387,
         top_core_KE_n4386, top_core_KE_n4385, top_core_KE_n4384,
         top_core_KE_n4383, top_core_KE_n4382, top_core_KE_n4381,
         top_core_KE_n4380, top_core_KE_n4379, top_core_KE_n4378,
         top_core_KE_n4377, top_core_KE_n4376, top_core_KE_n4375,
         top_core_KE_n4374, top_core_KE_n4373, top_core_KE_n4372,
         top_core_KE_n4371, top_core_KE_n4370, top_core_KE_n4369,
         top_core_KE_n4368, top_core_KE_n4367, top_core_KE_n4366,
         top_core_KE_n4365, top_core_KE_n4364, top_core_KE_n4363,
         top_core_KE_n4362, top_core_KE_n4361, top_core_KE_n4360,
         top_core_KE_n4359, top_core_KE_n4358, top_core_KE_n4357,
         top_core_KE_n4356, top_core_KE_n4355, top_core_KE_n4354,
         top_core_KE_n4353, top_core_KE_n4352, top_core_KE_n4351,
         top_core_KE_n4350, top_core_KE_n4349, top_core_KE_n4348,
         top_core_KE_n4347, top_core_KE_n4346, top_core_KE_n4345,
         top_core_KE_n4344, top_core_KE_n4343, top_core_KE_n4342,
         top_core_KE_n4341, top_core_KE_n4340, top_core_KE_n4339,
         top_core_KE_n4338, top_core_KE_n4337, top_core_KE_n4336,
         top_core_KE_n4335, top_core_KE_n4334, top_core_KE_n4333,
         top_core_KE_n4332, top_core_KE_n4331, top_core_KE_n4330,
         top_core_KE_n4329, top_core_KE_n4328, top_core_KE_n4327,
         top_core_KE_n4326, top_core_KE_n4325, top_core_KE_n4324,
         top_core_KE_n4323, top_core_KE_n4322, top_core_KE_n4321,
         top_core_KE_n4320, top_core_KE_n4319, top_core_KE_n4318,
         top_core_KE_n4317, top_core_KE_n4316, top_core_KE_n4315,
         top_core_KE_n4314, top_core_KE_n4313, top_core_KE_n4312,
         top_core_KE_n4311, top_core_KE_n4310, top_core_KE_n4309,
         top_core_KE_n4308, top_core_KE_n4307, top_core_KE_n4306,
         top_core_KE_n4305, top_core_KE_n4304, top_core_KE_n4303,
         top_core_KE_n4302, top_core_KE_n4301, top_core_KE_n4300,
         top_core_KE_n4299, top_core_KE_n4298, top_core_KE_n4297,
         top_core_KE_n4296, top_core_KE_n4295, top_core_KE_n4294,
         top_core_KE_n4293, top_core_KE_n4292, top_core_KE_n4291,
         top_core_KE_n4290, top_core_KE_n4289, top_core_KE_n4288,
         top_core_KE_n4287, top_core_KE_n4286, top_core_KE_n4285,
         top_core_KE_n4284, top_core_KE_n4283, top_core_KE_n4282,
         top_core_KE_n4281, top_core_KE_n4280, top_core_KE_n4279,
         top_core_KE_n4278, top_core_KE_n4277, top_core_KE_n4276,
         top_core_KE_n4275, top_core_KE_n4274, top_core_KE_n4273,
         top_core_KE_n4272, top_core_KE_n4271, top_core_KE_n4270,
         top_core_KE_n4269, top_core_KE_n4268, top_core_KE_n4267,
         top_core_KE_n4266, top_core_KE_n4265, top_core_KE_n4264,
         top_core_KE_n4263, top_core_KE_n4262, top_core_KE_n4261,
         top_core_KE_n4260, top_core_KE_n4259, top_core_KE_n4258,
         top_core_KE_n4257, top_core_KE_n4256, top_core_KE_n4255,
         top_core_KE_n4254, top_core_KE_n4253, top_core_KE_n4252,
         top_core_KE_n4251, top_core_KE_n4250, top_core_KE_n4249,
         top_core_KE_n4248, top_core_KE_n4247, top_core_KE_n4246,
         top_core_KE_n4245, top_core_KE_n4244, top_core_KE_n4243,
         top_core_KE_n4242, top_core_KE_n4241, top_core_KE_n4240,
         top_core_KE_n4239, top_core_KE_n4238, top_core_KE_n4237,
         top_core_KE_n4236, top_core_KE_n4235, top_core_KE_n4234,
         top_core_KE_n4233, top_core_KE_n4232, top_core_KE_n4231,
         top_core_KE_n4230, top_core_KE_n4229, top_core_KE_n4228,
         top_core_KE_n4227, top_core_KE_n4226, top_core_KE_n4225,
         top_core_KE_n4224, top_core_KE_n4223, top_core_KE_n4222,
         top_core_KE_n4221, top_core_KE_n4220, top_core_KE_n4219,
         top_core_KE_n4218, top_core_KE_n4217, top_core_KE_n4216,
         top_core_KE_n4215, top_core_KE_n4214, top_core_KE_n4213,
         top_core_KE_n4212, top_core_KE_n4211, top_core_KE_n4210,
         top_core_KE_n4209, top_core_KE_n4208, top_core_KE_n4207,
         top_core_KE_n4206, top_core_KE_n4205, top_core_KE_n4204,
         top_core_KE_n4203, top_core_KE_n4202, top_core_KE_n4201,
         top_core_KE_n4200, top_core_KE_n4199, top_core_KE_n4198,
         top_core_KE_n4197, top_core_KE_n4196, top_core_KE_n4195,
         top_core_KE_n4194, top_core_KE_n4193, top_core_KE_n4192,
         top_core_KE_n4191, top_core_KE_n4190, top_core_KE_n4189,
         top_core_KE_n4188, top_core_KE_n4187, top_core_KE_n4186,
         top_core_KE_n4185, top_core_KE_n4184, top_core_KE_n4183,
         top_core_KE_n4182, top_core_KE_n4181, top_core_KE_n4180,
         top_core_KE_n4179, top_core_KE_n4178, top_core_KE_n4177,
         top_core_KE_n4176, top_core_KE_n4175, top_core_KE_n4174,
         top_core_KE_n4173, top_core_KE_n4172, top_core_KE_n4171,
         top_core_KE_n4170, top_core_KE_n4169, top_core_KE_n4168,
         top_core_KE_n4167, top_core_KE_n4166, top_core_KE_n4165,
         top_core_KE_n4164, top_core_KE_n4163, top_core_KE_n4162,
         top_core_KE_n4161, top_core_KE_n4160, top_core_KE_n4159,
         top_core_KE_n4158, top_core_KE_n4157, top_core_KE_n4156,
         top_core_KE_n4155, top_core_KE_n4154, top_core_KE_n4153,
         top_core_KE_n4152, top_core_KE_n4151, top_core_KE_n4150,
         top_core_KE_n4149, top_core_KE_n4148, top_core_KE_n4147,
         top_core_KE_n4146, top_core_KE_n4145, top_core_KE_n4144,
         top_core_KE_n4143, top_core_KE_n4142, top_core_KE_n4141,
         top_core_KE_n4140, top_core_KE_n4139, top_core_KE_n4138,
         top_core_KE_n4137, top_core_KE_n4136, top_core_KE_n4135,
         top_core_KE_n4134, top_core_KE_n4133, top_core_KE_n4132,
         top_core_KE_n4131, top_core_KE_n4130, top_core_KE_n4129,
         top_core_KE_n4128, top_core_KE_n4127, top_core_KE_n4126,
         top_core_KE_n4125, top_core_KE_n4124, top_core_KE_n4123,
         top_core_KE_n4122, top_core_KE_n4121, top_core_KE_n4120,
         top_core_KE_n4119, top_core_KE_n4118, top_core_KE_n4117,
         top_core_KE_n4116, top_core_KE_n4115, top_core_KE_n4114,
         top_core_KE_n4113, top_core_KE_n4112, top_core_KE_n4111,
         top_core_KE_n4110, top_core_KE_n4109, top_core_KE_n4108,
         top_core_KE_n4107, top_core_KE_n4106, top_core_KE_n4105,
         top_core_KE_n4104, top_core_KE_n4103, top_core_KE_n4102,
         top_core_KE_n4101, top_core_KE_n4100, top_core_KE_n4099,
         top_core_KE_n4098, top_core_KE_n4097, top_core_KE_n4096,
         top_core_KE_n4095, top_core_KE_n4094, top_core_KE_n4093,
         top_core_KE_n4092, top_core_KE_n4091, top_core_KE_n4090,
         top_core_KE_n4089, top_core_KE_n4088, top_core_KE_n4087,
         top_core_KE_n4086, top_core_KE_n4085, top_core_KE_n4084,
         top_core_KE_n4083, top_core_KE_n4082, top_core_KE_n4081,
         top_core_KE_n4080, top_core_KE_n4079, top_core_KE_n4078,
         top_core_KE_n4077, top_core_KE_n4076, top_core_KE_n4075,
         top_core_KE_n4074, top_core_KE_n4073, top_core_KE_n4072,
         top_core_KE_n4071, top_core_KE_n4070, top_core_KE_n4069,
         top_core_KE_n4068, top_core_KE_n4067, top_core_KE_n4066,
         top_core_KE_n4065, top_core_KE_n4064, top_core_KE_n4063,
         top_core_KE_n4062, top_core_KE_n4061, top_core_KE_n4060,
         top_core_KE_n4059, top_core_KE_n4058, top_core_KE_n4057,
         top_core_KE_n4056, top_core_KE_n4055, top_core_KE_n4054,
         top_core_KE_n4053, top_core_KE_n4052, top_core_KE_n4051,
         top_core_KE_n4050, top_core_KE_n4049, top_core_KE_n4048,
         top_core_KE_n4047, top_core_KE_n4046, top_core_KE_n4045,
         top_core_KE_n4044, top_core_KE_n4043, top_core_KE_n4042,
         top_core_KE_n4041, top_core_KE_n4040, top_core_KE_n4039,
         top_core_KE_n4038, top_core_KE_n4037, top_core_KE_n4036,
         top_core_KE_n4035, top_core_KE_n4034, top_core_KE_n4033,
         top_core_KE_n4032, top_core_KE_n4031, top_core_KE_n4030,
         top_core_KE_n4029, top_core_KE_n4028, top_core_KE_n4027,
         top_core_KE_n4026, top_core_KE_n4025, top_core_KE_n4024,
         top_core_KE_n4023, top_core_KE_n4022, top_core_KE_n4021,
         top_core_KE_n4020, top_core_KE_n4019, top_core_KE_n4018,
         top_core_KE_n4017, top_core_KE_n4016, top_core_KE_n4015,
         top_core_KE_n4014, top_core_KE_n4013, top_core_KE_n4012,
         top_core_KE_n4011, top_core_KE_n4010, top_core_KE_n4009,
         top_core_KE_n4008, top_core_KE_n4007, top_core_KE_n4006,
         top_core_KE_n4005, top_core_KE_n4004, top_core_KE_n4003,
         top_core_KE_n4002, top_core_KE_n4001, top_core_KE_n4000,
         top_core_KE_n3999, top_core_KE_n3998, top_core_KE_n3997,
         top_core_KE_n3996, top_core_KE_n3995, top_core_KE_n3994,
         top_core_KE_n3993, top_core_KE_n3992, top_core_KE_n3991,
         top_core_KE_n3990, top_core_KE_n3989, top_core_KE_n3988,
         top_core_KE_n3987, top_core_KE_n3986, top_core_KE_n3985,
         top_core_KE_n3984, top_core_KE_n3983, top_core_KE_n3982,
         top_core_KE_n3981, top_core_KE_n3980, top_core_KE_n3979,
         top_core_KE_n3978, top_core_KE_n3977, top_core_KE_n3976,
         top_core_KE_n3975, top_core_KE_n3974, top_core_KE_n3973,
         top_core_KE_n3972, top_core_KE_n3971, top_core_KE_n3970,
         top_core_KE_n3969, top_core_KE_n3968, top_core_KE_n3967,
         top_core_KE_n3966, top_core_KE_n3965, top_core_KE_n3964,
         top_core_KE_n3963, top_core_KE_n3962, top_core_KE_n3961,
         top_core_KE_n3960, top_core_KE_n3959, top_core_KE_n3958,
         top_core_KE_n3957, top_core_KE_n3956, top_core_KE_n3955,
         top_core_KE_n3954, top_core_KE_n3953, top_core_KE_n3952,
         top_core_KE_n3951, top_core_KE_n3950, top_core_KE_n3949,
         top_core_KE_n3948, top_core_KE_n3947, top_core_KE_n3946,
         top_core_KE_n3945, top_core_KE_n3944, top_core_KE_n3943,
         top_core_KE_n3942, top_core_KE_n3941, top_core_KE_n3940,
         top_core_KE_n3939, top_core_KE_n3938, top_core_KE_n3937,
         top_core_KE_n3936, top_core_KE_n3935, top_core_KE_n3934,
         top_core_KE_n3933, top_core_KE_n3932, top_core_KE_n3931,
         top_core_KE_n3930, top_core_KE_n3929, top_core_KE_n3928,
         top_core_KE_n3927, top_core_KE_n3926, top_core_KE_n3925,
         top_core_KE_n3924, top_core_KE_n3923, top_core_KE_n3922,
         top_core_KE_n3921, top_core_KE_n3920, top_core_KE_n3919,
         top_core_KE_n3918, top_core_KE_n3917, top_core_KE_n3916,
         top_core_KE_n3915, top_core_KE_n3914, top_core_KE_n3913,
         top_core_KE_n3912, top_core_KE_n3911, top_core_KE_n3910,
         top_core_KE_n3909, top_core_KE_n3908, top_core_KE_n3907,
         top_core_KE_n3906, top_core_KE_n3905, top_core_KE_n3904,
         top_core_KE_n3903, top_core_KE_n3902, top_core_KE_n3901,
         top_core_KE_n3900, top_core_KE_n3899, top_core_KE_n3898,
         top_core_KE_n3897, top_core_KE_n3896, top_core_KE_n3895,
         top_core_KE_n3894, top_core_KE_n3893, top_core_KE_n3892,
         top_core_KE_n3891, top_core_KE_n3890, top_core_KE_n3889,
         top_core_KE_n3888, top_core_KE_n3887, top_core_KE_n3886,
         top_core_KE_n3885, top_core_KE_n3884, top_core_KE_n3883,
         top_core_KE_n3882, top_core_KE_n3881, top_core_KE_n3880,
         top_core_KE_n3879, top_core_KE_n3878, top_core_KE_n3877,
         top_core_KE_n3876, top_core_KE_n3875, top_core_KE_n3874,
         top_core_KE_n3873, top_core_KE_n3872, top_core_KE_n3871,
         top_core_KE_n3870, top_core_KE_n3869, top_core_KE_n3868,
         top_core_KE_n3867, top_core_KE_n3866, top_core_KE_n3865,
         top_core_KE_n3864, top_core_KE_n3863, top_core_KE_n3862,
         top_core_KE_n3861, top_core_KE_n3860, top_core_KE_n3859,
         top_core_KE_n3858, top_core_KE_n3857, top_core_KE_n3856,
         top_core_KE_n3855, top_core_KE_n3854, top_core_KE_n3853,
         top_core_KE_n3852, top_core_KE_n3851, top_core_KE_n3850,
         top_core_KE_n3849, top_core_KE_n3848, top_core_KE_n3847,
         top_core_KE_n3846, top_core_KE_n3845, top_core_KE_n3844,
         top_core_KE_n3843, top_core_KE_n3842, top_core_KE_n3841,
         top_core_KE_n3840, top_core_KE_n3839, top_core_KE_n3838,
         top_core_KE_n3837, top_core_KE_n3836, top_core_KE_n3835,
         top_core_KE_n3834, top_core_KE_n3833, top_core_KE_n3832,
         top_core_KE_n3831, top_core_KE_n3830, top_core_KE_n3829,
         top_core_KE_n3828, top_core_KE_n3827, top_core_KE_n3826,
         top_core_KE_n3825, top_core_KE_n3824, top_core_KE_n3823,
         top_core_KE_n3822, top_core_KE_n3821, top_core_KE_n3820,
         top_core_KE_n3819, top_core_KE_n3818, top_core_KE_n3817,
         top_core_KE_n3816, top_core_KE_n3815, top_core_KE_n3814,
         top_core_KE_n3813, top_core_KE_n3812, top_core_KE_n3811,
         top_core_KE_n3810, top_core_KE_n3809, top_core_KE_n3808,
         top_core_KE_n3807, top_core_KE_n3806, top_core_KE_n3805,
         top_core_KE_n3804, top_core_KE_n3803, top_core_KE_n3802,
         top_core_KE_n3801, top_core_KE_n3800, top_core_KE_n3799,
         top_core_KE_n3798, top_core_KE_n3797, top_core_KE_n3796,
         top_core_KE_n3795, top_core_KE_n3794, top_core_KE_n3793,
         top_core_KE_n3792, top_core_KE_n3791, top_core_KE_n3790,
         top_core_KE_n3789, top_core_KE_n3788, top_core_KE_n3787,
         top_core_KE_n3786, top_core_KE_n3785, top_core_KE_n3784,
         top_core_KE_n3783, top_core_KE_n3782, top_core_KE_n3781,
         top_core_KE_n3780, top_core_KE_n3779, top_core_KE_n3778,
         top_core_KE_n3777, top_core_KE_n3776, top_core_KE_n3775,
         top_core_KE_n3774, top_core_KE_n3773, top_core_KE_n3772,
         top_core_KE_n3771, top_core_KE_n3770, top_core_KE_n3769,
         top_core_KE_n3768, top_core_KE_n3767, top_core_KE_n3766,
         top_core_KE_n3765, top_core_KE_n3764, top_core_KE_n3763,
         top_core_KE_n3762, top_core_KE_n3761, top_core_KE_n3760,
         top_core_KE_n3759, top_core_KE_n3758, top_core_KE_n3757,
         top_core_KE_n3756, top_core_KE_n3755, top_core_KE_n3754,
         top_core_KE_n3753, top_core_KE_n3752, top_core_KE_n3751,
         top_core_KE_n3750, top_core_KE_n3749, top_core_KE_n3748,
         top_core_KE_n3747, top_core_KE_n3746, top_core_KE_n3745,
         top_core_KE_n3744, top_core_KE_n3743, top_core_KE_n3742,
         top_core_KE_n3741, top_core_KE_n3740, top_core_KE_n3739,
         top_core_KE_n3738, top_core_KE_n3737, top_core_KE_n3736,
         top_core_KE_n3735, top_core_KE_n3734, top_core_KE_n3733,
         top_core_KE_n3732, top_core_KE_n3731, top_core_KE_n3730,
         top_core_KE_n3729, top_core_KE_n3728, top_core_KE_n3727,
         top_core_KE_n3726, top_core_KE_n3725, top_core_KE_n3724,
         top_core_KE_n3723, top_core_KE_n3722, top_core_KE_n3721,
         top_core_KE_n3720, top_core_KE_n3719, top_core_KE_n3718,
         top_core_KE_n3717, top_core_KE_n3716, top_core_KE_n3715,
         top_core_KE_n3714, top_core_KE_n3713, top_core_KE_n3712,
         top_core_KE_n3711, top_core_KE_n3710, top_core_KE_n3709,
         top_core_KE_n3708, top_core_KE_n3707, top_core_KE_n3706,
         top_core_KE_n3705, top_core_KE_n3704, top_core_KE_n3703,
         top_core_KE_n3702, top_core_KE_n3701, top_core_KE_n3700,
         top_core_KE_n3699, top_core_KE_n3698, top_core_KE_n3697,
         top_core_KE_n3696, top_core_KE_n3695, top_core_KE_n3694,
         top_core_KE_n3693, top_core_KE_n3692, top_core_KE_n3691,
         top_core_KE_n3690, top_core_KE_n3689, top_core_KE_n3688,
         top_core_KE_n3687, top_core_KE_n3686, top_core_KE_n3685,
         top_core_KE_n3684, top_core_KE_n3683, top_core_KE_n3682,
         top_core_KE_n3681, top_core_KE_n3680, top_core_KE_n3679,
         top_core_KE_n3678, top_core_KE_n3677, top_core_KE_n3676,
         top_core_KE_n3675, top_core_KE_n3674, top_core_KE_n3673,
         top_core_KE_n3672, top_core_KE_n3671, top_core_KE_n3670,
         top_core_KE_n3669, top_core_KE_n3668, top_core_KE_n3667,
         top_core_KE_n3666, top_core_KE_n3665, top_core_KE_n3664,
         top_core_KE_n3663, top_core_KE_n3662, top_core_KE_n3661,
         top_core_KE_n3660, top_core_KE_n3659, top_core_KE_n3658,
         top_core_KE_n3657, top_core_KE_n3656, top_core_KE_n3655,
         top_core_KE_n3654, top_core_KE_n3653, top_core_KE_n3652,
         top_core_KE_n3651, top_core_KE_n3650, top_core_KE_n3649,
         top_core_KE_n3648, top_core_KE_n3647, top_core_KE_n3646,
         top_core_KE_n3645, top_core_KE_n3644, top_core_KE_n3643,
         top_core_KE_n3642, top_core_KE_n3641, top_core_KE_n3640,
         top_core_KE_n3639, top_core_KE_n3638, top_core_KE_n3637,
         top_core_KE_n3636, top_core_KE_n3635, top_core_KE_n3634,
         top_core_KE_n3633, top_core_KE_n3632, top_core_KE_n3631,
         top_core_KE_n3630, top_core_KE_n3629, top_core_KE_n3628,
         top_core_KE_n3627, top_core_KE_n3626, top_core_KE_n3625,
         top_core_KE_n3624, top_core_KE_n3623, top_core_KE_n3622,
         top_core_KE_n3621, top_core_KE_n3620, top_core_KE_n3619,
         top_core_KE_n3618, top_core_KE_n3617, top_core_KE_n3616,
         top_core_KE_n3615, top_core_KE_n3614, top_core_KE_n3613,
         top_core_KE_n3612, top_core_KE_n3611, top_core_KE_n3610,
         top_core_KE_n3609, top_core_KE_n3608, top_core_KE_n3607,
         top_core_KE_n3606, top_core_KE_n3605, top_core_KE_n3604,
         top_core_KE_n3603, top_core_KE_n3602, top_core_KE_n3601,
         top_core_KE_n3600, top_core_KE_n3599, top_core_KE_n3598,
         top_core_KE_n3597, top_core_KE_n3596, top_core_KE_n3595,
         top_core_KE_n3594, top_core_KE_n3593, top_core_KE_n3592,
         top_core_KE_n3591, top_core_KE_n3590, top_core_KE_n3589,
         top_core_KE_n3588, top_core_KE_n3587, top_core_KE_n3586,
         top_core_KE_n3585, top_core_KE_n3584, top_core_KE_n3583,
         top_core_KE_n3582, top_core_KE_n3581, top_core_KE_n3580,
         top_core_KE_n3579, top_core_KE_n3578, top_core_KE_n3577,
         top_core_KE_n3576, top_core_KE_n3575, top_core_KE_n3574,
         top_core_KE_n3573, top_core_KE_n3572, top_core_KE_n3571,
         top_core_KE_n3570, top_core_KE_n3569, top_core_KE_n3568,
         top_core_KE_n3567, top_core_KE_n3566, top_core_KE_n3565,
         top_core_KE_n3564, top_core_KE_n3563, top_core_KE_n3562,
         top_core_KE_n3561, top_core_KE_n3560, top_core_KE_n3559,
         top_core_KE_n3558, top_core_KE_n3557, top_core_KE_n3556,
         top_core_KE_n3555, top_core_KE_n3554, top_core_KE_n3553,
         top_core_KE_n3552, top_core_KE_n3551, top_core_KE_n3550,
         top_core_KE_n3549, top_core_KE_n3548, top_core_KE_n3547,
         top_core_KE_n3546, top_core_KE_n3545, top_core_KE_n3544,
         top_core_KE_n3543, top_core_KE_n3542, top_core_KE_n3541,
         top_core_KE_n3540, top_core_KE_n3539, top_core_KE_n3538,
         top_core_KE_n3537, top_core_KE_n3536, top_core_KE_n3535,
         top_core_KE_n3534, top_core_KE_n3533, top_core_KE_n3532,
         top_core_KE_n3531, top_core_KE_n3530, top_core_KE_n3529,
         top_core_KE_n3528, top_core_KE_n3527, top_core_KE_n3526,
         top_core_KE_n3525, top_core_KE_n3524, top_core_KE_n3523,
         top_core_KE_n3522, top_core_KE_n3521, top_core_KE_n3520,
         top_core_KE_n3519, top_core_KE_n3518, top_core_KE_n3517,
         top_core_KE_n3516, top_core_KE_n3515, top_core_KE_n3514,
         top_core_KE_n3513, top_core_KE_n3512, top_core_KE_n3511,
         top_core_KE_n3510, top_core_KE_n3509, top_core_KE_n3508,
         top_core_KE_n3507, top_core_KE_n3506, top_core_KE_n3505,
         top_core_KE_n3504, top_core_KE_n3503, top_core_KE_n3502,
         top_core_KE_n3501, top_core_KE_n3500, top_core_KE_n3499,
         top_core_KE_n3498, top_core_KE_n3497, top_core_KE_n3496,
         top_core_KE_n3495, top_core_KE_n3494, top_core_KE_n3493,
         top_core_KE_n3492, top_core_KE_n3491, top_core_KE_n3490,
         top_core_KE_n3489, top_core_KE_n3488, top_core_KE_n3487,
         top_core_KE_n3486, top_core_KE_n3485, top_core_KE_n3484,
         top_core_KE_n3483, top_core_KE_n3482, top_core_KE_n3481,
         top_core_KE_n3480, top_core_KE_n3479, top_core_KE_n3478,
         top_core_KE_n3477, top_core_KE_n3476, top_core_KE_n3475,
         top_core_KE_n3474, top_core_KE_n3473, top_core_KE_n3472,
         top_core_KE_n3471, top_core_KE_n3470, top_core_KE_n3469,
         top_core_KE_n3468, top_core_KE_n3467, top_core_KE_n3466,
         top_core_KE_n3465, top_core_KE_n3464, top_core_KE_n3463,
         top_core_KE_n3462, top_core_KE_n3461, top_core_KE_n3460,
         top_core_KE_n3459, top_core_KE_n3458, top_core_KE_n3457,
         top_core_KE_n3456, top_core_KE_n3455, top_core_KE_n3454,
         top_core_KE_n3453, top_core_KE_n3452, top_core_KE_n3451,
         top_core_KE_n3450, top_core_KE_n3449, top_core_KE_n3448,
         top_core_KE_n3447, top_core_KE_n3446, top_core_KE_n3445,
         top_core_KE_n3444, top_core_KE_n3443, top_core_KE_n3442,
         top_core_KE_n3441, top_core_KE_n3440, top_core_KE_n3439,
         top_core_KE_n3438, top_core_KE_n3437, top_core_KE_n3436,
         top_core_KE_n3435, top_core_KE_n3434, top_core_KE_n3433,
         top_core_KE_n3432, top_core_KE_n3431, top_core_KE_n3430,
         top_core_KE_n3429, top_core_KE_n3428, top_core_KE_n3427,
         top_core_KE_n3426, top_core_KE_n3425, top_core_KE_n3424,
         top_core_KE_n3423, top_core_KE_n3422, top_core_KE_n3421,
         top_core_KE_n3420, top_core_KE_n3419, top_core_KE_n3418,
         top_core_KE_n3417, top_core_KE_n3416, top_core_KE_n3415,
         top_core_KE_n3414, top_core_KE_n3413, top_core_KE_n3412,
         top_core_KE_n3411, top_core_KE_n3410, top_core_KE_n3409,
         top_core_KE_n3408, top_core_KE_n3407, top_core_KE_n3406,
         top_core_KE_n3405, top_core_KE_n3404, top_core_KE_n3403,
         top_core_KE_n3402, top_core_KE_n3401, top_core_KE_n3400,
         top_core_KE_n3399, top_core_KE_n3398, top_core_KE_n3397,
         top_core_KE_n3396, top_core_KE_n3395, top_core_KE_n3394,
         top_core_KE_n3393, top_core_KE_n3392, top_core_KE_n3391,
         top_core_KE_n3390, top_core_KE_n3389, top_core_KE_n3388,
         top_core_KE_n3387, top_core_KE_n3386, top_core_KE_n3385,
         top_core_KE_n3384, top_core_KE_n3383, top_core_KE_n3382,
         top_core_KE_n3381, top_core_KE_n3380, top_core_KE_n3379,
         top_core_KE_n3378, top_core_KE_n3377, top_core_KE_n3376,
         top_core_KE_n3375, top_core_KE_n3374, top_core_KE_n3373,
         top_core_KE_n3372, top_core_KE_n3371, top_core_KE_n3370,
         top_core_KE_n3369, top_core_KE_n3368, top_core_KE_n3367,
         top_core_KE_n3366, top_core_KE_n3365, top_core_KE_n3364,
         top_core_KE_n3363, top_core_KE_n3362, top_core_KE_n3361,
         top_core_KE_n3360, top_core_KE_n3359, top_core_KE_n3358,
         top_core_KE_n3357, top_core_KE_n3356, top_core_KE_n3355,
         top_core_KE_n3354, top_core_KE_n3353, top_core_KE_n3352,
         top_core_KE_n3351, top_core_KE_n3350, top_core_KE_n3349,
         top_core_KE_n3348, top_core_KE_n3347, top_core_KE_n3346,
         top_core_KE_n3345, top_core_KE_n3344, top_core_KE_n3343,
         top_core_KE_n3342, top_core_KE_n3341, top_core_KE_n3340,
         top_core_KE_n3339, top_core_KE_n3338, top_core_KE_n3337,
         top_core_KE_n3336, top_core_KE_n3335, top_core_KE_n3334,
         top_core_KE_n3333, top_core_KE_n3332, top_core_KE_n3331,
         top_core_KE_n3330, top_core_KE_n3329, top_core_KE_n3328,
         top_core_KE_n3327, top_core_KE_n3326, top_core_KE_n3325,
         top_core_KE_n3324, top_core_KE_n3323, top_core_KE_n3322,
         top_core_KE_n3321, top_core_KE_n3320, top_core_KE_n3319,
         top_core_KE_n3318, top_core_KE_n3317, top_core_KE_n3316,
         top_core_KE_n3315, top_core_KE_n3314, top_core_KE_n3313,
         top_core_KE_n3312, top_core_KE_n3311, top_core_KE_n3310,
         top_core_KE_n3309, top_core_KE_n3308, top_core_KE_n3307,
         top_core_KE_n3306, top_core_KE_n3305, top_core_KE_n3304,
         top_core_KE_n3303, top_core_KE_n3302, top_core_KE_n3301,
         top_core_KE_n3300, top_core_KE_n3299, top_core_KE_n3298,
         top_core_KE_n3297, top_core_KE_n3296, top_core_KE_n3295,
         top_core_KE_n3294, top_core_KE_n3293, top_core_KE_n3292,
         top_core_KE_n3291, top_core_KE_n3290, top_core_KE_n3289,
         top_core_KE_n3288, top_core_KE_n3287, top_core_KE_n3286,
         top_core_KE_n3285, top_core_KE_n3284, top_core_KE_n3283,
         top_core_KE_n3282, top_core_KE_n3281, top_core_KE_n3280,
         top_core_KE_n3279, top_core_KE_n3278, top_core_KE_n3277,
         top_core_KE_n3276, top_core_KE_n3275, top_core_KE_n3274,
         top_core_KE_n3273, top_core_KE_n3272, top_core_KE_n3271,
         top_core_KE_n3270, top_core_KE_n3269, top_core_KE_n3268,
         top_core_KE_n3267, top_core_KE_n3266, top_core_KE_n3265,
         top_core_KE_n3264, top_core_KE_n3263, top_core_KE_n3262,
         top_core_KE_n3261, top_core_KE_n3260, top_core_KE_n3259,
         top_core_KE_n3258, top_core_KE_n3257, top_core_KE_n3256,
         top_core_KE_n3255, top_core_KE_n3254, top_core_KE_n3253,
         top_core_KE_n3252, top_core_KE_n3251, top_core_KE_n3250,
         top_core_KE_n3249, top_core_KE_n3248, top_core_KE_n3247,
         top_core_KE_n3246, top_core_KE_n3245, top_core_KE_n3244,
         top_core_KE_n3243, top_core_KE_n3242, top_core_KE_n3241,
         top_core_KE_n3240, top_core_KE_n3239, top_core_KE_n3238,
         top_core_KE_n3237, top_core_KE_n3236, top_core_KE_n3235,
         top_core_KE_n3234, top_core_KE_n3233, top_core_KE_n3232,
         top_core_KE_n3231, top_core_KE_n3230, top_core_KE_n3229,
         top_core_KE_n3228, top_core_KE_n3227, top_core_KE_n3226,
         top_core_KE_n3225, top_core_KE_n3224, top_core_KE_n3223,
         top_core_KE_n3222, top_core_KE_n3221, top_core_KE_n3220,
         top_core_KE_n3219, top_core_KE_n3218, top_core_KE_n3217,
         top_core_KE_n3216, top_core_KE_n3215, top_core_KE_n3214,
         top_core_KE_n3213, top_core_KE_n3212, top_core_KE_n3211,
         top_core_KE_n3210, top_core_KE_n3209, top_core_KE_n3208,
         top_core_KE_n3207, top_core_KE_n3206, top_core_KE_n3205,
         top_core_KE_n3204, top_core_KE_n3203, top_core_KE_n3202,
         top_core_KE_n3201, top_core_KE_n3200, top_core_KE_n3199,
         top_core_KE_n3198, top_core_KE_n3197, top_core_KE_n3196,
         top_core_KE_n3195, top_core_KE_n3194, top_core_KE_n3193,
         top_core_KE_n3192, top_core_KE_n3191, top_core_KE_n3190,
         top_core_KE_n3189, top_core_KE_n3188, top_core_KE_n3187,
         top_core_KE_n3186, top_core_KE_n3185, top_core_KE_n3184,
         top_core_KE_n3183, top_core_KE_n3182, top_core_KE_n3181,
         top_core_KE_n3180, top_core_KE_n3179, top_core_KE_n3178,
         top_core_KE_n3177, top_core_KE_n3176, top_core_KE_n3175,
         top_core_KE_n3174, top_core_KE_n3173, top_core_KE_n3172,
         top_core_KE_n3171, top_core_KE_n3170, top_core_KE_n3169,
         top_core_KE_n3168, top_core_KE_n3167, top_core_KE_n3166,
         top_core_KE_n3165, top_core_KE_n3164, top_core_KE_n3163,
         top_core_KE_n3162, top_core_KE_n3161, top_core_KE_n3160,
         top_core_KE_n3159, top_core_KE_n3158, top_core_KE_n3157,
         top_core_KE_n3156, top_core_KE_n3155, top_core_KE_n3154,
         top_core_KE_n3153, top_core_KE_n3152, top_core_KE_n3151,
         top_core_KE_n3150, top_core_KE_n3149, top_core_KE_n3148,
         top_core_KE_n3147, top_core_KE_n3146, top_core_KE_n3145,
         top_core_KE_n3144, top_core_KE_n3143, top_core_KE_n3142,
         top_core_KE_n3141, top_core_KE_n3140, top_core_KE_n3139,
         top_core_KE_n3138, top_core_KE_n3137, top_core_KE_n3136,
         top_core_KE_n3135, top_core_KE_n3134, top_core_KE_n3133,
         top_core_KE_n3132, top_core_KE_n3131, top_core_KE_n3130,
         top_core_KE_n3129, top_core_KE_n3128, top_core_KE_n3127,
         top_core_KE_n3126, top_core_KE_n3125, top_core_KE_n3124,
         top_core_KE_n3123, top_core_KE_n3122, top_core_KE_n3121,
         top_core_KE_n3120, top_core_KE_n3119, top_core_KE_n3118,
         top_core_KE_n3117, top_core_KE_n3116, top_core_KE_n3115,
         top_core_KE_n3114, top_core_KE_n3113, top_core_KE_n3112,
         top_core_KE_n3111, top_core_KE_n3110, top_core_KE_n3109,
         top_core_KE_n3108, top_core_KE_n3107, top_core_KE_n3106,
         top_core_KE_n3105, top_core_KE_n3104, top_core_KE_n3103,
         top_core_KE_n3102, top_core_KE_n3101, top_core_KE_n3100,
         top_core_KE_n3099, top_core_KE_n3098, top_core_KE_n3097,
         top_core_KE_n3096, top_core_KE_n3095, top_core_KE_n3094,
         top_core_KE_n3093, top_core_KE_n3092, top_core_KE_n3091,
         top_core_KE_n3090, top_core_KE_n3089, top_core_KE_n3088,
         top_core_KE_n3087, top_core_KE_n3086, top_core_KE_n3085,
         top_core_KE_n3084, top_core_KE_n3083, top_core_KE_n3082,
         top_core_KE_n3081, top_core_KE_n3080, top_core_KE_n3079,
         top_core_KE_n3078, top_core_KE_n3077, top_core_KE_n3076,
         top_core_KE_n3075, top_core_KE_n3074, top_core_KE_n3073,
         top_core_KE_n3072, top_core_KE_n3071, top_core_KE_n3070,
         top_core_KE_n3069, top_core_KE_n3068, top_core_KE_n3067,
         top_core_KE_n3066, top_core_KE_n3065, top_core_KE_n3064,
         top_core_KE_n3063, top_core_KE_n3062, top_core_KE_n3061,
         top_core_KE_n3060, top_core_KE_n3059, top_core_KE_n3058,
         top_core_KE_n3057, top_core_KE_n3056, top_core_KE_n3055,
         top_core_KE_n3054, top_core_KE_n3053, top_core_KE_n3052,
         top_core_KE_n3051, top_core_KE_n3050, top_core_KE_n3049,
         top_core_KE_n3048, top_core_KE_n3047, top_core_KE_n3046,
         top_core_KE_n3045, top_core_KE_n3044, top_core_KE_n3043,
         top_core_KE_n3042, top_core_KE_n3041, top_core_KE_n3040,
         top_core_KE_n3039, top_core_KE_n3038, top_core_KE_n3037,
         top_core_KE_n3036, top_core_KE_n3035, top_core_KE_n3034,
         top_core_KE_n3033, top_core_KE_n3032, top_core_KE_n3031,
         top_core_KE_n3030, top_core_KE_n3029, top_core_KE_n3028,
         top_core_KE_n3027, top_core_KE_n3026, top_core_KE_n3025,
         top_core_KE_n3024, top_core_KE_n3023, top_core_KE_n3022,
         top_core_KE_n3021, top_core_KE_n3020, top_core_KE_n3019,
         top_core_KE_n3018, top_core_KE_n3017, top_core_KE_n3016,
         top_core_KE_n3015, top_core_KE_n3014, top_core_KE_n3013,
         top_core_KE_n3012, top_core_KE_n3011, top_core_KE_n3010,
         top_core_KE_n3009, top_core_KE_n3008, top_core_KE_n3007,
         top_core_KE_n3006, top_core_KE_n3005, top_core_KE_n3004,
         top_core_KE_n3003, top_core_KE_n3002, top_core_KE_n3001,
         top_core_KE_n3000, top_core_KE_n2999, top_core_KE_n2998,
         top_core_KE_n2997, top_core_KE_n2996, top_core_KE_n2995,
         top_core_KE_n2994, top_core_KE_n2993, top_core_KE_n2992,
         top_core_KE_n2991, top_core_KE_n2990, top_core_KE_n2989,
         top_core_KE_n2988, top_core_KE_n2987, top_core_KE_n2986,
         top_core_KE_n2985, top_core_KE_n2984, top_core_KE_n2983,
         top_core_KE_n2982, top_core_KE_n2981, top_core_KE_n2980,
         top_core_KE_n2979, top_core_KE_n2978, top_core_KE_n2977,
         top_core_KE_n2976, top_core_KE_n2975, top_core_KE_n2974,
         top_core_KE_n2973, top_core_KE_n2972, top_core_KE_n2971,
         top_core_KE_n2970, top_core_KE_n2969, top_core_KE_n2968,
         top_core_KE_n2967, top_core_KE_n2966, top_core_KE_n2965,
         top_core_KE_n2964, top_core_KE_n2963, top_core_KE_n2962,
         top_core_KE_n2961, top_core_KE_n2960, top_core_KE_n2959,
         top_core_KE_n2958, top_core_KE_n2957, top_core_KE_n2956,
         top_core_KE_n2955, top_core_KE_n2954, top_core_KE_n2953,
         top_core_KE_n2952, top_core_KE_n2951, top_core_KE_n2950,
         top_core_KE_n2949, top_core_KE_n2948, top_core_KE_n2947,
         top_core_KE_n2946, top_core_KE_n2945, top_core_KE_n2944,
         top_core_KE_n2943, top_core_KE_n2942, top_core_KE_n2941,
         top_core_KE_n2940, top_core_KE_n2939, top_core_KE_n2938,
         top_core_KE_n2937, top_core_KE_n2936, top_core_KE_n2935,
         top_core_KE_n2934, top_core_KE_n2933, top_core_KE_n2932,
         top_core_KE_n2931, top_core_KE_n2930, top_core_KE_n2929,
         top_core_KE_n2928, top_core_KE_n2927, top_core_KE_n2926,
         top_core_KE_n2925, top_core_KE_n2924, top_core_KE_n2923,
         top_core_KE_n2922, top_core_KE_n2921, top_core_KE_n2920,
         top_core_KE_n2919, top_core_KE_n2918, top_core_KE_n2917,
         top_core_KE_n2916, top_core_KE_n2915, top_core_KE_n2914,
         top_core_KE_n2913, top_core_KE_n2912, top_core_KE_n2911,
         top_core_KE_n2910, top_core_KE_n2909, top_core_KE_n2908,
         top_core_KE_n2907, top_core_KE_n2906, top_core_KE_n2905,
         top_core_KE_n2904, top_core_KE_n2903, top_core_KE_n2902,
         top_core_KE_n2901, top_core_KE_n2900, top_core_KE_n2899,
         top_core_KE_n2898, top_core_KE_n2897, top_core_KE_n2896,
         top_core_KE_n2895, top_core_KE_n2894, top_core_KE_n2893,
         top_core_KE_n2892, top_core_KE_n2891, top_core_KE_n2890,
         top_core_KE_n2889, top_core_KE_n2888, top_core_KE_n2887,
         top_core_KE_n2886, top_core_KE_n2885, top_core_KE_n2884,
         top_core_KE_n2883, top_core_KE_n2882, top_core_KE_n2881,
         top_core_KE_n2880, top_core_KE_n2879, top_core_KE_n2878,
         top_core_KE_n2877, top_core_KE_n2876, top_core_KE_n2875,
         top_core_KE_n2874, top_core_KE_n2873, top_core_KE_n2872,
         top_core_KE_n2871, top_core_KE_n2870, top_core_KE_n2869,
         top_core_KE_n2868, top_core_KE_n2867, top_core_KE_n2866,
         top_core_KE_n2865, top_core_KE_n2864, top_core_KE_n2863,
         top_core_KE_n2862, top_core_KE_n2861, top_core_KE_n2860,
         top_core_KE_n2859, top_core_KE_n2858, top_core_KE_n2857,
         top_core_KE_n2856, top_core_KE_n2855, top_core_KE_n2854,
         top_core_KE_n2853, top_core_KE_n2852, top_core_KE_n2851,
         top_core_KE_n2850, top_core_KE_n2849, top_core_KE_n2848,
         top_core_KE_n2847, top_core_KE_n2846, top_core_KE_n2845,
         top_core_KE_n2844, top_core_KE_n2843, top_core_KE_n2842,
         top_core_KE_n2841, top_core_KE_n2840, top_core_KE_n2839,
         top_core_KE_n2838, top_core_KE_n2837, top_core_KE_n2836,
         top_core_KE_n2835, top_core_KE_n2834, top_core_KE_n2833,
         top_core_KE_n2832, top_core_KE_n2831, top_core_KE_n2830,
         top_core_KE_n2829, top_core_KE_n2828, top_core_KE_n2827,
         top_core_KE_n2826, top_core_KE_n2825, top_core_KE_n2824,
         top_core_KE_n2823, top_core_KE_n2822, top_core_KE_n2821,
         top_core_KE_n2820, top_core_KE_n2819, top_core_KE_n2818,
         top_core_KE_n2817, top_core_KE_n2816, top_core_KE_n2815,
         top_core_KE_n2814, top_core_KE_n2813, top_core_KE_n2812,
         top_core_KE_n2811, top_core_KE_n2810, top_core_KE_n2809,
         top_core_KE_n2808, top_core_KE_n2807, top_core_KE_n2806,
         top_core_KE_n2805, top_core_KE_n2804, top_core_KE_n2803,
         top_core_KE_n2802, top_core_KE_n2801, top_core_KE_n2800,
         top_core_KE_n2799, top_core_KE_n2798, top_core_KE_n2797,
         top_core_KE_n2796, top_core_KE_n2795, top_core_KE_n2794,
         top_core_KE_n2793, top_core_KE_n2792, top_core_KE_n2791,
         top_core_KE_n2790, top_core_KE_n2789, top_core_KE_n2788,
         top_core_KE_n2787, top_core_KE_n2786, top_core_KE_n2785,
         top_core_KE_n2784, top_core_KE_n2783, top_core_KE_n2782,
         top_core_KE_n2781, top_core_KE_n2780, top_core_KE_n2779,
         top_core_KE_n2778, top_core_KE_n2777, top_core_KE_n2776,
         top_core_KE_n2775, top_core_KE_n2774, top_core_KE_n2773,
         top_core_KE_n2772, top_core_KE_n2771, top_core_KE_n2770,
         top_core_KE_n2769, top_core_KE_n2768, top_core_KE_n2767,
         top_core_KE_n2766, top_core_KE_n2765, top_core_KE_n2764,
         top_core_KE_n2763, top_core_KE_n2762, top_core_KE_n2761,
         top_core_KE_n2760, top_core_KE_n2759, top_core_KE_n2758,
         top_core_KE_n2757, top_core_KE_n2756, top_core_KE_n2755,
         top_core_KE_n2754, top_core_KE_n2753, top_core_KE_n2752,
         top_core_KE_n2751, top_core_KE_n2750, top_core_KE_n2749,
         top_core_KE_n2748, top_core_KE_n2747, top_core_KE_n2746,
         top_core_KE_n2745, top_core_KE_n2744, top_core_KE_n2743,
         top_core_KE_n2742, top_core_KE_n2741, top_core_KE_n2740,
         top_core_KE_n2739, top_core_KE_n2738, top_core_KE_n2737,
         top_core_KE_n2736, top_core_KE_n2735, top_core_KE_n2734,
         top_core_KE_n2733, top_core_KE_n2732, top_core_KE_n2731,
         top_core_KE_n2730, top_core_KE_n2729, top_core_KE_n2728,
         top_core_KE_n2727, top_core_KE_n2726, top_core_KE_n2725,
         top_core_KE_n2724, top_core_KE_n2723, top_core_KE_n2722,
         top_core_KE_n2721, top_core_KE_n2720, top_core_KE_n2719,
         top_core_KE_n2718, top_core_KE_n2717, top_core_KE_n2716,
         top_core_KE_n2715, top_core_KE_n2714, top_core_KE_n2712,
         top_core_KE_n2711, top_core_KE_n2710, top_core_KE_n2709,
         top_core_KE_n2708, top_core_KE_n2707, top_core_KE_n2705,
         top_core_KE_n2704, top_core_KE_n2703, top_core_KE_n2702,
         top_core_KE_n2701, top_core_KE_n2700, top_core_KE_n2699,
         top_core_KE_n2698, top_core_KE_n2697, top_core_KE_n2696,
         top_core_KE_n2695, top_core_KE_n2694, top_core_KE_n2693,
         top_core_KE_n2692, top_core_KE_n2691, top_core_KE_n2690,
         top_core_KE_n2689, top_core_KE_n2688, top_core_KE_n2687,
         top_core_KE_n2686, top_core_KE_n2685, top_core_KE_n2684,
         top_core_KE_n2683, top_core_KE_n2682, top_core_KE_n2681,
         top_core_KE_n2680, top_core_KE_n2679, top_core_KE_n2678,
         top_core_KE_n2677, top_core_KE_n2676, top_core_KE_n2675,
         top_core_KE_n2674, top_core_KE_n2673, top_core_KE_n2672,
         top_core_KE_n2671, top_core_KE_n2670, top_core_KE_n2669,
         top_core_KE_n2668, top_core_KE_n2667, top_core_KE_n2666,
         top_core_KE_n2665, top_core_KE_n2664, top_core_KE_n2663,
         top_core_KE_n2662, top_core_KE_n2661, top_core_KE_n2660,
         top_core_KE_n2659, top_core_KE_n2658, top_core_KE_n2657,
         top_core_KE_n2656, top_core_KE_n2655, top_core_KE_n2654,
         top_core_KE_n2653, top_core_KE_n2652, top_core_KE_n2651,
         top_core_KE_n2650, top_core_KE_n2649, top_core_KE_n2648,
         top_core_KE_n2647, top_core_KE_n2646, top_core_KE_n2645,
         top_core_KE_n2644, top_core_KE_n2643, top_core_KE_n2642,
         top_core_KE_n2641, top_core_KE_n2640, top_core_KE_n2639,
         top_core_KE_n2638, top_core_KE_n2637, top_core_KE_n2636,
         top_core_KE_n2635, top_core_KE_n2634, top_core_KE_n2633,
         top_core_KE_n2632, top_core_KE_n2631, top_core_KE_n2630,
         top_core_KE_n2629, top_core_KE_n2628, top_core_KE_n2627,
         top_core_KE_n2626, top_core_KE_n2625, top_core_KE_n2624,
         top_core_KE_n2623, top_core_KE_n2622, top_core_KE_n2621,
         top_core_KE_n2620, top_core_KE_n2619, top_core_KE_n2618,
         top_core_KE_n2617, top_core_KE_n2616, top_core_KE_n2615,
         top_core_KE_n2614, top_core_KE_n2613, top_core_KE_n2612,
         top_core_KE_n2611, top_core_KE_n2610, top_core_KE_n2609,
         top_core_KE_n2608, top_core_KE_n2607, top_core_KE_n2606,
         top_core_KE_n2605, top_core_KE_n2604, top_core_KE_n2603,
         top_core_KE_n2602, top_core_KE_n2601, top_core_KE_n2600,
         top_core_KE_n2599, top_core_KE_n2598, top_core_KE_n2597,
         top_core_KE_n2596, top_core_KE_n2595, top_core_KE_n2594,
         top_core_KE_n2593, top_core_KE_n2592, top_core_KE_n2591,
         top_core_KE_n2590, top_core_KE_n2589, top_core_KE_n2588,
         top_core_KE_n2587, top_core_KE_n2586, top_core_KE_n2585,
         top_core_KE_n2584, top_core_KE_n2583, top_core_KE_n2582,
         top_core_KE_n2581, top_core_KE_n2580, top_core_KE_n2579,
         top_core_KE_n2578, top_core_KE_n2577, top_core_KE_n2576,
         top_core_KE_n2575, top_core_KE_n2574, top_core_KE_n2573,
         top_core_KE_n2572, top_core_KE_n2571, top_core_KE_n2570,
         top_core_KE_n2569, top_core_KE_n2568, top_core_KE_n2567,
         top_core_KE_n2566, top_core_KE_n2565, top_core_KE_n2564,
         top_core_KE_n2563, top_core_KE_n2562, top_core_KE_n2561,
         top_core_KE_n2560, top_core_KE_n2559, top_core_KE_n2558,
         top_core_KE_n2557, top_core_KE_n2556, top_core_KE_n2555,
         top_core_KE_n2554, top_core_KE_n2553, top_core_KE_n2552,
         top_core_KE_n2551, top_core_KE_n2550, top_core_KE_n2549,
         top_core_KE_n2548, top_core_KE_n2547, top_core_KE_n2546,
         top_core_KE_n2545, top_core_KE_n2544, top_core_KE_n2543,
         top_core_KE_n2542, top_core_KE_n2541, top_core_KE_n2540,
         top_core_KE_n2539, top_core_KE_n2538, top_core_KE_n2537,
         top_core_KE_n2536, top_core_KE_n2535, top_core_KE_n2534,
         top_core_KE_n2533, top_core_KE_n2532, top_core_KE_n2531,
         top_core_KE_n2530, top_core_KE_n2529, top_core_KE_n2528,
         top_core_KE_n2527, top_core_KE_n2526, top_core_KE_n2525,
         top_core_KE_n2524, top_core_KE_n2523, top_core_KE_n2522,
         top_core_KE_n2521, top_core_KE_n2520, top_core_KE_n2519,
         top_core_KE_n2518, top_core_KE_n2517, top_core_KE_n2516,
         top_core_KE_n2515, top_core_KE_n2514, top_core_KE_n2513,
         top_core_KE_n2512, top_core_KE_n2511, top_core_KE_n2510,
         top_core_KE_n2509, top_core_KE_n2508, top_core_KE_n2507,
         top_core_KE_n2506, top_core_KE_n2504, top_core_KE_n2503,
         top_core_KE_n2502, top_core_KE_n2501, top_core_KE_n2500,
         top_core_KE_n2499, top_core_KE_n2498, top_core_KE_n2497,
         top_core_KE_n2496, top_core_KE_n2495, top_core_KE_n2494,
         top_core_KE_n2493, top_core_KE_n2492, top_core_KE_n2491,
         top_core_KE_n2490, top_core_KE_n2489, top_core_KE_n2488,
         top_core_KE_n2487, top_core_KE_n2486, top_core_KE_n2485,
         top_core_KE_n2484, top_core_KE_n2483, top_core_KE_n2482,
         top_core_KE_n2481, top_core_KE_n2480, top_core_KE_n2479,
         top_core_KE_n2478, top_core_KE_n2477, top_core_KE_n2476,
         top_core_KE_n2475, top_core_KE_n2474, top_core_KE_n2473,
         top_core_KE_n2472, top_core_KE_n2471, top_core_KE_n2470,
         top_core_KE_n2469, top_core_KE_n2468, top_core_KE_n2467,
         top_core_KE_n2466, top_core_KE_n2465, top_core_KE_n2464,
         top_core_KE_n2463, top_core_KE_n2462, top_core_KE_n2461,
         top_core_KE_n2460, top_core_KE_n2459, top_core_KE_n2458,
         top_core_KE_n2457, top_core_KE_n2456, top_core_KE_n2455,
         top_core_KE_n2454, top_core_KE_n2453, top_core_KE_n2452,
         top_core_KE_n2451, top_core_KE_n2450, top_core_KE_n2449,
         top_core_KE_n2448, top_core_KE_n2447, top_core_KE_n2446,
         top_core_KE_n2445, top_core_KE_n2444, top_core_KE_n2443,
         top_core_KE_n2442, top_core_KE_n2441, top_core_KE_n2440,
         top_core_KE_n2439, top_core_KE_n2438, top_core_KE_n2437,
         top_core_KE_n2436, top_core_KE_n2435, top_core_KE_n2434,
         top_core_KE_n2433, top_core_KE_n2432, top_core_KE_n2431,
         top_core_KE_n2430, top_core_KE_n2429, top_core_KE_n2428,
         top_core_KE_n2427, top_core_KE_n2426, top_core_KE_n2425,
         top_core_KE_n2424, top_core_KE_n2423, top_core_KE_n2422,
         top_core_KE_n2421, top_core_KE_n2420, top_core_KE_n2419,
         top_core_KE_n2418, top_core_KE_n2417, top_core_KE_n2416,
         top_core_KE_n2415, top_core_KE_n2414, top_core_KE_n2413,
         top_core_KE_n2412, top_core_KE_n2411, top_core_KE_n2410,
         top_core_KE_n2409, top_core_KE_n2408, top_core_KE_n2407,
         top_core_KE_n2406, top_core_KE_n2405, top_core_KE_n2404,
         top_core_KE_n2403, top_core_KE_n2402, top_core_KE_n2401,
         top_core_KE_n2400, top_core_KE_n2399, top_core_KE_n2398,
         top_core_KE_n2397, top_core_KE_n2396, top_core_KE_n2395,
         top_core_KE_n2394, top_core_KE_n2393, top_core_KE_n2392,
         top_core_KE_n2391, top_core_KE_n2390, top_core_KE_n2389,
         top_core_KE_n2388, top_core_KE_n2387, top_core_KE_n2386,
         top_core_KE_n2385, top_core_KE_n2384, top_core_KE_n2383,
         top_core_KE_n2382, top_core_KE_n2381, top_core_KE_n2380,
         top_core_KE_n2379, top_core_KE_n2378, top_core_KE_n2377,
         top_core_KE_n2376, top_core_KE_n2375, top_core_KE_n2374,
         top_core_KE_n2373, top_core_KE_n2372, top_core_KE_n2371,
         top_core_KE_n2370, top_core_KE_n2369, top_core_KE_n2368,
         top_core_KE_n2367, top_core_KE_n2366, top_core_KE_n2365,
         top_core_KE_n2364, top_core_KE_n2363, top_core_KE_n2362,
         top_core_KE_n2361, top_core_KE_n2360, top_core_KE_n2359,
         top_core_KE_n2358, top_core_KE_n2357, top_core_KE_n2356,
         top_core_KE_n2355, top_core_KE_n2354, top_core_KE_n2353,
         top_core_KE_n2352, top_core_KE_n2351, top_core_KE_n2350,
         top_core_KE_n2349, top_core_KE_n2348, top_core_KE_n2347,
         top_core_KE_n2346, top_core_KE_n2345, top_core_KE_n2344,
         top_core_KE_n2343, top_core_KE_n2342, top_core_KE_n2341,
         top_core_KE_n2340, top_core_KE_n2339, top_core_KE_n2338,
         top_core_KE_n2337, top_core_KE_n2336, top_core_KE_n2335,
         top_core_KE_n2334, top_core_KE_n2333, top_core_KE_n2332,
         top_core_KE_n2331, top_core_KE_n2330, top_core_KE_n2329,
         top_core_KE_n2328, top_core_KE_n2327, top_core_KE_n2326,
         top_core_KE_n2325, top_core_KE_n2324, top_core_KE_n2323,
         top_core_KE_n2322, top_core_KE_n2321, top_core_KE_n2320,
         top_core_KE_n2319, top_core_KE_n2318, top_core_KE_n2317,
         top_core_KE_n2316, top_core_KE_n2315, top_core_KE_n2314,
         top_core_KE_n2313, top_core_KE_n2312, top_core_KE_n2311,
         top_core_KE_n2310, top_core_KE_n2309, top_core_KE_n2308,
         top_core_KE_n2307, top_core_KE_n2306, top_core_KE_n2305,
         top_core_KE_n2304, top_core_KE_n2303, top_core_KE_n2302,
         top_core_KE_n2301, top_core_KE_n2300, top_core_KE_n2299,
         top_core_KE_n2298, top_core_KE_n2297, top_core_KE_n2296,
         top_core_KE_n2295, top_core_KE_n2294, top_core_KE_n2293,
         top_core_KE_n2292, top_core_KE_n2291, top_core_KE_n2290,
         top_core_KE_n2289, top_core_KE_n2288, top_core_KE_n2287,
         top_core_KE_n2286, top_core_KE_n2285, top_core_KE_n2284,
         top_core_KE_n2283, top_core_KE_n2282, top_core_KE_n2281,
         top_core_KE_n2280, top_core_KE_n2279, top_core_KE_n2278,
         top_core_KE_n2277, top_core_KE_n2276, top_core_KE_n2275,
         top_core_KE_n2274, top_core_KE_n2273, top_core_KE_n2272,
         top_core_KE_n2271, top_core_KE_n2270, top_core_KE_n2269,
         top_core_KE_n2268, top_core_KE_n2267, top_core_KE_n2266,
         top_core_KE_n2265, top_core_KE_n2264, top_core_KE_n2263,
         top_core_KE_n2262, top_core_KE_n2261, top_core_KE_n2260,
         top_core_KE_n2259, top_core_KE_n2258, top_core_KE_n2257,
         top_core_KE_n2256, top_core_KE_n2255, top_core_KE_n2254,
         top_core_KE_n2253, top_core_KE_n2252, top_core_KE_n2251,
         top_core_KE_n2250, top_core_KE_n2249, top_core_KE_n2248,
         top_core_KE_n2247, top_core_KE_n2246, top_core_KE_n2245,
         top_core_KE_n2244, top_core_KE_n2243, top_core_KE_n2242,
         top_core_KE_n2241, top_core_KE_n2240, top_core_KE_n2239,
         top_core_KE_n2238, top_core_KE_n2237, top_core_KE_n2236,
         top_core_KE_n2235, top_core_KE_n2234, top_core_KE_n2233,
         top_core_KE_n2232, top_core_KE_n2231, top_core_KE_n2230,
         top_core_KE_n2229, top_core_KE_n2228, top_core_KE_n2227,
         top_core_KE_n2226, top_core_KE_n2225, top_core_KE_n2224,
         top_core_KE_n2223, top_core_KE_n2222, top_core_KE_n2221,
         top_core_KE_n2220, top_core_KE_n2219, top_core_KE_n2218,
         top_core_KE_n2217, top_core_KE_n2216, top_core_KE_n2215,
         top_core_KE_n2214, top_core_KE_n2213, top_core_KE_n2212,
         top_core_KE_n2211, top_core_KE_n2210, top_core_KE_n2209,
         top_core_KE_n2208, top_core_KE_n2207, top_core_KE_n2206,
         top_core_KE_n2205, top_core_KE_n2204, top_core_KE_n2203,
         top_core_KE_n2202, top_core_KE_n2201, top_core_KE_n2200,
         top_core_KE_n2199, top_core_KE_n2198, top_core_KE_n2197,
         top_core_KE_n2196, top_core_KE_n2195, top_core_KE_n2194,
         top_core_KE_n2193, top_core_KE_n2192, top_core_KE_n2191,
         top_core_KE_n2190, top_core_KE_n2189, top_core_KE_n2188,
         top_core_KE_n2187, top_core_KE_n2186, top_core_KE_n2185,
         top_core_KE_n2184, top_core_KE_n2183, top_core_KE_n2182,
         top_core_KE_n2181, top_core_KE_n2180, top_core_KE_n2179,
         top_core_KE_n2178, top_core_KE_n2176, top_core_KE_n2175,
         top_core_KE_n2174, top_core_KE_n2173, top_core_KE_n2172,
         top_core_KE_n2171, top_core_KE_n2170, top_core_KE_n2169,
         top_core_KE_n2168, top_core_KE_n2167, top_core_KE_n2166,
         top_core_KE_n2165, top_core_KE_n2164, top_core_KE_n2163,
         top_core_KE_n2162, top_core_KE_n2161, top_core_KE_n2160,
         top_core_KE_n2159, top_core_KE_n2158, top_core_KE_n2157,
         top_core_KE_n2156, top_core_KE_n2155, top_core_KE_n2154,
         top_core_KE_n2153, top_core_KE_n2152, top_core_KE_n2151,
         top_core_KE_n2150, top_core_KE_n2149, top_core_KE_n2148,
         top_core_KE_n2147, top_core_KE_n2146, top_core_KE_n2145,
         top_core_KE_n2144, top_core_KE_n2143, top_core_KE_n2142,
         top_core_KE_n2141, top_core_KE_n2140, top_core_KE_n2139,
         top_core_KE_n2138, top_core_KE_n2137, top_core_KE_n2136,
         top_core_KE_n2135, top_core_KE_n2134, top_core_KE_n2133,
         top_core_KE_n2132, top_core_KE_n2131, top_core_KE_n2130,
         top_core_KE_n2129, top_core_KE_n2128, top_core_KE_n2127,
         top_core_KE_n2126, top_core_KE_n2125, top_core_KE_n2124,
         top_core_KE_n2123, top_core_KE_n2122, top_core_KE_n2121,
         top_core_KE_n2120, top_core_KE_n2119, top_core_KE_n2118,
         top_core_KE_n2117, top_core_KE_n2116, top_core_KE_n2115,
         top_core_KE_n2114, top_core_KE_n2113, top_core_KE_n2112,
         top_core_KE_n2111, top_core_KE_n2110, top_core_KE_n2109,
         top_core_KE_n2108, top_core_KE_n2107, top_core_KE_n2106,
         top_core_KE_n2105, top_core_KE_n2104, top_core_KE_n2103,
         top_core_KE_n2102, top_core_KE_n2101, top_core_KE_n2100,
         top_core_KE_n2099, top_core_KE_n2098, top_core_KE_n2097,
         top_core_KE_n2096, top_core_KE_n2095, top_core_KE_n2094,
         top_core_KE_n2093, top_core_KE_n2092, top_core_KE_n2091,
         top_core_KE_n2090, top_core_KE_n2089, top_core_KE_n2088,
         top_core_KE_n2087, top_core_KE_n2086, top_core_KE_n2085,
         top_core_KE_n2084, top_core_KE_n2083, top_core_KE_n2082,
         top_core_KE_n2081, top_core_KE_n2080, top_core_KE_n2079,
         top_core_KE_n2078, top_core_KE_n2077, top_core_KE_n2076,
         top_core_KE_n2075, top_core_KE_n2074, top_core_KE_n2073,
         top_core_KE_n2072, top_core_KE_n2071, top_core_KE_n2070,
         top_core_KE_n2069, top_core_KE_n2068, top_core_KE_n2067,
         top_core_KE_n2066, top_core_KE_n2065, top_core_KE_n2064,
         top_core_KE_n2063, top_core_KE_n2062, top_core_KE_n2061,
         top_core_KE_n2060, top_core_KE_n2059, top_core_KE_n2058,
         top_core_KE_n2057, top_core_KE_n2056, top_core_KE_n2055,
         top_core_KE_n2054, top_core_KE_n2053, top_core_KE_n2052,
         top_core_KE_n2051, top_core_KE_n2050, top_core_KE_n2049,
         top_core_KE_n2048, top_core_KE_n2047, top_core_KE_n2046,
         top_core_KE_n2045, top_core_KE_n2044, top_core_KE_n2043,
         top_core_KE_n2042, top_core_KE_n2041, top_core_KE_n2040,
         top_core_KE_n2039, top_core_KE_n2038, top_core_KE_n2037,
         top_core_KE_n2036, top_core_KE_n2035, top_core_KE_n2034,
         top_core_KE_n2033, top_core_KE_n2032, top_core_KE_n2031,
         top_core_KE_n2030, top_core_KE_n2029, top_core_KE_n2028,
         top_core_KE_n2027, top_core_KE_n2026, top_core_KE_n2025,
         top_core_KE_n2024, top_core_KE_n2023, top_core_KE_n2022,
         top_core_KE_n2021, top_core_KE_n2020, top_core_KE_n2019,
         top_core_KE_n2018, top_core_KE_n2017, top_core_KE_n2016,
         top_core_KE_n2015, top_core_KE_n2014, top_core_KE_n2013,
         top_core_KE_n2012, top_core_KE_n2011, top_core_KE_n2010,
         top_core_KE_n2009, top_core_KE_n2008, top_core_KE_n2007,
         top_core_KE_n2006, top_core_KE_n2005, top_core_KE_n2004,
         top_core_KE_n2003, top_core_KE_n2002, top_core_KE_n2001,
         top_core_KE_n2000, top_core_KE_n1999, top_core_KE_n1998,
         top_core_KE_n1997, top_core_KE_n1996, top_core_KE_n1995,
         top_core_KE_n1994, top_core_KE_n1993, top_core_KE_n1992,
         top_core_KE_n1991, top_core_KE_n1990, top_core_KE_n1989,
         top_core_KE_n1988, top_core_KE_n1987, top_core_KE_n1986,
         top_core_KE_n1985, top_core_KE_n1984, top_core_KE_n1983,
         top_core_KE_n1982, top_core_KE_n1981, top_core_KE_n1980,
         top_core_KE_n1979, top_core_KE_n1978, top_core_KE_n1977,
         top_core_KE_n1976, top_core_KE_n1975, top_core_KE_n1974,
         top_core_KE_n1973, top_core_KE_n1972, top_core_KE_n1971,
         top_core_KE_n1970, top_core_KE_n1969, top_core_KE_n1968,
         top_core_KE_n1967, top_core_KE_n1966, top_core_KE_n1965,
         top_core_KE_n1964, top_core_KE_n1963, top_core_KE_n1962,
         top_core_KE_n1961, top_core_KE_n1960, top_core_KE_n1959,
         top_core_KE_n1958, top_core_KE_n1957, top_core_KE_n1956,
         top_core_KE_n1955, top_core_KE_n1954, top_core_KE_n1953,
         top_core_KE_n1952, top_core_KE_n1951, top_core_KE_n1950,
         top_core_KE_n1949, top_core_KE_n1948, top_core_KE_n1947,
         top_core_KE_n1946, top_core_KE_n1945, top_core_KE_n1944,
         top_core_KE_n1943, top_core_KE_n1942, top_core_KE_n1941,
         top_core_KE_n1940, top_core_KE_n1939, top_core_KE_n1938,
         top_core_KE_n1937, top_core_KE_n1936, top_core_KE_n1935,
         top_core_KE_n1934, top_core_KE_n1933, top_core_KE_n1932,
         top_core_KE_n1931, top_core_KE_n1930, top_core_KE_n1929,
         top_core_KE_n1928, top_core_KE_n1927, top_core_KE_n1926,
         top_core_KE_n1925, top_core_KE_n1924, top_core_KE_n1923,
         top_core_KE_n1922, top_core_KE_n1921, top_core_KE_n1920,
         top_core_KE_n1919, top_core_KE_n1918, top_core_KE_n1917,
         top_core_KE_n1916, top_core_KE_n1915, top_core_KE_n1914,
         top_core_KE_n1913, top_core_KE_n1912, top_core_KE_n1911,
         top_core_KE_n1910, top_core_KE_n1909, top_core_KE_n1908,
         top_core_KE_n1907, top_core_KE_n1906, top_core_KE_n1905,
         top_core_KE_n1904, top_core_KE_n1903, top_core_KE_n1902,
         top_core_KE_n1901, top_core_KE_n1900, top_core_KE_n1899,
         top_core_KE_n1898, top_core_KE_n1897, top_core_KE_n1896,
         top_core_KE_n1895, top_core_KE_n1894, top_core_KE_n1893,
         top_core_KE_n1892, top_core_KE_n1891, top_core_KE_n1890,
         top_core_KE_n1889, top_core_KE_n1888, top_core_KE_n1887,
         top_core_KE_n1886, top_core_KE_n1885, top_core_KE_n1884,
         top_core_KE_n1883, top_core_KE_n1882, top_core_KE_n1881,
         top_core_KE_n1880, top_core_KE_n1879, top_core_KE_n1878,
         top_core_KE_n1877, top_core_KE_n1876, top_core_KE_n1875,
         top_core_KE_n1874, top_core_KE_n1873, top_core_KE_n1871,
         top_core_KE_n1870, top_core_KE_n1869, top_core_KE_n1868,
         top_core_KE_n1867, top_core_KE_n1866, top_core_KE_n1865,
         top_core_KE_n1864, top_core_KE_n1863, top_core_KE_n1862,
         top_core_KE_n1861, top_core_KE_n1860, top_core_KE_n1859,
         top_core_KE_n1858, top_core_KE_n1857, top_core_KE_n1856,
         top_core_KE_n1855, top_core_KE_n1854, top_core_KE_n1853,
         top_core_KE_n1852, top_core_KE_n1851, top_core_KE_n1850,
         top_core_KE_n1849, top_core_KE_n1848, top_core_KE_n1847,
         top_core_KE_n1846, top_core_KE_n1845, top_core_KE_n1844,
         top_core_KE_n1843, top_core_KE_n1842, top_core_KE_n1841,
         top_core_KE_n1840, top_core_KE_n1839, top_core_KE_n1838,
         top_core_KE_n1837, top_core_KE_n1836, top_core_KE_n1835,
         top_core_KE_n1834, top_core_KE_n1833, top_core_KE_n1832,
         top_core_KE_n1831, top_core_KE_n1830, top_core_KE_n1829,
         top_core_KE_n1828, top_core_KE_n1827, top_core_KE_n1826,
         top_core_KE_n1825, top_core_KE_n1824, top_core_KE_n1823,
         top_core_KE_n1822, top_core_KE_n1821, top_core_KE_n1820,
         top_core_KE_n1819, top_core_KE_n1818, top_core_KE_n1817,
         top_core_KE_n1816, top_core_KE_n1815, top_core_KE_n1814,
         top_core_KE_n1813, top_core_KE_n1812, top_core_KE_n1811,
         top_core_KE_n1810, top_core_KE_n1809, top_core_KE_n1808,
         top_core_KE_n1807, top_core_KE_n1806, top_core_KE_n1805,
         top_core_KE_n1804, top_core_KE_n1803, top_core_KE_n1802,
         top_core_KE_n1801, top_core_KE_n1800, top_core_KE_n1799,
         top_core_KE_n1798, top_core_KE_n1797, top_core_KE_n1796,
         top_core_KE_n1795, top_core_KE_n1794, top_core_KE_n1793,
         top_core_KE_n1792, top_core_KE_n1791, top_core_KE_n1790,
         top_core_KE_n1789, top_core_KE_n1788, top_core_KE_n1787,
         top_core_KE_n1786, top_core_KE_n1785, top_core_KE_n1784,
         top_core_KE_n1783, top_core_KE_n1782, top_core_KE_n1781,
         top_core_KE_n1780, top_core_KE_n1779, top_core_KE_n1778,
         top_core_KE_n1777, top_core_KE_n1776, top_core_KE_n1775,
         top_core_KE_n1774, top_core_KE_n1773, top_core_KE_n1772,
         top_core_KE_n1771, top_core_KE_n1770, top_core_KE_n1769,
         top_core_KE_n1768, top_core_KE_n1767, top_core_KE_n1766,
         top_core_KE_n1765, top_core_KE_n1764, top_core_KE_n1763,
         top_core_KE_n1762, top_core_KE_n1761, top_core_KE_n1760,
         top_core_KE_n1759, top_core_KE_n1758, top_core_KE_n1757,
         top_core_KE_n1756, top_core_KE_n1755, top_core_KE_n1754,
         top_core_KE_n1753, top_core_KE_n1752, top_core_KE_n1751,
         top_core_KE_n1750, top_core_KE_n1749, top_core_KE_n1748,
         top_core_KE_n1747, top_core_KE_n1746, top_core_KE_n1745,
         top_core_KE_n1744, top_core_KE_n1743, top_core_KE_n1742,
         top_core_KE_n1741, top_core_KE_n1740, top_core_KE_n1739,
         top_core_KE_n1738, top_core_KE_n1737, top_core_KE_n1736,
         top_core_KE_n1735, top_core_KE_n1734, top_core_KE_n1733,
         top_core_KE_n1732, top_core_KE_n1731, top_core_KE_n1730,
         top_core_KE_n1729, top_core_KE_n1728, top_core_KE_n1727,
         top_core_KE_n1726, top_core_KE_n1725, top_core_KE_n1724,
         top_core_KE_n1723, top_core_KE_n1722, top_core_KE_n1721,
         top_core_KE_n1720, top_core_KE_n1719, top_core_KE_n1718,
         top_core_KE_n1717, top_core_KE_n1716, top_core_KE_n1715,
         top_core_KE_n1714, top_core_KE_n1713, top_core_KE_n1712,
         top_core_KE_n1711, top_core_KE_n1710, top_core_KE_n1709,
         top_core_KE_n1708, top_core_KE_n1707, top_core_KE_n1706,
         top_core_KE_n1705, top_core_KE_n1704, top_core_KE_n1703,
         top_core_KE_n1702, top_core_KE_n1701, top_core_KE_n1700,
         top_core_KE_n1699, top_core_KE_n1698, top_core_KE_n1697,
         top_core_KE_n1696, top_core_KE_n1695, top_core_KE_n1694,
         top_core_KE_n1693, top_core_KE_n1692, top_core_KE_n1691,
         top_core_KE_n1690, top_core_KE_n1689, top_core_KE_n1688,
         top_core_KE_n1687, top_core_KE_n1686, top_core_KE_n1685,
         top_core_KE_n1684, top_core_KE_n1683, top_core_KE_n1682,
         top_core_KE_n1681, top_core_KE_n1680, top_core_KE_n1679,
         top_core_KE_n1678, top_core_KE_n1677, top_core_KE_n1676,
         top_core_KE_n1675, top_core_KE_n1674, top_core_KE_n1673,
         top_core_KE_n1672, top_core_KE_n1671, top_core_KE_n1670,
         top_core_KE_n1669, top_core_KE_n1668, top_core_KE_n1667,
         top_core_KE_n1666, top_core_KE_n1665, top_core_KE_n1664,
         top_core_KE_n1663, top_core_KE_n1662, top_core_KE_n1661,
         top_core_KE_n1660, top_core_KE_n1659, top_core_KE_n1658,
         top_core_KE_n1657, top_core_KE_n1656, top_core_KE_n1655,
         top_core_KE_n1654, top_core_KE_n1653, top_core_KE_n1652,
         top_core_KE_n1651, top_core_KE_n1650, top_core_KE_n1649,
         top_core_KE_n1648, top_core_KE_n1647, top_core_KE_n1646,
         top_core_KE_n1645, top_core_KE_n1644, top_core_KE_n1643,
         top_core_KE_n1642, top_core_KE_n1641, top_core_KE_n1640,
         top_core_KE_n1639, top_core_KE_n1638, top_core_KE_n1637,
         top_core_KE_n1636, top_core_KE_n1635, top_core_KE_n1634,
         top_core_KE_n1633, top_core_KE_n1632, top_core_KE_n1631,
         top_core_KE_n1630, top_core_KE_n1629, top_core_KE_n1628,
         top_core_KE_n1627, top_core_KE_n1626, top_core_KE_n1625,
         top_core_KE_n1624, top_core_KE_n1623, top_core_KE_n1622,
         top_core_KE_n1621, top_core_KE_n1620, top_core_KE_n1619,
         top_core_KE_n1618, top_core_KE_n1617, top_core_KE_n1616,
         top_core_KE_n1615, top_core_KE_n1614, top_core_KE_n1613,
         top_core_KE_n1612, top_core_KE_n1611, top_core_KE_n1610,
         top_core_KE_n1609, top_core_KE_n1608, top_core_KE_n1607,
         top_core_KE_n1606, top_core_KE_n1605, top_core_KE_n1604,
         top_core_KE_n1603, top_core_KE_n1602, top_core_KE_n1601,
         top_core_KE_n1600, top_core_KE_n1599, top_core_KE_n1598,
         top_core_KE_n1597, top_core_KE_n1596, top_core_KE_n1595,
         top_core_KE_n1594, top_core_KE_n1593, top_core_KE_n1592,
         top_core_KE_n1591, top_core_KE_n1590, top_core_KE_n1589,
         top_core_KE_n1588, top_core_KE_n1587, top_core_KE_n1586,
         top_core_KE_n1585, top_core_KE_n1584, top_core_KE_n1583,
         top_core_KE_n1582, top_core_KE_n1581, top_core_KE_n1580,
         top_core_KE_n1579, top_core_KE_n1578, top_core_KE_n1577,
         top_core_KE_n1576, top_core_KE_n1575, top_core_KE_n1574,
         top_core_KE_n1573, top_core_KE_n1572, top_core_KE_n1571,
         top_core_KE_n1570, top_core_KE_n1569, top_core_KE_n1568,
         top_core_KE_n1567, top_core_KE_n1566, top_core_KE_n1565,
         top_core_KE_n1564, top_core_KE_n1563, top_core_KE_n1562,
         top_core_KE_n1561, top_core_KE_n1560, top_core_KE_n1559,
         top_core_KE_n1558, top_core_KE_n1557, top_core_KE_n1556,
         top_core_KE_n1555, top_core_KE_n1554, top_core_KE_n1553,
         top_core_KE_n1552, top_core_KE_n1551, top_core_KE_n1550,
         top_core_KE_n1549, top_core_KE_n1548, top_core_KE_n1547,
         top_core_KE_n1546, top_core_KE_n1545, top_core_KE_n1544,
         top_core_KE_n1543, top_core_KE_n1542, top_core_KE_n1541,
         top_core_KE_n1540, top_core_KE_n1539, top_core_KE_n1538,
         top_core_KE_n1537, top_core_KE_n1536, top_core_KE_n1535,
         top_core_KE_n1534, top_core_KE_n1533, top_core_KE_n1532,
         top_core_KE_n1531, top_core_KE_n1530, top_core_KE_n1529,
         top_core_KE_n1528, top_core_KE_n1527, top_core_KE_n1526,
         top_core_KE_n1525, top_core_KE_n1524, top_core_KE_n1523,
         top_core_KE_n1522, top_core_KE_n1521, top_core_KE_n1520,
         top_core_KE_n1519, top_core_KE_n1518, top_core_KE_n1517,
         top_core_KE_n1516, top_core_KE_n1515, top_core_KE_n1514,
         top_core_KE_n1513, top_core_KE_n1512, top_core_KE_n1511,
         top_core_KE_n1510, top_core_KE_n1509, top_core_KE_n1508,
         top_core_KE_n1507, top_core_KE_n1506, top_core_KE_n1505,
         top_core_KE_n1504, top_core_KE_n1503, top_core_KE_n1502,
         top_core_KE_n1501, top_core_KE_n1500, top_core_KE_n1499,
         top_core_KE_n1498, top_core_KE_n1497, top_core_KE_n1496,
         top_core_KE_n1495, top_core_KE_n1494, top_core_KE_n1493,
         top_core_KE_n1492, top_core_KE_n1491, top_core_KE_n1490,
         top_core_KE_n1489, top_core_KE_n1488, top_core_KE_n1487,
         top_core_KE_n1486, top_core_KE_n1485, top_core_KE_n1484,
         top_core_KE_n1483, top_core_KE_n1482, top_core_KE_n1481,
         top_core_KE_n1480, top_core_KE_n1479, top_core_KE_n1478,
         top_core_KE_n1477, top_core_KE_n1476, top_core_KE_n1475,
         top_core_KE_n1474, top_core_KE_n1473, top_core_KE_n1472,
         top_core_KE_n1471, top_core_KE_n1470, top_core_KE_n1469,
         top_core_KE_n1468, top_core_KE_n1467, top_core_KE_n1466,
         top_core_KE_n1465, top_core_KE_n1464, top_core_KE_n1463,
         top_core_KE_n1462, top_core_KE_n1461, top_core_KE_n1460,
         top_core_KE_n1459, top_core_KE_n1458, top_core_KE_n1457,
         top_core_KE_n1456, top_core_KE_n1455, top_core_KE_n1454,
         top_core_KE_n1453, top_core_KE_n1452, top_core_KE_n1451,
         top_core_KE_n1450, top_core_KE_n1449, top_core_KE_n1448,
         top_core_KE_n1447, top_core_KE_n1446, top_core_KE_n1445,
         top_core_KE_n1444, top_core_KE_n1443, top_core_KE_n1442,
         top_core_KE_n1441, top_core_KE_n1440, top_core_KE_n1439,
         top_core_KE_n1438, top_core_KE_n1437, top_core_KE_n1436,
         top_core_KE_n1435, top_core_KE_n1434, top_core_KE_n1433,
         top_core_KE_n1432, top_core_KE_n1431, top_core_KE_n1430,
         top_core_KE_n1429, top_core_KE_n1428, top_core_KE_n1427,
         top_core_KE_n1426, top_core_KE_n1425, top_core_KE_n1424,
         top_core_KE_n1423, top_core_KE_n1422, top_core_KE_n1421,
         top_core_KE_n1420, top_core_KE_n1419, top_core_KE_n1418,
         top_core_KE_n1417, top_core_KE_n1416, top_core_KE_n1415,
         top_core_KE_n1414, top_core_KE_n1413, top_core_KE_n1412,
         top_core_KE_n1411, top_core_KE_n1410, top_core_KE_n1409,
         top_core_KE_n1408, top_core_KE_n1407, top_core_KE_n1406,
         top_core_KE_n1405, top_core_KE_n1404, top_core_KE_n1403,
         top_core_KE_n1402, top_core_KE_n1401, top_core_KE_n1400,
         top_core_KE_n1399, top_core_KE_n1398, top_core_KE_n1397,
         top_core_KE_n1396, top_core_KE_n1395, top_core_KE_n1394,
         top_core_KE_n1393, top_core_KE_n1392, top_core_KE_n1391,
         top_core_KE_n1390, top_core_KE_n1389, top_core_KE_n1388,
         top_core_KE_n1387, top_core_KE_n1386, top_core_KE_n1385,
         top_core_KE_n1384, top_core_KE_n1383, top_core_KE_n1382,
         top_core_KE_n1381, top_core_KE_n1380, top_core_KE_n1379,
         top_core_KE_n1378, top_core_KE_n1377, top_core_KE_n1376,
         top_core_KE_n1375, top_core_KE_n1374, top_core_KE_n1373,
         top_core_KE_n1372, top_core_KE_n1371, top_core_KE_n1370,
         top_core_KE_n1369, top_core_KE_n1368, top_core_KE_n1367,
         top_core_KE_n1366, top_core_KE_n1365, top_core_KE_n1364,
         top_core_KE_n1363, top_core_KE_n1362, top_core_KE_n1361,
         top_core_KE_n1360, top_core_KE_n1359, top_core_KE_n1358,
         top_core_KE_n1357, top_core_KE_n1356, top_core_KE_n1355,
         top_core_KE_n1354, top_core_KE_n1353, top_core_KE_n1352,
         top_core_KE_n1351, top_core_KE_n1350, top_core_KE_n1349,
         top_core_KE_n1348, top_core_KE_n1347, top_core_KE_n1346,
         top_core_KE_n1345, top_core_KE_n1344, top_core_KE_n1343,
         top_core_KE_n1342, top_core_KE_n1341, top_core_KE_n1340,
         top_core_KE_n1339, top_core_KE_n1338, top_core_KE_n1337,
         top_core_KE_n1336, top_core_KE_n1335, top_core_KE_n1334,
         top_core_KE_n1333, top_core_KE_n1332, top_core_KE_n1331,
         top_core_KE_n1330, top_core_KE_n1329, top_core_KE_n1328,
         top_core_KE_n1327, top_core_KE_n1326, top_core_KE_n1325,
         top_core_KE_n1324, top_core_KE_n1323, top_core_KE_n1322,
         top_core_KE_n1321, top_core_KE_n1320, top_core_KE_n1319,
         top_core_KE_n1318, top_core_KE_n1317, top_core_KE_n1316,
         top_core_KE_n1315, top_core_KE_n1314, top_core_KE_n1313,
         top_core_KE_n1312, top_core_KE_n1311, top_core_KE_n1310,
         top_core_KE_n1309, top_core_KE_n1308, top_core_KE_n1307,
         top_core_KE_n1306, top_core_KE_n1305, top_core_KE_n1304,
         top_core_KE_n1303, top_core_KE_n1302, top_core_KE_n1301,
         top_core_KE_n1300, top_core_KE_n1299, top_core_KE_n1298,
         top_core_KE_n1297, top_core_KE_n1296, top_core_KE_n1295,
         top_core_KE_n1294, top_core_KE_n1293, top_core_KE_n1292,
         top_core_KE_n1291, top_core_KE_n1290, top_core_KE_n1289,
         top_core_KE_n1288, top_core_KE_n1287, top_core_KE_n1286,
         top_core_KE_n1285, top_core_KE_n1284, top_core_KE_n1283,
         top_core_KE_n1282, top_core_KE_n1281, top_core_KE_n1280,
         top_core_KE_n1279, top_core_KE_n1278, top_core_KE_n1277,
         top_core_KE_n1276, top_core_KE_n1275, top_core_KE_n1274,
         top_core_KE_n1273, top_core_KE_n1272, top_core_KE_n1271,
         top_core_KE_n1270, top_core_KE_n1269, top_core_KE_n1268,
         top_core_KE_n1267, top_core_KE_n1266, top_core_KE_n1265,
         top_core_KE_n1264, top_core_KE_n1263, top_core_KE_n1262,
         top_core_KE_n1261, top_core_KE_n1260, top_core_KE_n1259,
         top_core_KE_n1258, top_core_KE_n1257, top_core_KE_n1256,
         top_core_KE_n1255, top_core_KE_n1254, top_core_KE_n1253,
         top_core_KE_n1252, top_core_KE_n1251, top_core_KE_n1250,
         top_core_KE_n1249, top_core_KE_n1248, top_core_KE_n1247,
         top_core_KE_n1246, top_core_KE_n1245, top_core_KE_n1244,
         top_core_KE_n1243, top_core_KE_n1242, top_core_KE_n1241,
         top_core_KE_n1240, top_core_KE_n1239, top_core_KE_n1238,
         top_core_KE_n1237, top_core_KE_n1236, top_core_KE_n1235,
         top_core_KE_n1234, top_core_KE_n1233, top_core_KE_n1232,
         top_core_KE_n1231, top_core_KE_n1230, top_core_KE_n1229,
         top_core_KE_n1228, top_core_KE_n1227, top_core_KE_n1226,
         top_core_KE_n1225, top_core_KE_n1224, top_core_KE_n1223,
         top_core_KE_n1222, top_core_KE_n1221, top_core_KE_n1220,
         top_core_KE_n1219, top_core_KE_n1218, top_core_KE_n1217,
         top_core_KE_n1216, top_core_KE_n1215, top_core_KE_n1214,
         top_core_KE_n1213, top_core_KE_n1212, top_core_KE_n1211,
         top_core_KE_n1210, top_core_KE_n1209, top_core_KE_n1208,
         top_core_KE_n1207, top_core_KE_n1206, top_core_KE_n1205,
         top_core_KE_n1204, top_core_KE_n1203, top_core_KE_n1202,
         top_core_KE_n1201, top_core_KE_n1200, top_core_KE_n1199,
         top_core_KE_n1198, top_core_KE_n1197, top_core_KE_n1196,
         top_core_KE_n1195, top_core_KE_n1194, top_core_KE_n1193,
         top_core_KE_n1192, top_core_KE_n1191, top_core_KE_n1190,
         top_core_KE_n1189, top_core_KE_n1188, top_core_KE_n1187,
         top_core_KE_n1186, top_core_KE_n1185, top_core_KE_n1184,
         top_core_KE_n1183, top_core_KE_n1182, top_core_KE_n1181,
         top_core_KE_n1180, top_core_KE_n1179, top_core_KE_n1178,
         top_core_KE_n1177, top_core_KE_n1176, top_core_KE_n1175,
         top_core_KE_n1174, top_core_KE_n1173, top_core_KE_n1172,
         top_core_KE_n1171, top_core_KE_n1170, top_core_KE_n1169,
         top_core_KE_n1168, top_core_KE_n1167, top_core_KE_n1166,
         top_core_KE_n1165, top_core_KE_n1164, top_core_KE_n1163,
         top_core_KE_n1162, top_core_KE_n1161, top_core_KE_n1160,
         top_core_KE_n1159, top_core_KE_n1158, top_core_KE_n1157,
         top_core_KE_n1156, top_core_KE_n1155, top_core_KE_n1154,
         top_core_KE_n1153, top_core_KE_n1152, top_core_KE_n1151,
         top_core_KE_n1150, top_core_KE_n1149, top_core_KE_n1148,
         top_core_KE_n1147, top_core_KE_n1146, top_core_KE_n1145,
         top_core_KE_n1144, top_core_KE_n1143, top_core_KE_n1142,
         top_core_KE_n1141, top_core_KE_n1140, top_core_KE_n1139,
         top_core_KE_n1138, top_core_KE_n1137, top_core_KE_n1136,
         top_core_KE_n1135, top_core_KE_n1134, top_core_KE_n1133,
         top_core_KE_n1132, top_core_KE_n1131, top_core_KE_n1130,
         top_core_KE_n1129, top_core_KE_n1128, top_core_KE_n1127,
         top_core_KE_n1126, top_core_KE_n1125, top_core_KE_n1124,
         top_core_KE_n1123, top_core_KE_n1122, top_core_KE_n1121,
         top_core_KE_n1120, top_core_KE_n1119, top_core_KE_n1118,
         top_core_KE_n1117, top_core_KE_n1116, top_core_KE_n1115,
         top_core_KE_n1114, top_core_KE_n1113, top_core_KE_n1112,
         top_core_KE_n1111, top_core_KE_n1110, top_core_KE_n1109,
         top_core_KE_n1108, top_core_KE_n1107, top_core_KE_n1106,
         top_core_KE_n1105, top_core_KE_n1104, top_core_KE_n1103,
         top_core_KE_n1102, top_core_KE_n1101, top_core_KE_n1100,
         top_core_KE_n1099, top_core_KE_n1098, top_core_KE_n1097,
         top_core_KE_n1096, top_core_KE_n1095, top_core_KE_n1094,
         top_core_KE_n1093, top_core_KE_n1092, top_core_KE_n1091,
         top_core_KE_n1090, top_core_KE_n1089, top_core_KE_n1088,
         top_core_KE_n1087, top_core_KE_n1086, top_core_KE_n1085,
         top_core_KE_n1084, top_core_KE_n1083, top_core_KE_n1082,
         top_core_KE_n1081, top_core_KE_n1080, top_core_KE_n1079,
         top_core_KE_n1078, top_core_KE_n1077, top_core_KE_n1076,
         top_core_KE_n1075, top_core_KE_n1074, top_core_KE_n1073,
         top_core_KE_n1072, top_core_KE_n1071, top_core_KE_n1070,
         top_core_KE_n1069, top_core_KE_n1068, top_core_KE_n1067,
         top_core_KE_n1066, top_core_KE_n1065, top_core_KE_n1064,
         top_core_KE_n1063, top_core_KE_n1062, top_core_KE_n1061,
         top_core_KE_n1060, top_core_KE_n1059, top_core_KE_n1058,
         top_core_KE_n1057, top_core_KE_n1056, top_core_KE_n1055,
         top_core_KE_n1054, top_core_KE_n1053, top_core_KE_n1052,
         top_core_KE_n1051, top_core_KE_n1050, top_core_KE_n1049,
         top_core_KE_n1048, top_core_KE_n1047, top_core_KE_n1046,
         top_core_KE_n1045, top_core_KE_n1044, top_core_KE_n1043,
         top_core_KE_n1042, top_core_KE_n1041, top_core_KE_n1040,
         top_core_KE_n1039, top_core_KE_n1038, top_core_KE_n1037,
         top_core_KE_n1036, top_core_KE_n1035, top_core_KE_n1034,
         top_core_KE_n1033, top_core_KE_n1032, top_core_KE_n1031,
         top_core_KE_n1030, top_core_KE_n1029, top_core_KE_n1028,
         top_core_KE_n1027, top_core_KE_n1026, top_core_KE_n1025,
         top_core_KE_n1024, top_core_KE_n1023, top_core_KE_n1022,
         top_core_KE_n1021, top_core_KE_n1020, top_core_KE_n1019,
         top_core_KE_n1018, top_core_KE_n1017, top_core_KE_n1016,
         top_core_KE_n1015, top_core_KE_n1014, top_core_KE_n1013,
         top_core_KE_n1012, top_core_KE_n1011, top_core_KE_n1010,
         top_core_KE_n1009, top_core_KE_n1008, top_core_KE_n1007,
         top_core_KE_n1006, top_core_KE_n1005, top_core_KE_n1004,
         top_core_KE_n1003, top_core_KE_n1002, top_core_KE_n1001,
         top_core_KE_n1000, top_core_KE_n999, top_core_KE_n998,
         top_core_KE_n997, top_core_KE_n996, top_core_KE_n995,
         top_core_KE_n994, top_core_KE_n993, top_core_KE_n992,
         top_core_KE_n991, top_core_KE_n990, top_core_KE_n989,
         top_core_KE_n988, top_core_KE_n987, top_core_KE_n986,
         top_core_KE_n985, top_core_KE_n984, top_core_KE_n983,
         top_core_KE_n982, top_core_KE_n981, top_core_KE_n980,
         top_core_KE_n979, top_core_KE_n978, top_core_KE_n977,
         top_core_KE_n976, top_core_KE_n975, top_core_KE_n974,
         top_core_KE_n973, top_core_KE_n972, top_core_KE_n971,
         top_core_KE_n970, top_core_KE_n969, top_core_KE_n968,
         top_core_KE_n967, top_core_KE_n966, top_core_KE_n965,
         top_core_KE_n964, top_core_KE_n963, top_core_KE_n962,
         top_core_KE_n961, top_core_KE_n960, top_core_KE_n959,
         top_core_KE_n958, top_core_KE_n957, top_core_KE_n956,
         top_core_KE_n955, top_core_KE_n954, top_core_KE_n953,
         top_core_KE_n952, top_core_KE_n951, top_core_KE_n950,
         top_core_KE_n949, top_core_KE_n948, top_core_KE_n947,
         top_core_KE_n946, top_core_KE_n945, top_core_KE_n944,
         top_core_KE_n943, top_core_KE_n942, top_core_KE_n941,
         top_core_KE_n940, top_core_KE_n939, top_core_KE_n938,
         top_core_KE_n937, top_core_KE_n936, top_core_KE_n935,
         top_core_KE_n934, top_core_KE_n933, top_core_KE_n932,
         top_core_KE_n931, top_core_KE_n930, top_core_KE_n929,
         top_core_KE_n928, top_core_KE_n927, top_core_KE_n926,
         top_core_KE_n925, top_core_KE_n924, top_core_KE_n923,
         top_core_KE_n922, top_core_KE_n921, top_core_KE_n920,
         top_core_KE_n919, top_core_KE_n918, top_core_KE_n917,
         top_core_KE_n916, top_core_KE_n915, top_core_KE_n914,
         top_core_KE_n913, top_core_KE_n912, top_core_KE_n911,
         top_core_KE_n910, top_core_KE_n909, top_core_KE_n907,
         top_core_KE_n906, top_core_KE_n903, top_core_KE_n902,
         top_core_KE_n901, top_core_KE_n900, top_core_KE_n899,
         top_core_KE_n898, top_core_KE_n897, top_core_KE_n896,
         top_core_KE_n895, top_core_KE_n894, top_core_KE_n892,
         top_core_KE_n891, top_core_KE_n890, top_core_KE_n889,
         top_core_KE_n888, top_core_KE_n887, top_core_KE_n886,
         top_core_KE_n885, top_core_KE_n884, top_core_KE_n883,
         top_core_KE_n882, top_core_KE_n881, top_core_KE_n880,
         top_core_KE_n879, top_core_KE_n878, top_core_KE_n877,
         top_core_KE_n876, top_core_KE_n875, top_core_KE_n874,
         top_core_KE_n873, top_core_KE_n872, top_core_KE_n871,
         top_core_KE_n870, top_core_KE_n869, top_core_KE_n868,
         top_core_KE_n867, top_core_KE_n866, top_core_KE_n865,
         top_core_KE_n864, top_core_KE_n863, top_core_KE_n862,
         top_core_KE_n861, top_core_KE_n860, top_core_KE_n859,
         top_core_KE_n858, top_core_KE_n857, top_core_KE_n856,
         top_core_KE_n855, top_core_KE_n854, top_core_KE_n853,
         top_core_KE_n852, top_core_KE_n851, top_core_KE_n850,
         top_core_KE_n849, top_core_KE_n848, top_core_KE_n847,
         top_core_KE_n846, top_core_KE_n845, top_core_KE_n844,
         top_core_KE_n843, top_core_KE_n842, top_core_KE_n841,
         top_core_KE_n840, top_core_KE_n839, top_core_KE_n838,
         top_core_KE_n837, top_core_KE_n836, top_core_KE_n835,
         top_core_KE_n834, top_core_KE_n833, top_core_KE_n832,
         top_core_KE_n831, top_core_KE_n830, top_core_KE_n829,
         top_core_KE_n828, top_core_KE_n827, top_core_KE_n826,
         top_core_KE_n825, top_core_KE_n824, top_core_KE_n823,
         top_core_KE_n822, top_core_KE_n821, top_core_KE_n820,
         top_core_KE_n819, top_core_KE_n818, top_core_KE_n817,
         top_core_KE_n816, top_core_KE_n815, top_core_KE_n814,
         top_core_KE_n813, top_core_KE_n812, top_core_KE_n811,
         top_core_KE_n810, top_core_KE_n809, top_core_KE_n808,
         top_core_KE_n807, top_core_KE_n806, top_core_KE_n805,
         top_core_KE_n804, top_core_KE_n803, top_core_KE_n802,
         top_core_KE_n801, top_core_KE_n800, top_core_KE_n799,
         top_core_KE_n798, top_core_KE_n797, top_core_KE_n796,
         top_core_KE_n795, top_core_KE_n794, top_core_KE_n793,
         top_core_KE_n792, top_core_KE_n791, top_core_KE_n790,
         top_core_KE_n789, top_core_KE_n788, top_core_KE_n787,
         top_core_KE_n786, top_core_KE_n785, top_core_KE_n784,
         top_core_KE_n783, top_core_KE_n782, top_core_KE_n781,
         top_core_KE_n780, top_core_KE_n779, top_core_KE_n778,
         top_core_KE_n777, top_core_KE_n776, top_core_KE_n775,
         top_core_KE_n774, top_core_KE_n773, top_core_KE_n772,
         top_core_KE_n771, top_core_KE_n770, top_core_KE_n769,
         top_core_KE_n768, top_core_KE_n767, top_core_KE_n766,
         top_core_KE_n765, top_core_KE_n764, top_core_KE_n763,
         top_core_KE_n762, top_core_KE_n761, top_core_KE_n760,
         top_core_KE_n759, top_core_KE_n758, top_core_KE_n757,
         top_core_KE_n756, top_core_KE_n755, top_core_KE_n754,
         top_core_KE_n753, top_core_KE_n752, top_core_KE_n751,
         top_core_KE_n750, top_core_KE_n749, top_core_KE_n748,
         top_core_KE_n747, top_core_KE_n746, top_core_KE_n745,
         top_core_KE_n744, top_core_KE_n743, top_core_KE_n741,
         top_core_KE_n728, top_core_KE_n658, top_core_KE_n657,
         top_core_KE_n656, top_core_KE_n655, top_core_KE_n654,
         top_core_KE_n653, top_core_KE_n652, top_core_KE_n651,
         top_core_KE_n650, top_core_KE_n649, top_core_KE_n648,
         top_core_KE_n647, top_core_KE_n646, top_core_KE_n645,
         top_core_KE_n644, top_core_KE_n643, top_core_KE_n642,
         top_core_KE_n641, top_core_KE_n640, top_core_KE_n639,
         top_core_KE_n638, top_core_KE_n637, top_core_KE_n636,
         top_core_KE_n635, top_core_KE_N1, top_core_KE_N0,
         top_core_KE_prev_key1_reg_0_, top_core_KE_prev_key1_reg_1_,
         top_core_KE_prev_key1_reg_2_, top_core_KE_prev_key1_reg_3_,
         top_core_KE_prev_key1_reg_4_, top_core_KE_prev_key1_reg_5_,
         top_core_KE_prev_key1_reg_6_, top_core_KE_prev_key1_reg_7_,
         top_core_KE_prev_key1_reg_8_, top_core_KE_prev_key1_reg_9_,
         top_core_KE_prev_key1_reg_10_, top_core_KE_prev_key1_reg_11_,
         top_core_KE_prev_key1_reg_12_, top_core_KE_prev_key1_reg_13_,
         top_core_KE_prev_key1_reg_14_, top_core_KE_prev_key1_reg_15_,
         top_core_KE_prev_key1_reg_16_, top_core_KE_prev_key1_reg_17_,
         top_core_KE_prev_key1_reg_18_, top_core_KE_prev_key1_reg_19_,
         top_core_KE_prev_key1_reg_20_, top_core_KE_prev_key1_reg_21_,
         top_core_KE_prev_key1_reg_22_, top_core_KE_prev_key1_reg_23_,
         top_core_KE_prev_key1_reg_24_, top_core_KE_prev_key1_reg_25_,
         top_core_KE_prev_key1_reg_26_, top_core_KE_prev_key1_reg_27_,
         top_core_KE_prev_key1_reg_28_, top_core_KE_prev_key1_reg_29_,
         top_core_KE_prev_key1_reg_30_, top_core_KE_prev_key1_reg_31_,
         top_core_KE_prev_key1_reg_32_, top_core_KE_prev_key1_reg_33_,
         top_core_KE_prev_key1_reg_34_, top_core_KE_prev_key1_reg_35_,
         top_core_KE_prev_key1_reg_36_, top_core_KE_prev_key1_reg_37_,
         top_core_KE_prev_key1_reg_38_, top_core_KE_prev_key1_reg_39_,
         top_core_KE_prev_key1_reg_40_, top_core_KE_prev_key1_reg_41_,
         top_core_KE_prev_key1_reg_42_, top_core_KE_prev_key1_reg_43_,
         top_core_KE_prev_key1_reg_44_, top_core_KE_prev_key1_reg_45_,
         top_core_KE_prev_key1_reg_46_, top_core_KE_prev_key1_reg_47_,
         top_core_KE_prev_key1_reg_48_, top_core_KE_prev_key1_reg_49_,
         top_core_KE_prev_key1_reg_50_, top_core_KE_prev_key1_reg_51_,
         top_core_KE_prev_key1_reg_52_, top_core_KE_prev_key1_reg_53_,
         top_core_KE_prev_key1_reg_54_, top_core_KE_prev_key1_reg_55_,
         top_core_KE_prev_key1_reg_56_, top_core_KE_prev_key1_reg_57_,
         top_core_KE_prev_key1_reg_58_, top_core_KE_prev_key1_reg_59_,
         top_core_KE_prev_key1_reg_60_, top_core_KE_prev_key1_reg_61_,
         top_core_KE_prev_key1_reg_62_, top_core_KE_prev_key1_reg_63_,
         top_core_KE_prev_key1_reg_64_, top_core_KE_prev_key1_reg_65_,
         top_core_KE_prev_key1_reg_66_, top_core_KE_prev_key1_reg_67_,
         top_core_KE_prev_key1_reg_68_, top_core_KE_prev_key1_reg_69_,
         top_core_KE_prev_key1_reg_70_, top_core_KE_prev_key1_reg_71_,
         top_core_KE_prev_key1_reg_72_, top_core_KE_prev_key1_reg_73_,
         top_core_KE_prev_key1_reg_74_, top_core_KE_prev_key1_reg_75_,
         top_core_KE_prev_key1_reg_76_, top_core_KE_prev_key1_reg_77_,
         top_core_KE_prev_key1_reg_78_, top_core_KE_prev_key1_reg_79_,
         top_core_KE_prev_key1_reg_80_, top_core_KE_prev_key1_reg_81_,
         top_core_KE_prev_key1_reg_82_, top_core_KE_prev_key1_reg_83_,
         top_core_KE_prev_key1_reg_84_, top_core_KE_prev_key1_reg_85_,
         top_core_KE_prev_key1_reg_86_, top_core_KE_prev_key1_reg_87_,
         top_core_KE_prev_key1_reg_88_, top_core_KE_prev_key1_reg_89_,
         top_core_KE_prev_key1_reg_90_, top_core_KE_prev_key1_reg_91_,
         top_core_KE_prev_key1_reg_92_, top_core_KE_prev_key1_reg_93_,
         top_core_KE_prev_key1_reg_94_, top_core_KE_prev_key1_reg_95_,
         top_core_KE_prev_key1_reg_96_, top_core_KE_prev_key1_reg_97_,
         top_core_KE_prev_key1_reg_98_, top_core_KE_prev_key1_reg_99_,
         top_core_KE_prev_key1_reg_100_, top_core_KE_prev_key1_reg_101_,
         top_core_KE_prev_key1_reg_102_, top_core_KE_prev_key1_reg_103_,
         top_core_KE_prev_key1_reg_104_, top_core_KE_prev_key1_reg_105_,
         top_core_KE_prev_key1_reg_106_, top_core_KE_prev_key1_reg_107_,
         top_core_KE_prev_key1_reg_108_, top_core_KE_prev_key1_reg_109_,
         top_core_KE_prev_key1_reg_110_, top_core_KE_prev_key1_reg_111_,
         top_core_KE_prev_key1_reg_112_, top_core_KE_prev_key1_reg_113_,
         top_core_KE_prev_key1_reg_114_, top_core_KE_prev_key1_reg_115_,
         top_core_KE_prev_key1_reg_116_, top_core_KE_prev_key1_reg_117_,
         top_core_KE_prev_key1_reg_118_, top_core_KE_prev_key1_reg_119_,
         top_core_KE_prev_key1_reg_120_, top_core_KE_prev_key1_reg_121_,
         top_core_KE_prev_key1_reg_122_, top_core_KE_prev_key1_reg_123_,
         top_core_KE_prev_key1_reg_124_, top_core_KE_prev_key1_reg_125_,
         top_core_KE_prev_key1_reg_126_, top_core_KE_prev_key1_reg_127_,
         top_core_KE_prev_key0_reg_0_, top_core_KE_prev_key0_reg_1_,
         top_core_KE_prev_key0_reg_2_, top_core_KE_prev_key0_reg_3_,
         top_core_KE_prev_key0_reg_4_, top_core_KE_prev_key0_reg_5_,
         top_core_KE_prev_key0_reg_6_, top_core_KE_prev_key0_reg_7_,
         top_core_KE_prev_key0_reg_8_, top_core_KE_prev_key0_reg_9_,
         top_core_KE_prev_key0_reg_10_, top_core_KE_prev_key0_reg_11_,
         top_core_KE_prev_key0_reg_12_, top_core_KE_prev_key0_reg_13_,
         top_core_KE_prev_key0_reg_14_, top_core_KE_prev_key0_reg_15_,
         top_core_KE_prev_key0_reg_16_, top_core_KE_prev_key0_reg_17_,
         top_core_KE_prev_key0_reg_18_, top_core_KE_prev_key0_reg_19_,
         top_core_KE_prev_key0_reg_20_, top_core_KE_prev_key0_reg_21_,
         top_core_KE_prev_key0_reg_22_, top_core_KE_prev_key0_reg_23_,
         top_core_KE_prev_key0_reg_24_, top_core_KE_prev_key0_reg_25_,
         top_core_KE_prev_key0_reg_26_, top_core_KE_prev_key0_reg_27_,
         top_core_KE_prev_key0_reg_28_, top_core_KE_prev_key0_reg_29_,
         top_core_KE_prev_key0_reg_30_, top_core_KE_prev_key0_reg_31_,
         top_core_KE_prev_key0_reg_32_, top_core_KE_prev_key0_reg_33_,
         top_core_KE_prev_key0_reg_34_, top_core_KE_prev_key0_reg_35_,
         top_core_KE_prev_key0_reg_36_, top_core_KE_prev_key0_reg_37_,
         top_core_KE_prev_key0_reg_38_, top_core_KE_prev_key0_reg_39_,
         top_core_KE_prev_key0_reg_40_, top_core_KE_prev_key0_reg_41_,
         top_core_KE_prev_key0_reg_42_, top_core_KE_prev_key0_reg_43_,
         top_core_KE_prev_key0_reg_44_, top_core_KE_prev_key0_reg_45_,
         top_core_KE_prev_key0_reg_46_, top_core_KE_prev_key0_reg_47_,
         top_core_KE_prev_key0_reg_48_, top_core_KE_prev_key0_reg_49_,
         top_core_KE_prev_key0_reg_50_, top_core_KE_prev_key0_reg_51_,
         top_core_KE_prev_key0_reg_52_, top_core_KE_prev_key0_reg_53_,
         top_core_KE_prev_key0_reg_54_, top_core_KE_prev_key0_reg_55_,
         top_core_KE_prev_key0_reg_56_, top_core_KE_prev_key0_reg_57_,
         top_core_KE_prev_key0_reg_58_, top_core_KE_prev_key0_reg_59_,
         top_core_KE_prev_key0_reg_60_, top_core_KE_prev_key0_reg_61_,
         top_core_KE_prev_key0_reg_62_, top_core_KE_prev_key0_reg_63_,
         top_core_KE_prev_key0_reg_88_, top_core_KE_prev_key0_reg_89_,
         top_core_KE_prev_key0_reg_90_, top_core_KE_prev_key0_reg_91_,
         top_core_KE_prev_key0_reg_92_, top_core_KE_prev_key0_reg_93_,
         top_core_KE_prev_key0_reg_94_, top_core_KE_prev_key0_reg_95_,
         top_core_KE_prev_key0_reg_96_, top_core_KE_prev_key0_reg_97_,
         top_core_KE_prev_key0_reg_98_, top_core_KE_prev_key0_reg_99_,
         top_core_KE_prev_key0_reg_100_, top_core_KE_prev_key0_reg_101_,
         top_core_KE_prev_key0_reg_102_, top_core_KE_prev_key0_reg_103_,
         top_core_KE_prev_key0_reg_104_, top_core_KE_prev_key0_reg_105_,
         top_core_KE_prev_key0_reg_106_, top_core_KE_prev_key0_reg_107_,
         top_core_KE_prev_key0_reg_108_, top_core_KE_prev_key0_reg_109_,
         top_core_KE_prev_key0_reg_110_, top_core_KE_prev_key0_reg_111_,
         top_core_KE_prev_key0_reg_112_, top_core_KE_prev_key0_reg_113_,
         top_core_KE_prev_key0_reg_114_, top_core_KE_prev_key0_reg_115_,
         top_core_KE_prev_key0_reg_116_, top_core_KE_prev_key0_reg_117_,
         top_core_KE_prev_key0_reg_118_, top_core_KE_prev_key0_reg_119_,
         top_core_KE_prev_key0_reg_120_, top_core_KE_prev_key0_reg_121_,
         top_core_KE_prev_key0_reg_122_, top_core_KE_prev_key0_reg_123_,
         top_core_KE_prev_key0_reg_124_, top_core_KE_prev_key0_reg_125_,
         top_core_KE_prev_key0_reg_126_, top_core_KE_prev_key0_reg_127_,
         top_core_KE_round_ctr_reg_0_, top_core_KE_round_ctr_reg_1_,
         top_core_KE_round_ctr_reg_2_, top_core_KE_round_ctr_reg_3_,
         top_core_KE_key_mem_ctrl_reg_0_, top_core_KE_key_mem_ctrl_reg_1_,
         top_core_KE_rcon_reg_0_, top_core_KE_rcon_reg_1_,
         top_core_KE_rcon_reg_2_, top_core_KE_rcon_reg_3_,
         top_core_KE_rcon_reg_4_, top_core_KE_rcon_reg_5_,
         top_core_KE_rcon_reg_6_, top_core_KE_rcon_reg_7_,
         top_core_KE_key_mem_14__0_, top_core_KE_key_mem_14__1_,
         top_core_KE_key_mem_14__2_, top_core_KE_key_mem_14__3_,
         top_core_KE_key_mem_14__4_, top_core_KE_key_mem_14__5_,
         top_core_KE_key_mem_14__6_, top_core_KE_key_mem_14__7_,
         top_core_KE_key_mem_14__8_, top_core_KE_key_mem_14__9_,
         top_core_KE_key_mem_14__10_, top_core_KE_key_mem_14__11_,
         top_core_KE_key_mem_14__12_, top_core_KE_key_mem_14__13_,
         top_core_KE_key_mem_14__14_, top_core_KE_key_mem_14__15_,
         top_core_KE_key_mem_14__16_, top_core_KE_key_mem_14__17_,
         top_core_KE_key_mem_14__18_, top_core_KE_key_mem_14__19_,
         top_core_KE_key_mem_14__20_, top_core_KE_key_mem_14__21_,
         top_core_KE_key_mem_14__22_, top_core_KE_key_mem_14__23_,
         top_core_KE_key_mem_14__24_, top_core_KE_key_mem_14__25_,
         top_core_KE_key_mem_14__26_, top_core_KE_key_mem_14__27_,
         top_core_KE_key_mem_14__28_, top_core_KE_key_mem_14__29_,
         top_core_KE_key_mem_14__30_, top_core_KE_key_mem_14__31_,
         top_core_KE_key_mem_14__32_, top_core_KE_key_mem_14__33_,
         top_core_KE_key_mem_14__34_, top_core_KE_key_mem_14__35_,
         top_core_KE_key_mem_14__36_, top_core_KE_key_mem_14__37_,
         top_core_KE_key_mem_14__38_, top_core_KE_key_mem_14__39_,
         top_core_KE_key_mem_14__40_, top_core_KE_key_mem_14__41_,
         top_core_KE_key_mem_14__42_, top_core_KE_key_mem_14__43_,
         top_core_KE_key_mem_14__44_, top_core_KE_key_mem_14__45_,
         top_core_KE_key_mem_14__46_, top_core_KE_key_mem_14__47_,
         top_core_KE_key_mem_14__48_, top_core_KE_key_mem_14__49_,
         top_core_KE_key_mem_14__50_, top_core_KE_key_mem_14__51_,
         top_core_KE_key_mem_14__52_, top_core_KE_key_mem_14__53_,
         top_core_KE_key_mem_14__54_, top_core_KE_key_mem_14__55_,
         top_core_KE_key_mem_14__56_, top_core_KE_key_mem_14__57_,
         top_core_KE_key_mem_14__58_, top_core_KE_key_mem_14__59_,
         top_core_KE_key_mem_14__60_, top_core_KE_key_mem_14__61_,
         top_core_KE_key_mem_14__62_, top_core_KE_key_mem_14__63_,
         top_core_KE_key_mem_14__64_, top_core_KE_key_mem_14__65_,
         top_core_KE_key_mem_14__66_, top_core_KE_key_mem_14__67_,
         top_core_KE_key_mem_14__68_, top_core_KE_key_mem_14__69_,
         top_core_KE_key_mem_14__70_, top_core_KE_key_mem_14__71_,
         top_core_KE_key_mem_14__72_, top_core_KE_key_mem_14__73_,
         top_core_KE_key_mem_14__74_, top_core_KE_key_mem_14__75_,
         top_core_KE_key_mem_14__76_, top_core_KE_key_mem_14__77_,
         top_core_KE_key_mem_14__78_, top_core_KE_key_mem_14__79_,
         top_core_KE_key_mem_14__80_, top_core_KE_key_mem_14__81_,
         top_core_KE_key_mem_14__82_, top_core_KE_key_mem_14__83_,
         top_core_KE_key_mem_14__84_, top_core_KE_key_mem_14__85_,
         top_core_KE_key_mem_14__86_, top_core_KE_key_mem_14__87_,
         top_core_KE_key_mem_14__88_, top_core_KE_key_mem_14__89_,
         top_core_KE_key_mem_14__90_, top_core_KE_key_mem_14__91_,
         top_core_KE_key_mem_14__92_, top_core_KE_key_mem_14__93_,
         top_core_KE_key_mem_14__94_, top_core_KE_key_mem_14__95_,
         top_core_KE_key_mem_14__96_, top_core_KE_key_mem_14__97_,
         top_core_KE_key_mem_14__98_, top_core_KE_key_mem_14__99_,
         top_core_KE_key_mem_14__100_, top_core_KE_key_mem_14__101_,
         top_core_KE_key_mem_14__102_, top_core_KE_key_mem_14__103_,
         top_core_KE_key_mem_14__104_, top_core_KE_key_mem_14__105_,
         top_core_KE_key_mem_14__106_, top_core_KE_key_mem_14__107_,
         top_core_KE_key_mem_14__108_, top_core_KE_key_mem_14__109_,
         top_core_KE_key_mem_14__110_, top_core_KE_key_mem_14__111_,
         top_core_KE_key_mem_14__112_, top_core_KE_key_mem_14__113_,
         top_core_KE_key_mem_14__114_, top_core_KE_key_mem_14__115_,
         top_core_KE_key_mem_14__116_, top_core_KE_key_mem_14__117_,
         top_core_KE_key_mem_14__118_, top_core_KE_key_mem_14__119_,
         top_core_KE_key_mem_14__120_, top_core_KE_key_mem_14__121_,
         top_core_KE_key_mem_14__122_, top_core_KE_key_mem_14__123_,
         top_core_KE_key_mem_14__124_, top_core_KE_key_mem_14__125_,
         top_core_KE_key_mem_14__126_, top_core_KE_key_mem_14__127_,
         top_core_KE_key_mem_14__128_, top_core_KE_key_mem_13__0_,
         top_core_KE_key_mem_13__1_, top_core_KE_key_mem_13__2_,
         top_core_KE_key_mem_13__3_, top_core_KE_key_mem_13__4_,
         top_core_KE_key_mem_13__5_, top_core_KE_key_mem_13__6_,
         top_core_KE_key_mem_13__7_, top_core_KE_key_mem_13__8_,
         top_core_KE_key_mem_13__9_, top_core_KE_key_mem_13__10_,
         top_core_KE_key_mem_13__11_, top_core_KE_key_mem_13__12_,
         top_core_KE_key_mem_13__13_, top_core_KE_key_mem_13__14_,
         top_core_KE_key_mem_13__15_, top_core_KE_key_mem_13__16_,
         top_core_KE_key_mem_13__17_, top_core_KE_key_mem_13__18_,
         top_core_KE_key_mem_13__19_, top_core_KE_key_mem_13__20_,
         top_core_KE_key_mem_13__21_, top_core_KE_key_mem_13__22_,
         top_core_KE_key_mem_13__23_, top_core_KE_key_mem_13__24_,
         top_core_KE_key_mem_13__25_, top_core_KE_key_mem_13__26_,
         top_core_KE_key_mem_13__27_, top_core_KE_key_mem_13__28_,
         top_core_KE_key_mem_13__29_, top_core_KE_key_mem_13__30_,
         top_core_KE_key_mem_13__31_, top_core_KE_key_mem_13__32_,
         top_core_KE_key_mem_13__33_, top_core_KE_key_mem_13__34_,
         top_core_KE_key_mem_13__35_, top_core_KE_key_mem_13__36_,
         top_core_KE_key_mem_13__37_, top_core_KE_key_mem_13__38_,
         top_core_KE_key_mem_13__39_, top_core_KE_key_mem_13__40_,
         top_core_KE_key_mem_13__41_, top_core_KE_key_mem_13__42_,
         top_core_KE_key_mem_13__43_, top_core_KE_key_mem_13__44_,
         top_core_KE_key_mem_13__45_, top_core_KE_key_mem_13__46_,
         top_core_KE_key_mem_13__47_, top_core_KE_key_mem_13__48_,
         top_core_KE_key_mem_13__49_, top_core_KE_key_mem_13__50_,
         top_core_KE_key_mem_13__51_, top_core_KE_key_mem_13__52_,
         top_core_KE_key_mem_13__53_, top_core_KE_key_mem_13__54_,
         top_core_KE_key_mem_13__55_, top_core_KE_key_mem_13__56_,
         top_core_KE_key_mem_13__57_, top_core_KE_key_mem_13__58_,
         top_core_KE_key_mem_13__59_, top_core_KE_key_mem_13__60_,
         top_core_KE_key_mem_13__61_, top_core_KE_key_mem_13__62_,
         top_core_KE_key_mem_13__63_, top_core_KE_key_mem_13__64_,
         top_core_KE_key_mem_13__65_, top_core_KE_key_mem_13__66_,
         top_core_KE_key_mem_13__67_, top_core_KE_key_mem_13__68_,
         top_core_KE_key_mem_13__69_, top_core_KE_key_mem_13__70_,
         top_core_KE_key_mem_13__71_, top_core_KE_key_mem_13__72_,
         top_core_KE_key_mem_13__73_, top_core_KE_key_mem_13__74_,
         top_core_KE_key_mem_13__75_, top_core_KE_key_mem_13__76_,
         top_core_KE_key_mem_13__77_, top_core_KE_key_mem_13__78_,
         top_core_KE_key_mem_13__79_, top_core_KE_key_mem_13__80_,
         top_core_KE_key_mem_13__81_, top_core_KE_key_mem_13__82_,
         top_core_KE_key_mem_13__83_, top_core_KE_key_mem_13__84_,
         top_core_KE_key_mem_13__85_, top_core_KE_key_mem_13__86_,
         top_core_KE_key_mem_13__87_, top_core_KE_key_mem_13__88_,
         top_core_KE_key_mem_13__89_, top_core_KE_key_mem_13__90_,
         top_core_KE_key_mem_13__91_, top_core_KE_key_mem_13__92_,
         top_core_KE_key_mem_13__93_, top_core_KE_key_mem_13__94_,
         top_core_KE_key_mem_13__95_, top_core_KE_key_mem_13__96_,
         top_core_KE_key_mem_13__97_, top_core_KE_key_mem_13__98_,
         top_core_KE_key_mem_13__99_, top_core_KE_key_mem_13__100_,
         top_core_KE_key_mem_13__101_, top_core_KE_key_mem_13__102_,
         top_core_KE_key_mem_13__103_, top_core_KE_key_mem_13__104_,
         top_core_KE_key_mem_13__105_, top_core_KE_key_mem_13__106_,
         top_core_KE_key_mem_13__107_, top_core_KE_key_mem_13__108_,
         top_core_KE_key_mem_13__109_, top_core_KE_key_mem_13__110_,
         top_core_KE_key_mem_13__111_, top_core_KE_key_mem_13__112_,
         top_core_KE_key_mem_13__113_, top_core_KE_key_mem_13__114_,
         top_core_KE_key_mem_13__115_, top_core_KE_key_mem_13__116_,
         top_core_KE_key_mem_13__117_, top_core_KE_key_mem_13__118_,
         top_core_KE_key_mem_13__119_, top_core_KE_key_mem_13__120_,
         top_core_KE_key_mem_13__121_, top_core_KE_key_mem_13__122_,
         top_core_KE_key_mem_13__123_, top_core_KE_key_mem_13__124_,
         top_core_KE_key_mem_13__125_, top_core_KE_key_mem_13__126_,
         top_core_KE_key_mem_13__127_, top_core_KE_key_mem_13__128_,
         top_core_KE_key_mem_12__0_, top_core_KE_key_mem_12__1_,
         top_core_KE_key_mem_12__2_, top_core_KE_key_mem_12__3_,
         top_core_KE_key_mem_12__4_, top_core_KE_key_mem_12__5_,
         top_core_KE_key_mem_12__6_, top_core_KE_key_mem_12__7_,
         top_core_KE_key_mem_12__8_, top_core_KE_key_mem_12__9_,
         top_core_KE_key_mem_12__10_, top_core_KE_key_mem_12__11_,
         top_core_KE_key_mem_12__12_, top_core_KE_key_mem_12__13_,
         top_core_KE_key_mem_12__14_, top_core_KE_key_mem_12__15_,
         top_core_KE_key_mem_12__16_, top_core_KE_key_mem_12__17_,
         top_core_KE_key_mem_12__18_, top_core_KE_key_mem_12__19_,
         top_core_KE_key_mem_12__20_, top_core_KE_key_mem_12__21_,
         top_core_KE_key_mem_12__22_, top_core_KE_key_mem_12__23_,
         top_core_KE_key_mem_12__24_, top_core_KE_key_mem_12__25_,
         top_core_KE_key_mem_12__26_, top_core_KE_key_mem_12__27_,
         top_core_KE_key_mem_12__28_, top_core_KE_key_mem_12__29_,
         top_core_KE_key_mem_12__30_, top_core_KE_key_mem_12__31_,
         top_core_KE_key_mem_12__32_, top_core_KE_key_mem_12__33_,
         top_core_KE_key_mem_12__34_, top_core_KE_key_mem_12__35_,
         top_core_KE_key_mem_12__36_, top_core_KE_key_mem_12__37_,
         top_core_KE_key_mem_12__38_, top_core_KE_key_mem_12__39_,
         top_core_KE_key_mem_12__40_, top_core_KE_key_mem_12__41_,
         top_core_KE_key_mem_12__42_, top_core_KE_key_mem_12__43_,
         top_core_KE_key_mem_12__44_, top_core_KE_key_mem_12__45_,
         top_core_KE_key_mem_12__46_, top_core_KE_key_mem_12__47_,
         top_core_KE_key_mem_12__48_, top_core_KE_key_mem_12__49_,
         top_core_KE_key_mem_12__50_, top_core_KE_key_mem_12__51_,
         top_core_KE_key_mem_12__52_, top_core_KE_key_mem_12__53_,
         top_core_KE_key_mem_12__54_, top_core_KE_key_mem_12__55_,
         top_core_KE_key_mem_12__56_, top_core_KE_key_mem_12__57_,
         top_core_KE_key_mem_12__58_, top_core_KE_key_mem_12__59_,
         top_core_KE_key_mem_12__60_, top_core_KE_key_mem_12__61_,
         top_core_KE_key_mem_12__62_, top_core_KE_key_mem_12__63_,
         top_core_KE_key_mem_12__64_, top_core_KE_key_mem_12__65_,
         top_core_KE_key_mem_12__66_, top_core_KE_key_mem_12__67_,
         top_core_KE_key_mem_12__68_, top_core_KE_key_mem_12__69_,
         top_core_KE_key_mem_12__70_, top_core_KE_key_mem_12__71_,
         top_core_KE_key_mem_12__72_, top_core_KE_key_mem_12__73_,
         top_core_KE_key_mem_12__74_, top_core_KE_key_mem_12__75_,
         top_core_KE_key_mem_12__76_, top_core_KE_key_mem_12__77_,
         top_core_KE_key_mem_12__78_, top_core_KE_key_mem_12__79_,
         top_core_KE_key_mem_12__80_, top_core_KE_key_mem_12__81_,
         top_core_KE_key_mem_12__82_, top_core_KE_key_mem_12__83_,
         top_core_KE_key_mem_12__84_, top_core_KE_key_mem_12__85_,
         top_core_KE_key_mem_12__86_, top_core_KE_key_mem_12__87_,
         top_core_KE_key_mem_12__88_, top_core_KE_key_mem_12__89_,
         top_core_KE_key_mem_12__90_, top_core_KE_key_mem_12__91_,
         top_core_KE_key_mem_12__92_, top_core_KE_key_mem_12__93_,
         top_core_KE_key_mem_12__94_, top_core_KE_key_mem_12__95_,
         top_core_KE_key_mem_12__96_, top_core_KE_key_mem_12__97_,
         top_core_KE_key_mem_12__98_, top_core_KE_key_mem_12__99_,
         top_core_KE_key_mem_12__100_, top_core_KE_key_mem_12__101_,
         top_core_KE_key_mem_12__102_, top_core_KE_key_mem_12__103_,
         top_core_KE_key_mem_12__104_, top_core_KE_key_mem_12__105_,
         top_core_KE_key_mem_12__106_, top_core_KE_key_mem_12__107_,
         top_core_KE_key_mem_12__108_, top_core_KE_key_mem_12__109_,
         top_core_KE_key_mem_12__110_, top_core_KE_key_mem_12__111_,
         top_core_KE_key_mem_12__112_, top_core_KE_key_mem_12__113_,
         top_core_KE_key_mem_12__114_, top_core_KE_key_mem_12__115_,
         top_core_KE_key_mem_12__116_, top_core_KE_key_mem_12__117_,
         top_core_KE_key_mem_12__118_, top_core_KE_key_mem_12__119_,
         top_core_KE_key_mem_12__120_, top_core_KE_key_mem_12__121_,
         top_core_KE_key_mem_12__122_, top_core_KE_key_mem_12__123_,
         top_core_KE_key_mem_12__124_, top_core_KE_key_mem_12__125_,
         top_core_KE_key_mem_12__126_, top_core_KE_key_mem_12__127_,
         top_core_KE_key_mem_12__128_, top_core_KE_key_mem_11__0_,
         top_core_KE_key_mem_11__1_, top_core_KE_key_mem_11__2_,
         top_core_KE_key_mem_11__3_, top_core_KE_key_mem_11__4_,
         top_core_KE_key_mem_11__5_, top_core_KE_key_mem_11__6_,
         top_core_KE_key_mem_11__7_, top_core_KE_key_mem_11__8_,
         top_core_KE_key_mem_11__9_, top_core_KE_key_mem_11__10_,
         top_core_KE_key_mem_11__11_, top_core_KE_key_mem_11__12_,
         top_core_KE_key_mem_11__13_, top_core_KE_key_mem_11__14_,
         top_core_KE_key_mem_11__15_, top_core_KE_key_mem_11__16_,
         top_core_KE_key_mem_11__17_, top_core_KE_key_mem_11__18_,
         top_core_KE_key_mem_11__19_, top_core_KE_key_mem_11__20_,
         top_core_KE_key_mem_11__21_, top_core_KE_key_mem_11__22_,
         top_core_KE_key_mem_11__23_, top_core_KE_key_mem_11__24_,
         top_core_KE_key_mem_11__25_, top_core_KE_key_mem_11__26_,
         top_core_KE_key_mem_11__27_, top_core_KE_key_mem_11__28_,
         top_core_KE_key_mem_11__29_, top_core_KE_key_mem_11__30_,
         top_core_KE_key_mem_11__31_, top_core_KE_key_mem_11__32_,
         top_core_KE_key_mem_11__33_, top_core_KE_key_mem_11__34_,
         top_core_KE_key_mem_11__35_, top_core_KE_key_mem_11__36_,
         top_core_KE_key_mem_11__37_, top_core_KE_key_mem_11__38_,
         top_core_KE_key_mem_11__39_, top_core_KE_key_mem_11__40_,
         top_core_KE_key_mem_11__41_, top_core_KE_key_mem_11__42_,
         top_core_KE_key_mem_11__43_, top_core_KE_key_mem_11__44_,
         top_core_KE_key_mem_11__45_, top_core_KE_key_mem_11__46_,
         top_core_KE_key_mem_11__47_, top_core_KE_key_mem_11__48_,
         top_core_KE_key_mem_11__49_, top_core_KE_key_mem_11__50_,
         top_core_KE_key_mem_11__51_, top_core_KE_key_mem_11__52_,
         top_core_KE_key_mem_11__53_, top_core_KE_key_mem_11__54_,
         top_core_KE_key_mem_11__55_, top_core_KE_key_mem_11__56_,
         top_core_KE_key_mem_11__57_, top_core_KE_key_mem_11__58_,
         top_core_KE_key_mem_11__59_, top_core_KE_key_mem_11__60_,
         top_core_KE_key_mem_11__61_, top_core_KE_key_mem_11__62_,
         top_core_KE_key_mem_11__63_, top_core_KE_key_mem_11__64_,
         top_core_KE_key_mem_11__65_, top_core_KE_key_mem_11__66_,
         top_core_KE_key_mem_11__67_, top_core_KE_key_mem_11__68_,
         top_core_KE_key_mem_11__69_, top_core_KE_key_mem_11__70_,
         top_core_KE_key_mem_11__71_, top_core_KE_key_mem_11__72_,
         top_core_KE_key_mem_11__73_, top_core_KE_key_mem_11__74_,
         top_core_KE_key_mem_11__75_, top_core_KE_key_mem_11__76_,
         top_core_KE_key_mem_11__77_, top_core_KE_key_mem_11__78_,
         top_core_KE_key_mem_11__79_, top_core_KE_key_mem_11__80_,
         top_core_KE_key_mem_11__81_, top_core_KE_key_mem_11__82_,
         top_core_KE_key_mem_11__83_, top_core_KE_key_mem_11__84_,
         top_core_KE_key_mem_11__85_, top_core_KE_key_mem_11__86_,
         top_core_KE_key_mem_11__87_, top_core_KE_key_mem_11__88_,
         top_core_KE_key_mem_11__89_, top_core_KE_key_mem_11__90_,
         top_core_KE_key_mem_11__91_, top_core_KE_key_mem_11__92_,
         top_core_KE_key_mem_11__93_, top_core_KE_key_mem_11__94_,
         top_core_KE_key_mem_11__95_, top_core_KE_key_mem_11__96_,
         top_core_KE_key_mem_11__97_, top_core_KE_key_mem_11__98_,
         top_core_KE_key_mem_11__99_, top_core_KE_key_mem_11__100_,
         top_core_KE_key_mem_11__101_, top_core_KE_key_mem_11__102_,
         top_core_KE_key_mem_11__103_, top_core_KE_key_mem_11__104_,
         top_core_KE_key_mem_11__105_, top_core_KE_key_mem_11__106_,
         top_core_KE_key_mem_11__107_, top_core_KE_key_mem_11__108_,
         top_core_KE_key_mem_11__109_, top_core_KE_key_mem_11__110_,
         top_core_KE_key_mem_11__111_, top_core_KE_key_mem_11__112_,
         top_core_KE_key_mem_11__113_, top_core_KE_key_mem_11__114_,
         top_core_KE_key_mem_11__115_, top_core_KE_key_mem_11__116_,
         top_core_KE_key_mem_11__117_, top_core_KE_key_mem_11__118_,
         top_core_KE_key_mem_11__119_, top_core_KE_key_mem_11__120_,
         top_core_KE_key_mem_11__121_, top_core_KE_key_mem_11__122_,
         top_core_KE_key_mem_11__123_, top_core_KE_key_mem_11__124_,
         top_core_KE_key_mem_11__125_, top_core_KE_key_mem_11__126_,
         top_core_KE_key_mem_11__127_, top_core_KE_key_mem_11__128_,
         top_core_KE_key_mem_10__0_, top_core_KE_key_mem_10__1_,
         top_core_KE_key_mem_10__2_, top_core_KE_key_mem_10__3_,
         top_core_KE_key_mem_10__4_, top_core_KE_key_mem_10__5_,
         top_core_KE_key_mem_10__6_, top_core_KE_key_mem_10__7_,
         top_core_KE_key_mem_10__8_, top_core_KE_key_mem_10__9_,
         top_core_KE_key_mem_10__10_, top_core_KE_key_mem_10__11_,
         top_core_KE_key_mem_10__12_, top_core_KE_key_mem_10__13_,
         top_core_KE_key_mem_10__14_, top_core_KE_key_mem_10__15_,
         top_core_KE_key_mem_10__16_, top_core_KE_key_mem_10__17_,
         top_core_KE_key_mem_10__18_, top_core_KE_key_mem_10__19_,
         top_core_KE_key_mem_10__20_, top_core_KE_key_mem_10__21_,
         top_core_KE_key_mem_10__22_, top_core_KE_key_mem_10__23_,
         top_core_KE_key_mem_10__24_, top_core_KE_key_mem_10__25_,
         top_core_KE_key_mem_10__26_, top_core_KE_key_mem_10__27_,
         top_core_KE_key_mem_10__28_, top_core_KE_key_mem_10__29_,
         top_core_KE_key_mem_10__30_, top_core_KE_key_mem_10__31_,
         top_core_KE_key_mem_10__32_, top_core_KE_key_mem_10__33_,
         top_core_KE_key_mem_10__34_, top_core_KE_key_mem_10__35_,
         top_core_KE_key_mem_10__36_, top_core_KE_key_mem_10__37_,
         top_core_KE_key_mem_10__38_, top_core_KE_key_mem_10__39_,
         top_core_KE_key_mem_10__40_, top_core_KE_key_mem_10__41_,
         top_core_KE_key_mem_10__42_, top_core_KE_key_mem_10__43_,
         top_core_KE_key_mem_10__44_, top_core_KE_key_mem_10__45_,
         top_core_KE_key_mem_10__46_, top_core_KE_key_mem_10__47_,
         top_core_KE_key_mem_10__48_, top_core_KE_key_mem_10__49_,
         top_core_KE_key_mem_10__50_, top_core_KE_key_mem_10__51_,
         top_core_KE_key_mem_10__52_, top_core_KE_key_mem_10__53_,
         top_core_KE_key_mem_10__54_, top_core_KE_key_mem_10__55_,
         top_core_KE_key_mem_10__56_, top_core_KE_key_mem_10__57_,
         top_core_KE_key_mem_10__58_, top_core_KE_key_mem_10__59_,
         top_core_KE_key_mem_10__60_, top_core_KE_key_mem_10__61_,
         top_core_KE_key_mem_10__62_, top_core_KE_key_mem_10__63_,
         top_core_KE_key_mem_10__64_, top_core_KE_key_mem_10__65_,
         top_core_KE_key_mem_10__66_, top_core_KE_key_mem_10__67_,
         top_core_KE_key_mem_10__68_, top_core_KE_key_mem_10__69_,
         top_core_KE_key_mem_10__70_, top_core_KE_key_mem_10__71_,
         top_core_KE_key_mem_10__72_, top_core_KE_key_mem_10__73_,
         top_core_KE_key_mem_10__74_, top_core_KE_key_mem_10__75_,
         top_core_KE_key_mem_10__76_, top_core_KE_key_mem_10__77_,
         top_core_KE_key_mem_10__78_, top_core_KE_key_mem_10__79_,
         top_core_KE_key_mem_10__80_, top_core_KE_key_mem_10__81_,
         top_core_KE_key_mem_10__82_, top_core_KE_key_mem_10__83_,
         top_core_KE_key_mem_10__84_, top_core_KE_key_mem_10__85_,
         top_core_KE_key_mem_10__86_, top_core_KE_key_mem_10__87_,
         top_core_KE_key_mem_10__88_, top_core_KE_key_mem_10__89_,
         top_core_KE_key_mem_10__90_, top_core_KE_key_mem_10__91_,
         top_core_KE_key_mem_10__92_, top_core_KE_key_mem_10__93_,
         top_core_KE_key_mem_10__94_, top_core_KE_key_mem_10__95_,
         top_core_KE_key_mem_10__96_, top_core_KE_key_mem_10__97_,
         top_core_KE_key_mem_10__98_, top_core_KE_key_mem_10__99_,
         top_core_KE_key_mem_10__100_, top_core_KE_key_mem_10__101_,
         top_core_KE_key_mem_10__102_, top_core_KE_key_mem_10__103_,
         top_core_KE_key_mem_10__104_, top_core_KE_key_mem_10__105_,
         top_core_KE_key_mem_10__106_, top_core_KE_key_mem_10__107_,
         top_core_KE_key_mem_10__108_, top_core_KE_key_mem_10__109_,
         top_core_KE_key_mem_10__110_, top_core_KE_key_mem_10__111_,
         top_core_KE_key_mem_10__112_, top_core_KE_key_mem_10__113_,
         top_core_KE_key_mem_10__114_, top_core_KE_key_mem_10__115_,
         top_core_KE_key_mem_10__116_, top_core_KE_key_mem_10__117_,
         top_core_KE_key_mem_10__118_, top_core_KE_key_mem_10__119_,
         top_core_KE_key_mem_10__120_, top_core_KE_key_mem_10__121_,
         top_core_KE_key_mem_10__122_, top_core_KE_key_mem_10__123_,
         top_core_KE_key_mem_10__124_, top_core_KE_key_mem_10__125_,
         top_core_KE_key_mem_10__126_, top_core_KE_key_mem_10__127_,
         top_core_KE_key_mem_10__128_, top_core_KE_key_mem_9__0_,
         top_core_KE_key_mem_9__1_, top_core_KE_key_mem_9__2_,
         top_core_KE_key_mem_9__3_, top_core_KE_key_mem_9__4_,
         top_core_KE_key_mem_9__5_, top_core_KE_key_mem_9__6_,
         top_core_KE_key_mem_9__7_, top_core_KE_key_mem_9__8_,
         top_core_KE_key_mem_9__9_, top_core_KE_key_mem_9__10_,
         top_core_KE_key_mem_9__11_, top_core_KE_key_mem_9__12_,
         top_core_KE_key_mem_9__13_, top_core_KE_key_mem_9__14_,
         top_core_KE_key_mem_9__15_, top_core_KE_key_mem_9__16_,
         top_core_KE_key_mem_9__17_, top_core_KE_key_mem_9__18_,
         top_core_KE_key_mem_9__19_, top_core_KE_key_mem_9__20_,
         top_core_KE_key_mem_9__21_, top_core_KE_key_mem_9__22_,
         top_core_KE_key_mem_9__23_, top_core_KE_key_mem_9__24_,
         top_core_KE_key_mem_9__25_, top_core_KE_key_mem_9__26_,
         top_core_KE_key_mem_9__27_, top_core_KE_key_mem_9__28_,
         top_core_KE_key_mem_9__29_, top_core_KE_key_mem_9__30_,
         top_core_KE_key_mem_9__31_, top_core_KE_key_mem_9__32_,
         top_core_KE_key_mem_9__33_, top_core_KE_key_mem_9__34_,
         top_core_KE_key_mem_9__35_, top_core_KE_key_mem_9__36_,
         top_core_KE_key_mem_9__37_, top_core_KE_key_mem_9__38_,
         top_core_KE_key_mem_9__39_, top_core_KE_key_mem_9__40_,
         top_core_KE_key_mem_9__41_, top_core_KE_key_mem_9__42_,
         top_core_KE_key_mem_9__43_, top_core_KE_key_mem_9__44_,
         top_core_KE_key_mem_9__45_, top_core_KE_key_mem_9__46_,
         top_core_KE_key_mem_9__47_, top_core_KE_key_mem_9__48_,
         top_core_KE_key_mem_9__49_, top_core_KE_key_mem_9__50_,
         top_core_KE_key_mem_9__51_, top_core_KE_key_mem_9__52_,
         top_core_KE_key_mem_9__53_, top_core_KE_key_mem_9__54_,
         top_core_KE_key_mem_9__55_, top_core_KE_key_mem_9__56_,
         top_core_KE_key_mem_9__57_, top_core_KE_key_mem_9__58_,
         top_core_KE_key_mem_9__59_, top_core_KE_key_mem_9__60_,
         top_core_KE_key_mem_9__61_, top_core_KE_key_mem_9__62_,
         top_core_KE_key_mem_9__63_, top_core_KE_key_mem_9__64_,
         top_core_KE_key_mem_9__65_, top_core_KE_key_mem_9__66_,
         top_core_KE_key_mem_9__67_, top_core_KE_key_mem_9__68_,
         top_core_KE_key_mem_9__69_, top_core_KE_key_mem_9__70_,
         top_core_KE_key_mem_9__71_, top_core_KE_key_mem_9__72_,
         top_core_KE_key_mem_9__73_, top_core_KE_key_mem_9__74_,
         top_core_KE_key_mem_9__75_, top_core_KE_key_mem_9__76_,
         top_core_KE_key_mem_9__77_, top_core_KE_key_mem_9__78_,
         top_core_KE_key_mem_9__79_, top_core_KE_key_mem_9__80_,
         top_core_KE_key_mem_9__81_, top_core_KE_key_mem_9__82_,
         top_core_KE_key_mem_9__83_, top_core_KE_key_mem_9__84_,
         top_core_KE_key_mem_9__85_, top_core_KE_key_mem_9__86_,
         top_core_KE_key_mem_9__87_, top_core_KE_key_mem_9__88_,
         top_core_KE_key_mem_9__89_, top_core_KE_key_mem_9__90_,
         top_core_KE_key_mem_9__91_, top_core_KE_key_mem_9__92_,
         top_core_KE_key_mem_9__93_, top_core_KE_key_mem_9__94_,
         top_core_KE_key_mem_9__95_, top_core_KE_key_mem_9__96_,
         top_core_KE_key_mem_9__97_, top_core_KE_key_mem_9__98_,
         top_core_KE_key_mem_9__99_, top_core_KE_key_mem_9__100_,
         top_core_KE_key_mem_9__101_, top_core_KE_key_mem_9__102_,
         top_core_KE_key_mem_9__103_, top_core_KE_key_mem_9__104_,
         top_core_KE_key_mem_9__105_, top_core_KE_key_mem_9__106_,
         top_core_KE_key_mem_9__107_, top_core_KE_key_mem_9__108_,
         top_core_KE_key_mem_9__109_, top_core_KE_key_mem_9__110_,
         top_core_KE_key_mem_9__111_, top_core_KE_key_mem_9__112_,
         top_core_KE_key_mem_9__113_, top_core_KE_key_mem_9__114_,
         top_core_KE_key_mem_9__115_, top_core_KE_key_mem_9__116_,
         top_core_KE_key_mem_9__117_, top_core_KE_key_mem_9__118_,
         top_core_KE_key_mem_9__119_, top_core_KE_key_mem_9__120_,
         top_core_KE_key_mem_9__121_, top_core_KE_key_mem_9__122_,
         top_core_KE_key_mem_9__123_, top_core_KE_key_mem_9__124_,
         top_core_KE_key_mem_9__125_, top_core_KE_key_mem_9__126_,
         top_core_KE_key_mem_9__127_, top_core_KE_key_mem_9__128_,
         top_core_KE_key_mem_8__0_, top_core_KE_key_mem_8__1_,
         top_core_KE_key_mem_8__2_, top_core_KE_key_mem_8__3_,
         top_core_KE_key_mem_8__4_, top_core_KE_key_mem_8__5_,
         top_core_KE_key_mem_8__6_, top_core_KE_key_mem_8__7_,
         top_core_KE_key_mem_8__8_, top_core_KE_key_mem_8__9_,
         top_core_KE_key_mem_8__10_, top_core_KE_key_mem_8__11_,
         top_core_KE_key_mem_8__12_, top_core_KE_key_mem_8__13_,
         top_core_KE_key_mem_8__14_, top_core_KE_key_mem_8__15_,
         top_core_KE_key_mem_8__16_, top_core_KE_key_mem_8__17_,
         top_core_KE_key_mem_8__18_, top_core_KE_key_mem_8__19_,
         top_core_KE_key_mem_8__20_, top_core_KE_key_mem_8__21_,
         top_core_KE_key_mem_8__22_, top_core_KE_key_mem_8__23_,
         top_core_KE_key_mem_8__24_, top_core_KE_key_mem_8__25_,
         top_core_KE_key_mem_8__26_, top_core_KE_key_mem_8__27_,
         top_core_KE_key_mem_8__28_, top_core_KE_key_mem_8__29_,
         top_core_KE_key_mem_8__30_, top_core_KE_key_mem_8__31_,
         top_core_KE_key_mem_8__32_, top_core_KE_key_mem_8__33_,
         top_core_KE_key_mem_8__34_, top_core_KE_key_mem_8__35_,
         top_core_KE_key_mem_8__36_, top_core_KE_key_mem_8__37_,
         top_core_KE_key_mem_8__38_, top_core_KE_key_mem_8__39_,
         top_core_KE_key_mem_8__40_, top_core_KE_key_mem_8__41_,
         top_core_KE_key_mem_8__42_, top_core_KE_key_mem_8__43_,
         top_core_KE_key_mem_8__44_, top_core_KE_key_mem_8__45_,
         top_core_KE_key_mem_8__46_, top_core_KE_key_mem_8__47_,
         top_core_KE_key_mem_8__48_, top_core_KE_key_mem_8__49_,
         top_core_KE_key_mem_8__50_, top_core_KE_key_mem_8__51_,
         top_core_KE_key_mem_8__52_, top_core_KE_key_mem_8__53_,
         top_core_KE_key_mem_8__54_, top_core_KE_key_mem_8__55_,
         top_core_KE_key_mem_8__56_, top_core_KE_key_mem_8__57_,
         top_core_KE_key_mem_8__58_, top_core_KE_key_mem_8__59_,
         top_core_KE_key_mem_8__60_, top_core_KE_key_mem_8__61_,
         top_core_KE_key_mem_8__62_, top_core_KE_key_mem_8__63_,
         top_core_KE_key_mem_8__64_, top_core_KE_key_mem_8__65_,
         top_core_KE_key_mem_8__66_, top_core_KE_key_mem_8__67_,
         top_core_KE_key_mem_8__68_, top_core_KE_key_mem_8__69_,
         top_core_KE_key_mem_8__70_, top_core_KE_key_mem_8__71_,
         top_core_KE_key_mem_8__72_, top_core_KE_key_mem_8__73_,
         top_core_KE_key_mem_8__74_, top_core_KE_key_mem_8__75_,
         top_core_KE_key_mem_8__76_, top_core_KE_key_mem_8__77_,
         top_core_KE_key_mem_8__78_, top_core_KE_key_mem_8__79_,
         top_core_KE_key_mem_8__80_, top_core_KE_key_mem_8__81_,
         top_core_KE_key_mem_8__82_, top_core_KE_key_mem_8__83_,
         top_core_KE_key_mem_8__84_, top_core_KE_key_mem_8__85_,
         top_core_KE_key_mem_8__86_, top_core_KE_key_mem_8__87_,
         top_core_KE_key_mem_8__88_, top_core_KE_key_mem_8__89_,
         top_core_KE_key_mem_8__90_, top_core_KE_key_mem_8__91_,
         top_core_KE_key_mem_8__92_, top_core_KE_key_mem_8__93_,
         top_core_KE_key_mem_8__94_, top_core_KE_key_mem_8__95_,
         top_core_KE_key_mem_8__96_, top_core_KE_key_mem_8__97_,
         top_core_KE_key_mem_8__98_, top_core_KE_key_mem_8__99_,
         top_core_KE_key_mem_8__100_, top_core_KE_key_mem_8__101_,
         top_core_KE_key_mem_8__102_, top_core_KE_key_mem_8__103_,
         top_core_KE_key_mem_8__104_, top_core_KE_key_mem_8__105_,
         top_core_KE_key_mem_8__106_, top_core_KE_key_mem_8__107_,
         top_core_KE_key_mem_8__108_, top_core_KE_key_mem_8__109_,
         top_core_KE_key_mem_8__110_, top_core_KE_key_mem_8__111_,
         top_core_KE_key_mem_8__112_, top_core_KE_key_mem_8__113_,
         top_core_KE_key_mem_8__114_, top_core_KE_key_mem_8__115_,
         top_core_KE_key_mem_8__116_, top_core_KE_key_mem_8__117_,
         top_core_KE_key_mem_8__118_, top_core_KE_key_mem_8__119_,
         top_core_KE_key_mem_8__120_, top_core_KE_key_mem_8__121_,
         top_core_KE_key_mem_8__122_, top_core_KE_key_mem_8__123_,
         top_core_KE_key_mem_8__124_, top_core_KE_key_mem_8__125_,
         top_core_KE_key_mem_8__126_, top_core_KE_key_mem_8__127_,
         top_core_KE_key_mem_8__128_, top_core_KE_key_mem_7__0_,
         top_core_KE_key_mem_7__1_, top_core_KE_key_mem_7__2_,
         top_core_KE_key_mem_7__3_, top_core_KE_key_mem_7__4_,
         top_core_KE_key_mem_7__5_, top_core_KE_key_mem_7__6_,
         top_core_KE_key_mem_7__7_, top_core_KE_key_mem_7__8_,
         top_core_KE_key_mem_7__9_, top_core_KE_key_mem_7__10_,
         top_core_KE_key_mem_7__11_, top_core_KE_key_mem_7__12_,
         top_core_KE_key_mem_7__13_, top_core_KE_key_mem_7__14_,
         top_core_KE_key_mem_7__15_, top_core_KE_key_mem_7__16_,
         top_core_KE_key_mem_7__17_, top_core_KE_key_mem_7__18_,
         top_core_KE_key_mem_7__19_, top_core_KE_key_mem_7__20_,
         top_core_KE_key_mem_7__21_, top_core_KE_key_mem_7__22_,
         top_core_KE_key_mem_7__23_, top_core_KE_key_mem_7__24_,
         top_core_KE_key_mem_7__25_, top_core_KE_key_mem_7__26_,
         top_core_KE_key_mem_7__27_, top_core_KE_key_mem_7__28_,
         top_core_KE_key_mem_7__29_, top_core_KE_key_mem_7__30_,
         top_core_KE_key_mem_7__31_, top_core_KE_key_mem_7__32_,
         top_core_KE_key_mem_7__33_, top_core_KE_key_mem_7__34_,
         top_core_KE_key_mem_7__35_, top_core_KE_key_mem_7__36_,
         top_core_KE_key_mem_7__37_, top_core_KE_key_mem_7__38_,
         top_core_KE_key_mem_7__39_, top_core_KE_key_mem_7__40_,
         top_core_KE_key_mem_7__41_, top_core_KE_key_mem_7__42_,
         top_core_KE_key_mem_7__43_, top_core_KE_key_mem_7__44_,
         top_core_KE_key_mem_7__45_, top_core_KE_key_mem_7__46_,
         top_core_KE_key_mem_7__47_, top_core_KE_key_mem_7__48_,
         top_core_KE_key_mem_7__49_, top_core_KE_key_mem_7__50_,
         top_core_KE_key_mem_7__51_, top_core_KE_key_mem_7__52_,
         top_core_KE_key_mem_7__53_, top_core_KE_key_mem_7__54_,
         top_core_KE_key_mem_7__55_, top_core_KE_key_mem_7__56_,
         top_core_KE_key_mem_7__57_, top_core_KE_key_mem_7__58_,
         top_core_KE_key_mem_7__59_, top_core_KE_key_mem_7__60_,
         top_core_KE_key_mem_7__61_, top_core_KE_key_mem_7__62_,
         top_core_KE_key_mem_7__63_, top_core_KE_key_mem_7__64_,
         top_core_KE_key_mem_7__65_, top_core_KE_key_mem_7__66_,
         top_core_KE_key_mem_7__67_, top_core_KE_key_mem_7__68_,
         top_core_KE_key_mem_7__69_, top_core_KE_key_mem_7__70_,
         top_core_KE_key_mem_7__71_, top_core_KE_key_mem_7__72_,
         top_core_KE_key_mem_7__73_, top_core_KE_key_mem_7__74_,
         top_core_KE_key_mem_7__75_, top_core_KE_key_mem_7__76_,
         top_core_KE_key_mem_7__77_, top_core_KE_key_mem_7__78_,
         top_core_KE_key_mem_7__79_, top_core_KE_key_mem_7__80_,
         top_core_KE_key_mem_7__81_, top_core_KE_key_mem_7__82_,
         top_core_KE_key_mem_7__83_, top_core_KE_key_mem_7__84_,
         top_core_KE_key_mem_7__85_, top_core_KE_key_mem_7__86_,
         top_core_KE_key_mem_7__87_, top_core_KE_key_mem_7__88_,
         top_core_KE_key_mem_7__89_, top_core_KE_key_mem_7__90_,
         top_core_KE_key_mem_7__91_, top_core_KE_key_mem_7__92_,
         top_core_KE_key_mem_7__93_, top_core_KE_key_mem_7__94_,
         top_core_KE_key_mem_7__95_, top_core_KE_key_mem_7__96_,
         top_core_KE_key_mem_7__97_, top_core_KE_key_mem_7__98_,
         top_core_KE_key_mem_7__99_, top_core_KE_key_mem_7__100_,
         top_core_KE_key_mem_7__101_, top_core_KE_key_mem_7__102_,
         top_core_KE_key_mem_7__103_, top_core_KE_key_mem_7__104_,
         top_core_KE_key_mem_7__105_, top_core_KE_key_mem_7__106_,
         top_core_KE_key_mem_7__107_, top_core_KE_key_mem_7__108_,
         top_core_KE_key_mem_7__109_, top_core_KE_key_mem_7__110_,
         top_core_KE_key_mem_7__111_, top_core_KE_key_mem_7__112_,
         top_core_KE_key_mem_7__113_, top_core_KE_key_mem_7__114_,
         top_core_KE_key_mem_7__115_, top_core_KE_key_mem_7__116_,
         top_core_KE_key_mem_7__117_, top_core_KE_key_mem_7__118_,
         top_core_KE_key_mem_7__119_, top_core_KE_key_mem_7__120_,
         top_core_KE_key_mem_7__121_, top_core_KE_key_mem_7__122_,
         top_core_KE_key_mem_7__123_, top_core_KE_key_mem_7__124_,
         top_core_KE_key_mem_7__125_, top_core_KE_key_mem_7__126_,
         top_core_KE_key_mem_7__127_, top_core_KE_key_mem_7__128_,
         top_core_KE_key_mem_6__0_, top_core_KE_key_mem_6__1_,
         top_core_KE_key_mem_6__2_, top_core_KE_key_mem_6__3_,
         top_core_KE_key_mem_6__4_, top_core_KE_key_mem_6__5_,
         top_core_KE_key_mem_6__6_, top_core_KE_key_mem_6__7_,
         top_core_KE_key_mem_6__8_, top_core_KE_key_mem_6__9_,
         top_core_KE_key_mem_6__10_, top_core_KE_key_mem_6__11_,
         top_core_KE_key_mem_6__12_, top_core_KE_key_mem_6__13_,
         top_core_KE_key_mem_6__14_, top_core_KE_key_mem_6__15_,
         top_core_KE_key_mem_6__16_, top_core_KE_key_mem_6__17_,
         top_core_KE_key_mem_6__18_, top_core_KE_key_mem_6__19_,
         top_core_KE_key_mem_6__20_, top_core_KE_key_mem_6__21_,
         top_core_KE_key_mem_6__22_, top_core_KE_key_mem_6__23_,
         top_core_KE_key_mem_6__24_, top_core_KE_key_mem_6__25_,
         top_core_KE_key_mem_6__26_, top_core_KE_key_mem_6__27_,
         top_core_KE_key_mem_6__28_, top_core_KE_key_mem_6__29_,
         top_core_KE_key_mem_6__30_, top_core_KE_key_mem_6__31_,
         top_core_KE_key_mem_6__32_, top_core_KE_key_mem_6__33_,
         top_core_KE_key_mem_6__34_, top_core_KE_key_mem_6__35_,
         top_core_KE_key_mem_6__36_, top_core_KE_key_mem_6__37_,
         top_core_KE_key_mem_6__38_, top_core_KE_key_mem_6__39_,
         top_core_KE_key_mem_6__40_, top_core_KE_key_mem_6__41_,
         top_core_KE_key_mem_6__42_, top_core_KE_key_mem_6__43_,
         top_core_KE_key_mem_6__44_, top_core_KE_key_mem_6__45_,
         top_core_KE_key_mem_6__46_, top_core_KE_key_mem_6__47_,
         top_core_KE_key_mem_6__48_, top_core_KE_key_mem_6__49_,
         top_core_KE_key_mem_6__50_, top_core_KE_key_mem_6__51_,
         top_core_KE_key_mem_6__52_, top_core_KE_key_mem_6__53_,
         top_core_KE_key_mem_6__54_, top_core_KE_key_mem_6__55_,
         top_core_KE_key_mem_6__56_, top_core_KE_key_mem_6__57_,
         top_core_KE_key_mem_6__58_, top_core_KE_key_mem_6__59_,
         top_core_KE_key_mem_6__60_, top_core_KE_key_mem_6__61_,
         top_core_KE_key_mem_6__62_, top_core_KE_key_mem_6__63_,
         top_core_KE_key_mem_6__64_, top_core_KE_key_mem_6__65_,
         top_core_KE_key_mem_6__66_, top_core_KE_key_mem_6__67_,
         top_core_KE_key_mem_6__68_, top_core_KE_key_mem_6__69_,
         top_core_KE_key_mem_6__70_, top_core_KE_key_mem_6__71_,
         top_core_KE_key_mem_6__72_, top_core_KE_key_mem_6__73_,
         top_core_KE_key_mem_6__74_, top_core_KE_key_mem_6__75_,
         top_core_KE_key_mem_6__76_, top_core_KE_key_mem_6__77_,
         top_core_KE_key_mem_6__78_, top_core_KE_key_mem_6__79_,
         top_core_KE_key_mem_6__80_, top_core_KE_key_mem_6__81_,
         top_core_KE_key_mem_6__82_, top_core_KE_key_mem_6__83_,
         top_core_KE_key_mem_6__84_, top_core_KE_key_mem_6__85_,
         top_core_KE_key_mem_6__86_, top_core_KE_key_mem_6__87_,
         top_core_KE_key_mem_6__88_, top_core_KE_key_mem_6__89_,
         top_core_KE_key_mem_6__90_, top_core_KE_key_mem_6__91_,
         top_core_KE_key_mem_6__92_, top_core_KE_key_mem_6__93_,
         top_core_KE_key_mem_6__94_, top_core_KE_key_mem_6__95_,
         top_core_KE_key_mem_6__96_, top_core_KE_key_mem_6__97_,
         top_core_KE_key_mem_6__98_, top_core_KE_key_mem_6__99_,
         top_core_KE_key_mem_6__100_, top_core_KE_key_mem_6__101_,
         top_core_KE_key_mem_6__102_, top_core_KE_key_mem_6__103_,
         top_core_KE_key_mem_6__104_, top_core_KE_key_mem_6__105_,
         top_core_KE_key_mem_6__106_, top_core_KE_key_mem_6__107_,
         top_core_KE_key_mem_6__108_, top_core_KE_key_mem_6__109_,
         top_core_KE_key_mem_6__110_, top_core_KE_key_mem_6__111_,
         top_core_KE_key_mem_6__112_, top_core_KE_key_mem_6__113_,
         top_core_KE_key_mem_6__114_, top_core_KE_key_mem_6__115_,
         top_core_KE_key_mem_6__116_, top_core_KE_key_mem_6__117_,
         top_core_KE_key_mem_6__118_, top_core_KE_key_mem_6__119_,
         top_core_KE_key_mem_6__120_, top_core_KE_key_mem_6__121_,
         top_core_KE_key_mem_6__122_, top_core_KE_key_mem_6__123_,
         top_core_KE_key_mem_6__124_, top_core_KE_key_mem_6__125_,
         top_core_KE_key_mem_6__126_, top_core_KE_key_mem_6__127_,
         top_core_KE_key_mem_6__128_, top_core_KE_key_mem_5__0_,
         top_core_KE_key_mem_5__1_, top_core_KE_key_mem_5__2_,
         top_core_KE_key_mem_5__3_, top_core_KE_key_mem_5__4_,
         top_core_KE_key_mem_5__5_, top_core_KE_key_mem_5__6_,
         top_core_KE_key_mem_5__7_, top_core_KE_key_mem_5__8_,
         top_core_KE_key_mem_5__9_, top_core_KE_key_mem_5__10_,
         top_core_KE_key_mem_5__11_, top_core_KE_key_mem_5__12_,
         top_core_KE_key_mem_5__13_, top_core_KE_key_mem_5__14_,
         top_core_KE_key_mem_5__15_, top_core_KE_key_mem_5__16_,
         top_core_KE_key_mem_5__17_, top_core_KE_key_mem_5__18_,
         top_core_KE_key_mem_5__19_, top_core_KE_key_mem_5__20_,
         top_core_KE_key_mem_5__21_, top_core_KE_key_mem_5__22_,
         top_core_KE_key_mem_5__23_, top_core_KE_key_mem_5__24_,
         top_core_KE_key_mem_5__25_, top_core_KE_key_mem_5__26_,
         top_core_KE_key_mem_5__27_, top_core_KE_key_mem_5__28_,
         top_core_KE_key_mem_5__29_, top_core_KE_key_mem_5__30_,
         top_core_KE_key_mem_5__31_, top_core_KE_key_mem_5__32_,
         top_core_KE_key_mem_5__33_, top_core_KE_key_mem_5__34_,
         top_core_KE_key_mem_5__35_, top_core_KE_key_mem_5__36_,
         top_core_KE_key_mem_5__37_, top_core_KE_key_mem_5__38_,
         top_core_KE_key_mem_5__39_, top_core_KE_key_mem_5__40_,
         top_core_KE_key_mem_5__41_, top_core_KE_key_mem_5__42_,
         top_core_KE_key_mem_5__43_, top_core_KE_key_mem_5__44_,
         top_core_KE_key_mem_5__45_, top_core_KE_key_mem_5__46_,
         top_core_KE_key_mem_5__47_, top_core_KE_key_mem_5__48_,
         top_core_KE_key_mem_5__49_, top_core_KE_key_mem_5__50_,
         top_core_KE_key_mem_5__51_, top_core_KE_key_mem_5__52_,
         top_core_KE_key_mem_5__53_, top_core_KE_key_mem_5__54_,
         top_core_KE_key_mem_5__55_, top_core_KE_key_mem_5__56_,
         top_core_KE_key_mem_5__57_, top_core_KE_key_mem_5__58_,
         top_core_KE_key_mem_5__59_, top_core_KE_key_mem_5__60_,
         top_core_KE_key_mem_5__61_, top_core_KE_key_mem_5__62_,
         top_core_KE_key_mem_5__63_, top_core_KE_key_mem_5__64_,
         top_core_KE_key_mem_5__65_, top_core_KE_key_mem_5__66_,
         top_core_KE_key_mem_5__67_, top_core_KE_key_mem_5__68_,
         top_core_KE_key_mem_5__69_, top_core_KE_key_mem_5__70_,
         top_core_KE_key_mem_5__71_, top_core_KE_key_mem_5__72_,
         top_core_KE_key_mem_5__73_, top_core_KE_key_mem_5__74_,
         top_core_KE_key_mem_5__75_, top_core_KE_key_mem_5__76_,
         top_core_KE_key_mem_5__77_, top_core_KE_key_mem_5__78_,
         top_core_KE_key_mem_5__79_, top_core_KE_key_mem_5__80_,
         top_core_KE_key_mem_5__81_, top_core_KE_key_mem_5__82_,
         top_core_KE_key_mem_5__83_, top_core_KE_key_mem_5__84_,
         top_core_KE_key_mem_5__85_, top_core_KE_key_mem_5__86_,
         top_core_KE_key_mem_5__87_, top_core_KE_key_mem_5__88_,
         top_core_KE_key_mem_5__89_, top_core_KE_key_mem_5__90_,
         top_core_KE_key_mem_5__91_, top_core_KE_key_mem_5__92_,
         top_core_KE_key_mem_5__93_, top_core_KE_key_mem_5__94_,
         top_core_KE_key_mem_5__95_, top_core_KE_key_mem_5__96_,
         top_core_KE_key_mem_5__97_, top_core_KE_key_mem_5__98_,
         top_core_KE_key_mem_5__99_, top_core_KE_key_mem_5__100_,
         top_core_KE_key_mem_5__101_, top_core_KE_key_mem_5__102_,
         top_core_KE_key_mem_5__103_, top_core_KE_key_mem_5__104_,
         top_core_KE_key_mem_5__105_, top_core_KE_key_mem_5__106_,
         top_core_KE_key_mem_5__107_, top_core_KE_key_mem_5__108_,
         top_core_KE_key_mem_5__109_, top_core_KE_key_mem_5__110_,
         top_core_KE_key_mem_5__111_, top_core_KE_key_mem_5__112_,
         top_core_KE_key_mem_5__113_, top_core_KE_key_mem_5__114_,
         top_core_KE_key_mem_5__115_, top_core_KE_key_mem_5__116_,
         top_core_KE_key_mem_5__117_, top_core_KE_key_mem_5__118_,
         top_core_KE_key_mem_5__119_, top_core_KE_key_mem_5__120_,
         top_core_KE_key_mem_5__121_, top_core_KE_key_mem_5__122_,
         top_core_KE_key_mem_5__123_, top_core_KE_key_mem_5__124_,
         top_core_KE_key_mem_5__125_, top_core_KE_key_mem_5__126_,
         top_core_KE_key_mem_5__127_, top_core_KE_key_mem_5__128_,
         top_core_KE_key_mem_4__0_, top_core_KE_key_mem_4__1_,
         top_core_KE_key_mem_4__2_, top_core_KE_key_mem_4__3_,
         top_core_KE_key_mem_4__4_, top_core_KE_key_mem_4__5_,
         top_core_KE_key_mem_4__6_, top_core_KE_key_mem_4__7_,
         top_core_KE_key_mem_4__8_, top_core_KE_key_mem_4__9_,
         top_core_KE_key_mem_4__10_, top_core_KE_key_mem_4__11_,
         top_core_KE_key_mem_4__12_, top_core_KE_key_mem_4__13_,
         top_core_KE_key_mem_4__14_, top_core_KE_key_mem_4__15_,
         top_core_KE_key_mem_4__16_, top_core_KE_key_mem_4__17_,
         top_core_KE_key_mem_4__18_, top_core_KE_key_mem_4__19_,
         top_core_KE_key_mem_4__20_, top_core_KE_key_mem_4__21_,
         top_core_KE_key_mem_4__22_, top_core_KE_key_mem_4__23_,
         top_core_KE_key_mem_4__24_, top_core_KE_key_mem_4__25_,
         top_core_KE_key_mem_4__26_, top_core_KE_key_mem_4__27_,
         top_core_KE_key_mem_4__28_, top_core_KE_key_mem_4__29_,
         top_core_KE_key_mem_4__30_, top_core_KE_key_mem_4__31_,
         top_core_KE_key_mem_4__32_, top_core_KE_key_mem_4__33_,
         top_core_KE_key_mem_4__34_, top_core_KE_key_mem_4__35_,
         top_core_KE_key_mem_4__36_, top_core_KE_key_mem_4__37_,
         top_core_KE_key_mem_4__38_, top_core_KE_key_mem_4__39_,
         top_core_KE_key_mem_4__40_, top_core_KE_key_mem_4__41_,
         top_core_KE_key_mem_4__42_, top_core_KE_key_mem_4__43_,
         top_core_KE_key_mem_4__44_, top_core_KE_key_mem_4__45_,
         top_core_KE_key_mem_4__46_, top_core_KE_key_mem_4__47_,
         top_core_KE_key_mem_4__48_, top_core_KE_key_mem_4__49_,
         top_core_KE_key_mem_4__50_, top_core_KE_key_mem_4__51_,
         top_core_KE_key_mem_4__52_, top_core_KE_key_mem_4__53_,
         top_core_KE_key_mem_4__54_, top_core_KE_key_mem_4__55_,
         top_core_KE_key_mem_4__56_, top_core_KE_key_mem_4__57_,
         top_core_KE_key_mem_4__58_, top_core_KE_key_mem_4__59_,
         top_core_KE_key_mem_4__60_, top_core_KE_key_mem_4__61_,
         top_core_KE_key_mem_4__62_, top_core_KE_key_mem_4__63_,
         top_core_KE_key_mem_4__64_, top_core_KE_key_mem_4__65_,
         top_core_KE_key_mem_4__66_, top_core_KE_key_mem_4__67_,
         top_core_KE_key_mem_4__68_, top_core_KE_key_mem_4__69_,
         top_core_KE_key_mem_4__70_, top_core_KE_key_mem_4__71_,
         top_core_KE_key_mem_4__72_, top_core_KE_key_mem_4__73_,
         top_core_KE_key_mem_4__74_, top_core_KE_key_mem_4__75_,
         top_core_KE_key_mem_4__76_, top_core_KE_key_mem_4__77_,
         top_core_KE_key_mem_4__78_, top_core_KE_key_mem_4__79_,
         top_core_KE_key_mem_4__80_, top_core_KE_key_mem_4__81_,
         top_core_KE_key_mem_4__82_, top_core_KE_key_mem_4__83_,
         top_core_KE_key_mem_4__84_, top_core_KE_key_mem_4__85_,
         top_core_KE_key_mem_4__86_, top_core_KE_key_mem_4__87_,
         top_core_KE_key_mem_4__88_, top_core_KE_key_mem_4__89_,
         top_core_KE_key_mem_4__90_, top_core_KE_key_mem_4__91_,
         top_core_KE_key_mem_4__92_, top_core_KE_key_mem_4__93_,
         top_core_KE_key_mem_4__94_, top_core_KE_key_mem_4__95_,
         top_core_KE_key_mem_4__96_, top_core_KE_key_mem_4__97_,
         top_core_KE_key_mem_4__98_, top_core_KE_key_mem_4__99_,
         top_core_KE_key_mem_4__100_, top_core_KE_key_mem_4__101_,
         top_core_KE_key_mem_4__102_, top_core_KE_key_mem_4__103_,
         top_core_KE_key_mem_4__104_, top_core_KE_key_mem_4__105_,
         top_core_KE_key_mem_4__106_, top_core_KE_key_mem_4__107_,
         top_core_KE_key_mem_4__108_, top_core_KE_key_mem_4__109_,
         top_core_KE_key_mem_4__110_, top_core_KE_key_mem_4__111_,
         top_core_KE_key_mem_4__112_, top_core_KE_key_mem_4__113_,
         top_core_KE_key_mem_4__114_, top_core_KE_key_mem_4__115_,
         top_core_KE_key_mem_4__116_, top_core_KE_key_mem_4__117_,
         top_core_KE_key_mem_4__118_, top_core_KE_key_mem_4__119_,
         top_core_KE_key_mem_4__120_, top_core_KE_key_mem_4__121_,
         top_core_KE_key_mem_4__122_, top_core_KE_key_mem_4__123_,
         top_core_KE_key_mem_4__124_, top_core_KE_key_mem_4__125_,
         top_core_KE_key_mem_4__126_, top_core_KE_key_mem_4__127_,
         top_core_KE_key_mem_4__128_, top_core_KE_key_mem_3__0_,
         top_core_KE_key_mem_3__1_, top_core_KE_key_mem_3__2_,
         top_core_KE_key_mem_3__3_, top_core_KE_key_mem_3__4_,
         top_core_KE_key_mem_3__5_, top_core_KE_key_mem_3__6_,
         top_core_KE_key_mem_3__7_, top_core_KE_key_mem_3__8_,
         top_core_KE_key_mem_3__9_, top_core_KE_key_mem_3__10_,
         top_core_KE_key_mem_3__11_, top_core_KE_key_mem_3__12_,
         top_core_KE_key_mem_3__13_, top_core_KE_key_mem_3__14_,
         top_core_KE_key_mem_3__15_, top_core_KE_key_mem_3__16_,
         top_core_KE_key_mem_3__17_, top_core_KE_key_mem_3__18_,
         top_core_KE_key_mem_3__19_, top_core_KE_key_mem_3__20_,
         top_core_KE_key_mem_3__21_, top_core_KE_key_mem_3__22_,
         top_core_KE_key_mem_3__23_, top_core_KE_key_mem_3__24_,
         top_core_KE_key_mem_3__25_, top_core_KE_key_mem_3__26_,
         top_core_KE_key_mem_3__27_, top_core_KE_key_mem_3__28_,
         top_core_KE_key_mem_3__29_, top_core_KE_key_mem_3__30_,
         top_core_KE_key_mem_3__31_, top_core_KE_key_mem_3__32_,
         top_core_KE_key_mem_3__33_, top_core_KE_key_mem_3__34_,
         top_core_KE_key_mem_3__35_, top_core_KE_key_mem_3__36_,
         top_core_KE_key_mem_3__37_, top_core_KE_key_mem_3__38_,
         top_core_KE_key_mem_3__39_, top_core_KE_key_mem_3__40_,
         top_core_KE_key_mem_3__41_, top_core_KE_key_mem_3__42_,
         top_core_KE_key_mem_3__43_, top_core_KE_key_mem_3__44_,
         top_core_KE_key_mem_3__45_, top_core_KE_key_mem_3__46_,
         top_core_KE_key_mem_3__47_, top_core_KE_key_mem_3__48_,
         top_core_KE_key_mem_3__49_, top_core_KE_key_mem_3__50_,
         top_core_KE_key_mem_3__51_, top_core_KE_key_mem_3__52_,
         top_core_KE_key_mem_3__53_, top_core_KE_key_mem_3__54_,
         top_core_KE_key_mem_3__55_, top_core_KE_key_mem_3__56_,
         top_core_KE_key_mem_3__57_, top_core_KE_key_mem_3__58_,
         top_core_KE_key_mem_3__59_, top_core_KE_key_mem_3__60_,
         top_core_KE_key_mem_3__61_, top_core_KE_key_mem_3__62_,
         top_core_KE_key_mem_3__63_, top_core_KE_key_mem_3__64_,
         top_core_KE_key_mem_3__65_, top_core_KE_key_mem_3__66_,
         top_core_KE_key_mem_3__67_, top_core_KE_key_mem_3__68_,
         top_core_KE_key_mem_3__69_, top_core_KE_key_mem_3__70_,
         top_core_KE_key_mem_3__71_, top_core_KE_key_mem_3__72_,
         top_core_KE_key_mem_3__73_, top_core_KE_key_mem_3__74_,
         top_core_KE_key_mem_3__75_, top_core_KE_key_mem_3__76_,
         top_core_KE_key_mem_3__77_, top_core_KE_key_mem_3__78_,
         top_core_KE_key_mem_3__79_, top_core_KE_key_mem_3__80_,
         top_core_KE_key_mem_3__81_, top_core_KE_key_mem_3__82_,
         top_core_KE_key_mem_3__83_, top_core_KE_key_mem_3__84_,
         top_core_KE_key_mem_3__85_, top_core_KE_key_mem_3__86_,
         top_core_KE_key_mem_3__87_, top_core_KE_key_mem_3__88_,
         top_core_KE_key_mem_3__89_, top_core_KE_key_mem_3__90_,
         top_core_KE_key_mem_3__91_, top_core_KE_key_mem_3__92_,
         top_core_KE_key_mem_3__93_, top_core_KE_key_mem_3__94_,
         top_core_KE_key_mem_3__95_, top_core_KE_key_mem_3__96_,
         top_core_KE_key_mem_3__97_, top_core_KE_key_mem_3__98_,
         top_core_KE_key_mem_3__99_, top_core_KE_key_mem_3__100_,
         top_core_KE_key_mem_3__101_, top_core_KE_key_mem_3__102_,
         top_core_KE_key_mem_3__103_, top_core_KE_key_mem_3__104_,
         top_core_KE_key_mem_3__105_, top_core_KE_key_mem_3__106_,
         top_core_KE_key_mem_3__107_, top_core_KE_key_mem_3__108_,
         top_core_KE_key_mem_3__109_, top_core_KE_key_mem_3__110_,
         top_core_KE_key_mem_3__111_, top_core_KE_key_mem_3__112_,
         top_core_KE_key_mem_3__113_, top_core_KE_key_mem_3__114_,
         top_core_KE_key_mem_3__115_, top_core_KE_key_mem_3__116_,
         top_core_KE_key_mem_3__117_, top_core_KE_key_mem_3__118_,
         top_core_KE_key_mem_3__119_, top_core_KE_key_mem_3__120_,
         top_core_KE_key_mem_3__121_, top_core_KE_key_mem_3__122_,
         top_core_KE_key_mem_3__123_, top_core_KE_key_mem_3__124_,
         top_core_KE_key_mem_3__125_, top_core_KE_key_mem_3__126_,
         top_core_KE_key_mem_3__127_, top_core_KE_key_mem_3__128_,
         top_core_KE_key_mem_2__0_, top_core_KE_key_mem_2__1_,
         top_core_KE_key_mem_2__2_, top_core_KE_key_mem_2__3_,
         top_core_KE_key_mem_2__4_, top_core_KE_key_mem_2__5_,
         top_core_KE_key_mem_2__6_, top_core_KE_key_mem_2__7_,
         top_core_KE_key_mem_2__8_, top_core_KE_key_mem_2__9_,
         top_core_KE_key_mem_2__10_, top_core_KE_key_mem_2__11_,
         top_core_KE_key_mem_2__12_, top_core_KE_key_mem_2__13_,
         top_core_KE_key_mem_2__14_, top_core_KE_key_mem_2__15_,
         top_core_KE_key_mem_2__16_, top_core_KE_key_mem_2__17_,
         top_core_KE_key_mem_2__18_, top_core_KE_key_mem_2__19_,
         top_core_KE_key_mem_2__20_, top_core_KE_key_mem_2__21_,
         top_core_KE_key_mem_2__22_, top_core_KE_key_mem_2__23_,
         top_core_KE_key_mem_2__24_, top_core_KE_key_mem_2__25_,
         top_core_KE_key_mem_2__26_, top_core_KE_key_mem_2__27_,
         top_core_KE_key_mem_2__28_, top_core_KE_key_mem_2__29_,
         top_core_KE_key_mem_2__30_, top_core_KE_key_mem_2__31_,
         top_core_KE_key_mem_2__32_, top_core_KE_key_mem_2__33_,
         top_core_KE_key_mem_2__34_, top_core_KE_key_mem_2__35_,
         top_core_KE_key_mem_2__36_, top_core_KE_key_mem_2__37_,
         top_core_KE_key_mem_2__38_, top_core_KE_key_mem_2__39_,
         top_core_KE_key_mem_2__40_, top_core_KE_key_mem_2__41_,
         top_core_KE_key_mem_2__42_, top_core_KE_key_mem_2__43_,
         top_core_KE_key_mem_2__44_, top_core_KE_key_mem_2__45_,
         top_core_KE_key_mem_2__46_, top_core_KE_key_mem_2__47_,
         top_core_KE_key_mem_2__48_, top_core_KE_key_mem_2__49_,
         top_core_KE_key_mem_2__50_, top_core_KE_key_mem_2__51_,
         top_core_KE_key_mem_2__52_, top_core_KE_key_mem_2__53_,
         top_core_KE_key_mem_2__54_, top_core_KE_key_mem_2__55_,
         top_core_KE_key_mem_2__56_, top_core_KE_key_mem_2__57_,
         top_core_KE_key_mem_2__58_, top_core_KE_key_mem_2__59_,
         top_core_KE_key_mem_2__60_, top_core_KE_key_mem_2__61_,
         top_core_KE_key_mem_2__62_, top_core_KE_key_mem_2__63_,
         top_core_KE_key_mem_2__64_, top_core_KE_key_mem_2__65_,
         top_core_KE_key_mem_2__66_, top_core_KE_key_mem_2__67_,
         top_core_KE_key_mem_2__68_, top_core_KE_key_mem_2__69_,
         top_core_KE_key_mem_2__70_, top_core_KE_key_mem_2__71_,
         top_core_KE_key_mem_2__72_, top_core_KE_key_mem_2__73_,
         top_core_KE_key_mem_2__74_, top_core_KE_key_mem_2__75_,
         top_core_KE_key_mem_2__76_, top_core_KE_key_mem_2__77_,
         top_core_KE_key_mem_2__78_, top_core_KE_key_mem_2__79_,
         top_core_KE_key_mem_2__80_, top_core_KE_key_mem_2__81_,
         top_core_KE_key_mem_2__82_, top_core_KE_key_mem_2__83_,
         top_core_KE_key_mem_2__84_, top_core_KE_key_mem_2__85_,
         top_core_KE_key_mem_2__86_, top_core_KE_key_mem_2__87_,
         top_core_KE_key_mem_2__88_, top_core_KE_key_mem_2__89_,
         top_core_KE_key_mem_2__90_, top_core_KE_key_mem_2__91_,
         top_core_KE_key_mem_2__92_, top_core_KE_key_mem_2__93_,
         top_core_KE_key_mem_2__94_, top_core_KE_key_mem_2__95_,
         top_core_KE_key_mem_2__96_, top_core_KE_key_mem_2__97_,
         top_core_KE_key_mem_2__98_, top_core_KE_key_mem_2__99_,
         top_core_KE_key_mem_2__100_, top_core_KE_key_mem_2__101_,
         top_core_KE_key_mem_2__102_, top_core_KE_key_mem_2__103_,
         top_core_KE_key_mem_2__104_, top_core_KE_key_mem_2__105_,
         top_core_KE_key_mem_2__106_, top_core_KE_key_mem_2__107_,
         top_core_KE_key_mem_2__108_, top_core_KE_key_mem_2__109_,
         top_core_KE_key_mem_2__110_, top_core_KE_key_mem_2__111_,
         top_core_KE_key_mem_2__112_, top_core_KE_key_mem_2__113_,
         top_core_KE_key_mem_2__114_, top_core_KE_key_mem_2__115_,
         top_core_KE_key_mem_2__116_, top_core_KE_key_mem_2__117_,
         top_core_KE_key_mem_2__118_, top_core_KE_key_mem_2__119_,
         top_core_KE_key_mem_2__120_, top_core_KE_key_mem_2__121_,
         top_core_KE_key_mem_2__122_, top_core_KE_key_mem_2__123_,
         top_core_KE_key_mem_2__124_, top_core_KE_key_mem_2__125_,
         top_core_KE_key_mem_2__126_, top_core_KE_key_mem_2__127_,
         top_core_KE_key_mem_2__128_, top_core_KE_key_mem_1__0_,
         top_core_KE_key_mem_1__1_, top_core_KE_key_mem_1__2_,
         top_core_KE_key_mem_1__3_, top_core_KE_key_mem_1__4_,
         top_core_KE_key_mem_1__5_, top_core_KE_key_mem_1__6_,
         top_core_KE_key_mem_1__7_, top_core_KE_key_mem_1__8_,
         top_core_KE_key_mem_1__9_, top_core_KE_key_mem_1__10_,
         top_core_KE_key_mem_1__11_, top_core_KE_key_mem_1__12_,
         top_core_KE_key_mem_1__13_, top_core_KE_key_mem_1__14_,
         top_core_KE_key_mem_1__15_, top_core_KE_key_mem_1__16_,
         top_core_KE_key_mem_1__17_, top_core_KE_key_mem_1__18_,
         top_core_KE_key_mem_1__19_, top_core_KE_key_mem_1__20_,
         top_core_KE_key_mem_1__21_, top_core_KE_key_mem_1__22_,
         top_core_KE_key_mem_1__23_, top_core_KE_key_mem_1__24_,
         top_core_KE_key_mem_1__25_, top_core_KE_key_mem_1__26_,
         top_core_KE_key_mem_1__27_, top_core_KE_key_mem_1__28_,
         top_core_KE_key_mem_1__29_, top_core_KE_key_mem_1__30_,
         top_core_KE_key_mem_1__31_, top_core_KE_key_mem_1__32_,
         top_core_KE_key_mem_1__33_, top_core_KE_key_mem_1__34_,
         top_core_KE_key_mem_1__35_, top_core_KE_key_mem_1__36_,
         top_core_KE_key_mem_1__37_, top_core_KE_key_mem_1__38_,
         top_core_KE_key_mem_1__39_, top_core_KE_key_mem_1__40_,
         top_core_KE_key_mem_1__41_, top_core_KE_key_mem_1__42_,
         top_core_KE_key_mem_1__43_, top_core_KE_key_mem_1__44_,
         top_core_KE_key_mem_1__45_, top_core_KE_key_mem_1__46_,
         top_core_KE_key_mem_1__47_, top_core_KE_key_mem_1__48_,
         top_core_KE_key_mem_1__49_, top_core_KE_key_mem_1__50_,
         top_core_KE_key_mem_1__51_, top_core_KE_key_mem_1__52_,
         top_core_KE_key_mem_1__53_, top_core_KE_key_mem_1__54_,
         top_core_KE_key_mem_1__55_, top_core_KE_key_mem_1__56_,
         top_core_KE_key_mem_1__57_, top_core_KE_key_mem_1__58_,
         top_core_KE_key_mem_1__59_, top_core_KE_key_mem_1__60_,
         top_core_KE_key_mem_1__61_, top_core_KE_key_mem_1__62_,
         top_core_KE_key_mem_1__63_, top_core_KE_key_mem_1__64_,
         top_core_KE_key_mem_1__65_, top_core_KE_key_mem_1__66_,
         top_core_KE_key_mem_1__67_, top_core_KE_key_mem_1__68_,
         top_core_KE_key_mem_1__69_, top_core_KE_key_mem_1__70_,
         top_core_KE_key_mem_1__71_, top_core_KE_key_mem_1__72_,
         top_core_KE_key_mem_1__73_, top_core_KE_key_mem_1__74_,
         top_core_KE_key_mem_1__75_, top_core_KE_key_mem_1__76_,
         top_core_KE_key_mem_1__77_, top_core_KE_key_mem_1__78_,
         top_core_KE_key_mem_1__79_, top_core_KE_key_mem_1__80_,
         top_core_KE_key_mem_1__81_, top_core_KE_key_mem_1__82_,
         top_core_KE_key_mem_1__83_, top_core_KE_key_mem_1__84_,
         top_core_KE_key_mem_1__85_, top_core_KE_key_mem_1__86_,
         top_core_KE_key_mem_1__87_, top_core_KE_key_mem_1__88_,
         top_core_KE_key_mem_1__89_, top_core_KE_key_mem_1__90_,
         top_core_KE_key_mem_1__91_, top_core_KE_key_mem_1__92_,
         top_core_KE_key_mem_1__93_, top_core_KE_key_mem_1__94_,
         top_core_KE_key_mem_1__95_, top_core_KE_key_mem_1__96_,
         top_core_KE_key_mem_1__97_, top_core_KE_key_mem_1__98_,
         top_core_KE_key_mem_1__99_, top_core_KE_key_mem_1__100_,
         top_core_KE_key_mem_1__101_, top_core_KE_key_mem_1__102_,
         top_core_KE_key_mem_1__103_, top_core_KE_key_mem_1__104_,
         top_core_KE_key_mem_1__105_, top_core_KE_key_mem_1__106_,
         top_core_KE_key_mem_1__107_, top_core_KE_key_mem_1__108_,
         top_core_KE_key_mem_1__109_, top_core_KE_key_mem_1__110_,
         top_core_KE_key_mem_1__111_, top_core_KE_key_mem_1__112_,
         top_core_KE_key_mem_1__113_, top_core_KE_key_mem_1__114_,
         top_core_KE_key_mem_1__115_, top_core_KE_key_mem_1__116_,
         top_core_KE_key_mem_1__117_, top_core_KE_key_mem_1__118_,
         top_core_KE_key_mem_1__119_, top_core_KE_key_mem_1__120_,
         top_core_KE_key_mem_1__121_, top_core_KE_key_mem_1__122_,
         top_core_KE_key_mem_1__123_, top_core_KE_key_mem_1__124_,
         top_core_KE_key_mem_1__125_, top_core_KE_key_mem_1__126_,
         top_core_KE_key_mem_1__127_, top_core_KE_key_mem_1__128_,
         top_core_KE_key_mem_0__0_, top_core_KE_key_mem_0__1_,
         top_core_KE_key_mem_0__2_, top_core_KE_key_mem_0__3_,
         top_core_KE_key_mem_0__4_, top_core_KE_key_mem_0__5_,
         top_core_KE_key_mem_0__6_, top_core_KE_key_mem_0__7_,
         top_core_KE_key_mem_0__8_, top_core_KE_key_mem_0__9_,
         top_core_KE_key_mem_0__10_, top_core_KE_key_mem_0__11_,
         top_core_KE_key_mem_0__12_, top_core_KE_key_mem_0__13_,
         top_core_KE_key_mem_0__14_, top_core_KE_key_mem_0__15_,
         top_core_KE_key_mem_0__16_, top_core_KE_key_mem_0__17_,
         top_core_KE_key_mem_0__18_, top_core_KE_key_mem_0__19_,
         top_core_KE_key_mem_0__20_, top_core_KE_key_mem_0__21_,
         top_core_KE_key_mem_0__22_, top_core_KE_key_mem_0__23_,
         top_core_KE_key_mem_0__24_, top_core_KE_key_mem_0__25_,
         top_core_KE_key_mem_0__26_, top_core_KE_key_mem_0__27_,
         top_core_KE_key_mem_0__28_, top_core_KE_key_mem_0__29_,
         top_core_KE_key_mem_0__30_, top_core_KE_key_mem_0__31_,
         top_core_KE_key_mem_0__32_, top_core_KE_key_mem_0__33_,
         top_core_KE_key_mem_0__34_, top_core_KE_key_mem_0__35_,
         top_core_KE_key_mem_0__36_, top_core_KE_key_mem_0__37_,
         top_core_KE_key_mem_0__38_, top_core_KE_key_mem_0__39_,
         top_core_KE_key_mem_0__40_, top_core_KE_key_mem_0__41_,
         top_core_KE_key_mem_0__42_, top_core_KE_key_mem_0__43_,
         top_core_KE_key_mem_0__44_, top_core_KE_key_mem_0__45_,
         top_core_KE_key_mem_0__46_, top_core_KE_key_mem_0__47_,
         top_core_KE_key_mem_0__48_, top_core_KE_key_mem_0__49_,
         top_core_KE_key_mem_0__50_, top_core_KE_key_mem_0__51_,
         top_core_KE_key_mem_0__52_, top_core_KE_key_mem_0__53_,
         top_core_KE_key_mem_0__54_, top_core_KE_key_mem_0__55_,
         top_core_KE_key_mem_0__56_, top_core_KE_key_mem_0__57_,
         top_core_KE_key_mem_0__58_, top_core_KE_key_mem_0__59_,
         top_core_KE_key_mem_0__60_, top_core_KE_key_mem_0__61_,
         top_core_KE_key_mem_0__62_, top_core_KE_key_mem_0__63_,
         top_core_KE_key_mem_0__64_, top_core_KE_key_mem_0__65_,
         top_core_KE_key_mem_0__66_, top_core_KE_key_mem_0__67_,
         top_core_KE_key_mem_0__68_, top_core_KE_key_mem_0__69_,
         top_core_KE_key_mem_0__70_, top_core_KE_key_mem_0__71_,
         top_core_KE_key_mem_0__72_, top_core_KE_key_mem_0__73_,
         top_core_KE_key_mem_0__74_, top_core_KE_key_mem_0__75_,
         top_core_KE_key_mem_0__76_, top_core_KE_key_mem_0__77_,
         top_core_KE_key_mem_0__78_, top_core_KE_key_mem_0__79_,
         top_core_KE_key_mem_0__80_, top_core_KE_key_mem_0__81_,
         top_core_KE_key_mem_0__82_, top_core_KE_key_mem_0__83_,
         top_core_KE_key_mem_0__84_, top_core_KE_key_mem_0__85_,
         top_core_KE_key_mem_0__86_, top_core_KE_key_mem_0__87_,
         top_core_KE_key_mem_0__88_, top_core_KE_key_mem_0__89_,
         top_core_KE_key_mem_0__90_, top_core_KE_key_mem_0__91_,
         top_core_KE_key_mem_0__92_, top_core_KE_key_mem_0__93_,
         top_core_KE_key_mem_0__94_, top_core_KE_key_mem_0__95_,
         top_core_KE_key_mem_0__96_, top_core_KE_key_mem_0__97_,
         top_core_KE_key_mem_0__98_, top_core_KE_key_mem_0__99_,
         top_core_KE_key_mem_0__100_, top_core_KE_key_mem_0__101_,
         top_core_KE_key_mem_0__102_, top_core_KE_key_mem_0__103_,
         top_core_KE_key_mem_0__104_, top_core_KE_key_mem_0__105_,
         top_core_KE_key_mem_0__106_, top_core_KE_key_mem_0__107_,
         top_core_KE_key_mem_0__108_, top_core_KE_key_mem_0__109_,
         top_core_KE_key_mem_0__110_, top_core_KE_key_mem_0__111_,
         top_core_KE_key_mem_0__112_, top_core_KE_key_mem_0__113_,
         top_core_KE_key_mem_0__114_, top_core_KE_key_mem_0__115_,
         top_core_KE_key_mem_0__116_, top_core_KE_key_mem_0__117_,
         top_core_KE_key_mem_0__118_, top_core_KE_key_mem_0__119_,
         top_core_KE_key_mem_0__120_, top_core_KE_key_mem_0__121_,
         top_core_KE_key_mem_0__122_, top_core_KE_key_mem_0__123_,
         top_core_KE_key_mem_0__124_, top_core_KE_key_mem_0__125_,
         top_core_KE_key_mem_0__126_, top_core_KE_key_mem_0__127_,
         top_core_KE_key_mem_0__128_, top_core_KE_Nk0_0_, top_core_KE_Nk0_1_,
         top_core_KE_Nk0_2_, top_core_KE_CipherKey0_0_,
         top_core_KE_CipherKey0_1_, top_core_KE_CipherKey0_2_,
         top_core_KE_CipherKey0_3_, top_core_KE_CipherKey0_4_,
         top_core_KE_CipherKey0_5_, top_core_KE_CipherKey0_6_,
         top_core_KE_CipherKey0_7_, top_core_KE_CipherKey0_8_,
         top_core_KE_CipherKey0_9_, top_core_KE_CipherKey0_10_,
         top_core_KE_CipherKey0_11_, top_core_KE_CipherKey0_12_,
         top_core_KE_CipherKey0_13_, top_core_KE_CipherKey0_14_,
         top_core_KE_CipherKey0_15_, top_core_KE_CipherKey0_16_,
         top_core_KE_CipherKey0_17_, top_core_KE_CipherKey0_18_,
         top_core_KE_CipherKey0_19_, top_core_KE_CipherKey0_20_,
         top_core_KE_CipherKey0_21_, top_core_KE_CipherKey0_22_,
         top_core_KE_CipherKey0_23_, top_core_KE_CipherKey0_24_,
         top_core_KE_CipherKey0_25_, top_core_KE_CipherKey0_26_,
         top_core_KE_CipherKey0_27_, top_core_KE_CipherKey0_28_,
         top_core_KE_CipherKey0_29_, top_core_KE_CipherKey0_30_,
         top_core_KE_CipherKey0_31_, top_core_KE_CipherKey0_32_,
         top_core_KE_CipherKey0_33_, top_core_KE_CipherKey0_34_,
         top_core_KE_CipherKey0_35_, top_core_KE_CipherKey0_36_,
         top_core_KE_CipherKey0_37_, top_core_KE_CipherKey0_38_,
         top_core_KE_CipherKey0_39_, top_core_KE_CipherKey0_40_,
         top_core_KE_CipherKey0_41_, top_core_KE_CipherKey0_42_,
         top_core_KE_CipherKey0_43_, top_core_KE_CipherKey0_44_,
         top_core_KE_CipherKey0_45_, top_core_KE_CipherKey0_46_,
         top_core_KE_CipherKey0_47_, top_core_KE_CipherKey0_48_,
         top_core_KE_CipherKey0_49_, top_core_KE_CipherKey0_50_,
         top_core_KE_CipherKey0_51_, top_core_KE_CipherKey0_52_,
         top_core_KE_CipherKey0_53_, top_core_KE_CipherKey0_54_,
         top_core_KE_CipherKey0_55_, top_core_KE_CipherKey0_56_,
         top_core_KE_CipherKey0_57_, top_core_KE_CipherKey0_58_,
         top_core_KE_CipherKey0_59_, top_core_KE_CipherKey0_60_,
         top_core_KE_CipherKey0_61_, top_core_KE_CipherKey0_62_,
         top_core_KE_CipherKey0_63_, top_core_KE_CipherKey0_64_,
         top_core_KE_CipherKey0_65_, top_core_KE_CipherKey0_66_,
         top_core_KE_CipherKey0_67_, top_core_KE_CipherKey0_68_,
         top_core_KE_CipherKey0_69_, top_core_KE_CipherKey0_70_,
         top_core_KE_CipherKey0_71_, top_core_KE_CipherKey0_72_,
         top_core_KE_CipherKey0_73_, top_core_KE_CipherKey0_74_,
         top_core_KE_CipherKey0_75_, top_core_KE_CipherKey0_76_,
         top_core_KE_CipherKey0_77_, top_core_KE_CipherKey0_78_,
         top_core_KE_CipherKey0_79_, top_core_KE_CipherKey0_80_,
         top_core_KE_CipherKey0_81_, top_core_KE_CipherKey0_82_,
         top_core_KE_CipherKey0_83_, top_core_KE_CipherKey0_84_,
         top_core_KE_CipherKey0_85_, top_core_KE_CipherKey0_86_,
         top_core_KE_CipherKey0_87_, top_core_KE_CipherKey0_88_,
         top_core_KE_CipherKey0_89_, top_core_KE_CipherKey0_90_,
         top_core_KE_CipherKey0_91_, top_core_KE_CipherKey0_92_,
         top_core_KE_CipherKey0_93_, top_core_KE_CipherKey0_94_,
         top_core_KE_CipherKey0_95_, top_core_KE_CipherKey0_96_,
         top_core_KE_CipherKey0_97_, top_core_KE_CipherKey0_98_,
         top_core_KE_CipherKey0_99_, top_core_KE_CipherKey0_100_,
         top_core_KE_CipherKey0_101_, top_core_KE_CipherKey0_102_,
         top_core_KE_CipherKey0_103_, top_core_KE_CipherKey0_104_,
         top_core_KE_CipherKey0_105_, top_core_KE_CipherKey0_106_,
         top_core_KE_CipherKey0_107_, top_core_KE_CipherKey0_108_,
         top_core_KE_CipherKey0_109_, top_core_KE_CipherKey0_110_,
         top_core_KE_CipherKey0_111_, top_core_KE_CipherKey0_112_,
         top_core_KE_CipherKey0_113_, top_core_KE_CipherKey0_114_,
         top_core_KE_CipherKey0_115_, top_core_KE_CipherKey0_116_,
         top_core_KE_CipherKey0_117_, top_core_KE_CipherKey0_118_,
         top_core_KE_CipherKey0_119_, top_core_KE_CipherKey0_120_,
         top_core_KE_CipherKey0_121_, top_core_KE_CipherKey0_122_,
         top_core_KE_CipherKey0_123_, top_core_KE_CipherKey0_124_,
         top_core_KE_CipherKey0_125_, top_core_KE_CipherKey0_126_,
         top_core_KE_CipherKey0_127_, top_core_KE_CipherKey0_128_,
         top_core_KE_CipherKey0_129_, top_core_KE_CipherKey0_130_,
         top_core_KE_CipherKey0_131_, top_core_KE_CipherKey0_132_,
         top_core_KE_CipherKey0_133_, top_core_KE_CipherKey0_134_,
         top_core_KE_CipherKey0_135_, top_core_KE_CipherKey0_136_,
         top_core_KE_CipherKey0_137_, top_core_KE_CipherKey0_138_,
         top_core_KE_CipherKey0_139_, top_core_KE_CipherKey0_140_,
         top_core_KE_CipherKey0_141_, top_core_KE_CipherKey0_142_,
         top_core_KE_CipherKey0_143_, top_core_KE_CipherKey0_144_,
         top_core_KE_CipherKey0_145_, top_core_KE_CipherKey0_146_,
         top_core_KE_CipherKey0_147_, top_core_KE_CipherKey0_148_,
         top_core_KE_CipherKey0_149_, top_core_KE_CipherKey0_150_,
         top_core_KE_CipherKey0_151_, top_core_KE_CipherKey0_152_,
         top_core_KE_CipherKey0_153_, top_core_KE_CipherKey0_154_,
         top_core_KE_CipherKey0_155_, top_core_KE_CipherKey0_156_,
         top_core_KE_CipherKey0_157_, top_core_KE_CipherKey0_158_,
         top_core_KE_CipherKey0_159_, top_core_KE_CipherKey0_160_,
         top_core_KE_CipherKey0_161_, top_core_KE_CipherKey0_162_,
         top_core_KE_CipherKey0_163_, top_core_KE_CipherKey0_164_,
         top_core_KE_CipherKey0_165_, top_core_KE_CipherKey0_166_,
         top_core_KE_CipherKey0_167_, top_core_KE_CipherKey0_168_,
         top_core_KE_CipherKey0_169_, top_core_KE_CipherKey0_170_,
         top_core_KE_CipherKey0_171_, top_core_KE_CipherKey0_172_,
         top_core_KE_CipherKey0_173_, top_core_KE_CipherKey0_174_,
         top_core_KE_CipherKey0_175_, top_core_KE_CipherKey0_176_,
         top_core_KE_CipherKey0_177_, top_core_KE_CipherKey0_178_,
         top_core_KE_CipherKey0_179_, top_core_KE_CipherKey0_180_,
         top_core_KE_CipherKey0_181_, top_core_KE_CipherKey0_182_,
         top_core_KE_CipherKey0_183_, top_core_KE_CipherKey0_184_,
         top_core_KE_CipherKey0_185_, top_core_KE_CipherKey0_186_,
         top_core_KE_CipherKey0_187_, top_core_KE_CipherKey0_188_,
         top_core_KE_CipherKey0_189_, top_core_KE_CipherKey0_190_,
         top_core_KE_CipherKey0_191_, top_core_KE_CipherKey0_192_,
         top_core_KE_CipherKey0_193_, top_core_KE_CipherKey0_194_,
         top_core_KE_CipherKey0_195_, top_core_KE_CipherKey0_196_,
         top_core_KE_CipherKey0_197_, top_core_KE_CipherKey0_198_,
         top_core_KE_CipherKey0_199_, top_core_KE_CipherKey0_200_,
         top_core_KE_CipherKey0_201_, top_core_KE_CipherKey0_202_,
         top_core_KE_CipherKey0_203_, top_core_KE_CipherKey0_204_,
         top_core_KE_CipherKey0_205_, top_core_KE_CipherKey0_206_,
         top_core_KE_CipherKey0_207_, top_core_KE_CipherKey0_208_,
         top_core_KE_CipherKey0_209_, top_core_KE_CipherKey0_210_,
         top_core_KE_CipherKey0_211_, top_core_KE_CipherKey0_212_,
         top_core_KE_CipherKey0_213_, top_core_KE_CipherKey0_214_,
         top_core_KE_CipherKey0_215_, top_core_KE_CipherKey0_216_,
         top_core_KE_CipherKey0_217_, top_core_KE_CipherKey0_218_,
         top_core_KE_CipherKey0_219_, top_core_KE_CipherKey0_220_,
         top_core_KE_CipherKey0_221_, top_core_KE_CipherKey0_222_,
         top_core_KE_CipherKey0_223_, top_core_KE_CipherKey0_224_,
         top_core_KE_CipherKey0_225_, top_core_KE_CipherKey0_226_,
         top_core_KE_CipherKey0_227_, top_core_KE_CipherKey0_228_,
         top_core_KE_CipherKey0_229_, top_core_KE_CipherKey0_230_,
         top_core_KE_CipherKey0_231_, top_core_KE_CipherKey0_232_,
         top_core_KE_CipherKey0_233_, top_core_KE_CipherKey0_234_,
         top_core_KE_CipherKey0_235_, top_core_KE_CipherKey0_236_,
         top_core_KE_CipherKey0_237_, top_core_KE_CipherKey0_238_,
         top_core_KE_CipherKey0_239_, top_core_KE_CipherKey0_240_,
         top_core_KE_CipherKey0_241_, top_core_KE_CipherKey0_242_,
         top_core_KE_CipherKey0_243_, top_core_KE_CipherKey0_244_,
         top_core_KE_CipherKey0_245_, top_core_KE_CipherKey0_246_,
         top_core_KE_CipherKey0_247_, top_core_KE_CipherKey0_248_,
         top_core_KE_CipherKey0_249_, top_core_KE_CipherKey0_250_,
         top_core_KE_CipherKey0_251_, top_core_KE_CipherKey0_252_,
         top_core_KE_CipherKey0_253_, top_core_KE_CipherKey0_254_,
         top_core_KE_CipherKey0_255_, top_core_KE_new_sboxw_192_0_,
         top_core_KE_new_sboxw_192_1_, top_core_KE_new_sboxw_192_2_,
         top_core_KE_new_sboxw_192_3_, top_core_KE_new_sboxw_192_4_,
         top_core_KE_new_sboxw_192_5_, top_core_KE_new_sboxw_192_6_,
         top_core_KE_new_sboxw_192_7_, top_core_KE_new_sboxw_192_8_,
         top_core_KE_new_sboxw_192_9_, top_core_KE_new_sboxw_192_10_,
         top_core_KE_new_sboxw_192_11_, top_core_KE_new_sboxw_192_12_,
         top_core_KE_new_sboxw_192_13_, top_core_KE_new_sboxw_192_14_,
         top_core_KE_new_sboxw_192_15_, top_core_KE_new_sboxw_192_16_,
         top_core_KE_new_sboxw_192_17_, top_core_KE_new_sboxw_192_18_,
         top_core_KE_new_sboxw_192_19_, top_core_KE_new_sboxw_192_20_,
         top_core_KE_new_sboxw_192_21_, top_core_KE_new_sboxw_192_22_,
         top_core_KE_new_sboxw_192_23_, top_core_KE_new_sboxw_192_24_,
         top_core_KE_new_sboxw_192_25_, top_core_KE_new_sboxw_192_26_,
         top_core_KE_new_sboxw_192_27_, top_core_KE_new_sboxw_192_28_,
         top_core_KE_new_sboxw_192_29_, top_core_KE_new_sboxw_192_30_,
         top_core_KE_new_sboxw_192_31_, top_core_KE_new_sboxw_0_,
         top_core_KE_new_sboxw_1_, top_core_KE_new_sboxw_2_,
         top_core_KE_new_sboxw_3_, top_core_KE_new_sboxw_4_,
         top_core_KE_new_sboxw_5_, top_core_KE_new_sboxw_6_,
         top_core_KE_new_sboxw_7_, top_core_KE_new_sboxw_8_,
         top_core_KE_new_sboxw_9_, top_core_KE_new_sboxw_10_,
         top_core_KE_new_sboxw_11_, top_core_KE_new_sboxw_12_,
         top_core_KE_new_sboxw_13_, top_core_KE_new_sboxw_14_,
         top_core_KE_new_sboxw_15_, top_core_KE_new_sboxw_16_,
         top_core_KE_new_sboxw_17_, top_core_KE_new_sboxw_18_,
         top_core_KE_new_sboxw_19_, top_core_KE_new_sboxw_20_,
         top_core_KE_new_sboxw_21_, top_core_KE_new_sboxw_22_,
         top_core_KE_new_sboxw_23_, top_core_KE_new_sboxw_24_,
         top_core_KE_new_sboxw_25_, top_core_KE_new_sboxw_26_,
         top_core_KE_new_sboxw_27_, top_core_KE_new_sboxw_28_,
         top_core_KE_new_sboxw_29_, top_core_KE_new_sboxw_30_,
         top_core_KE_new_sboxw_31_, top_core_io_div_16_n5,
         top_core_io_div_16_n3, top_core_io_div_16_n2, top_core_io_div_16_n1,
         top_core_io_div_16_N8, top_core_io_div_16_N7, top_core_io_div_16_c_1_,
         top_core_io_div_16_c_2_, top_core_EC_ss_n257, top_core_EC_ss_n256,
         top_core_EC_ss_n255, top_core_EC_ss_n254, top_core_EC_ss_n253,
         top_core_EC_ss_n252, top_core_EC_ss_n251, top_core_EC_ss_n250,
         top_core_EC_ss_n249, top_core_EC_ss_n248, top_core_EC_ss_n247,
         top_core_EC_ss_n246, top_core_EC_ss_n245, top_core_EC_ss_n244,
         top_core_EC_ss_n243, top_core_EC_ss_n242, top_core_EC_ss_n241,
         top_core_EC_ss_n240, top_core_EC_ss_n239, top_core_EC_ss_n238,
         top_core_EC_ss_n237, top_core_EC_ss_n236, top_core_EC_ss_n235,
         top_core_EC_ss_n234, top_core_EC_ss_n233, top_core_EC_ss_n232,
         top_core_EC_ss_n231, top_core_EC_ss_n230, top_core_EC_ss_n229,
         top_core_EC_ss_n228, top_core_EC_ss_n227, top_core_EC_ss_n226,
         top_core_EC_ss_n225, top_core_EC_ss_n224, top_core_EC_ss_n223,
         top_core_EC_ss_n222, top_core_EC_ss_n221, top_core_EC_ss_n220,
         top_core_EC_ss_n219, top_core_EC_ss_n218, top_core_EC_ss_n217,
         top_core_EC_ss_n216, top_core_EC_ss_n215, top_core_EC_ss_n214,
         top_core_EC_ss_n213, top_core_EC_ss_n212, top_core_EC_ss_n211,
         top_core_EC_ss_n210, top_core_EC_ss_n209, top_core_EC_ss_n208,
         top_core_EC_ss_n207, top_core_EC_ss_n206, top_core_EC_ss_n205,
         top_core_EC_ss_n204, top_core_EC_ss_n203, top_core_EC_ss_n202,
         top_core_EC_ss_n201, top_core_EC_ss_n200, top_core_EC_ss_n199,
         top_core_EC_ss_n198, top_core_EC_ss_n197, top_core_EC_ss_n196,
         top_core_EC_ss_n195, top_core_EC_ss_n194, top_core_EC_ss_n193,
         top_core_EC_ss_n192, top_core_EC_ss_n191, top_core_EC_ss_n190,
         top_core_EC_ss_n189, top_core_EC_ss_n188, top_core_EC_ss_n187,
         top_core_EC_ss_n186, top_core_EC_ss_n185, top_core_EC_ss_n184,
         top_core_EC_ss_n183, top_core_EC_ss_n182, top_core_EC_ss_n181,
         top_core_EC_ss_n180, top_core_EC_ss_n179, top_core_EC_ss_n178,
         top_core_EC_ss_n177, top_core_EC_ss_n176, top_core_EC_ss_n175,
         top_core_EC_ss_n174, top_core_EC_ss_n173, top_core_EC_ss_n172,
         top_core_EC_ss_n171, top_core_EC_ss_n170, top_core_EC_ss_n169,
         top_core_EC_ss_n168, top_core_EC_ss_n167, top_core_EC_ss_n166,
         top_core_EC_ss_n165, top_core_EC_ss_n164, top_core_EC_ss_n163,
         top_core_EC_ss_n162, top_core_EC_ss_n161, top_core_EC_ss_n160,
         top_core_EC_ss_n159, top_core_EC_ss_n158, top_core_EC_ss_n157,
         top_core_EC_ss_n156, top_core_EC_ss_n155, top_core_EC_ss_n154,
         top_core_EC_ss_n153, top_core_EC_ss_n152, top_core_EC_ss_n151,
         top_core_EC_ss_n150, top_core_EC_ss_n149, top_core_EC_ss_n148,
         top_core_EC_ss_n147, top_core_EC_ss_n146, top_core_EC_ss_n145,
         top_core_EC_ss_n144, top_core_EC_ss_n143, top_core_EC_ss_n142,
         top_core_EC_ss_n141, top_core_EC_ss_n140, top_core_EC_ss_n139,
         top_core_EC_ss_n138, top_core_EC_ss_n137, top_core_EC_ss_n136,
         top_core_EC_ss_n135, top_core_EC_ss_n134, top_core_EC_ss_n133,
         top_core_EC_ss_n132, top_core_EC_ss_n131, top_core_EC_ss_n130,
         top_core_EC_mc_n929, top_core_EC_mc_n928, top_core_EC_mc_n927,
         top_core_EC_mc_n926, top_core_EC_mc_n925, top_core_EC_mc_n924,
         top_core_EC_mc_n923, top_core_EC_mc_n922, top_core_EC_mc_n921,
         top_core_EC_mc_n920, top_core_EC_mc_n919, top_core_EC_mc_n918,
         top_core_EC_mc_n917, top_core_EC_mc_n916, top_core_EC_mc_n915,
         top_core_EC_mc_n914, top_core_EC_mc_n913, top_core_EC_mc_n912,
         top_core_EC_mc_n911, top_core_EC_mc_n910, top_core_EC_mc_n909,
         top_core_EC_mc_n908, top_core_EC_mc_n907, top_core_EC_mc_n906,
         top_core_EC_mc_n905, top_core_EC_mc_n904, top_core_EC_mc_n903,
         top_core_EC_mc_n902, top_core_EC_mc_n901, top_core_EC_mc_n900,
         top_core_EC_mc_n899, top_core_EC_mc_n898, top_core_EC_mc_n897,
         top_core_EC_mc_n896, top_core_EC_mc_n895, top_core_EC_mc_n894,
         top_core_EC_mc_n893, top_core_EC_mc_n892, top_core_EC_mc_n891,
         top_core_EC_mc_n890, top_core_EC_mc_n889, top_core_EC_mc_n888,
         top_core_EC_mc_n887, top_core_EC_mc_n886, top_core_EC_mc_n885,
         top_core_EC_mc_n884, top_core_EC_mc_n883, top_core_EC_mc_n882,
         top_core_EC_mc_n881, top_core_EC_mc_n880, top_core_EC_mc_n879,
         top_core_EC_mc_n878, top_core_EC_mc_n877, top_core_EC_mc_n876,
         top_core_EC_mc_n875, top_core_EC_mc_n874, top_core_EC_mc_n873,
         top_core_EC_mc_n872, top_core_EC_mc_n871, top_core_EC_mc_n870,
         top_core_EC_mc_n869, top_core_EC_mc_n868, top_core_EC_mc_n867,
         top_core_EC_mc_n866, top_core_EC_mc_n865, top_core_EC_mc_n864,
         top_core_EC_mc_n863, top_core_EC_mc_n862, top_core_EC_mc_n861,
         top_core_EC_mc_n860, top_core_EC_mc_n859, top_core_EC_mc_n858,
         top_core_EC_mc_n857, top_core_EC_mc_n856, top_core_EC_mc_n855,
         top_core_EC_mc_n854, top_core_EC_mc_n853, top_core_EC_mc_n852,
         top_core_EC_mc_n851, top_core_EC_mc_n850, top_core_EC_mc_n849,
         top_core_EC_mc_n848, top_core_EC_mc_n847, top_core_EC_mc_n846,
         top_core_EC_mc_n845, top_core_EC_mc_n844, top_core_EC_mc_n843,
         top_core_EC_mc_n842, top_core_EC_mc_n841, top_core_EC_mc_n840,
         top_core_EC_mc_n839, top_core_EC_mc_n838, top_core_EC_mc_n837,
         top_core_EC_mc_n836, top_core_EC_mc_n835, top_core_EC_mc_n834,
         top_core_EC_mc_n833, top_core_EC_mc_n832, top_core_EC_mc_n831,
         top_core_EC_mc_n830, top_core_EC_mc_n829, top_core_EC_mc_n828,
         top_core_EC_mc_n827, top_core_EC_mc_n826, top_core_EC_mc_n825,
         top_core_EC_mc_n824, top_core_EC_mc_n823, top_core_EC_mc_n822,
         top_core_EC_mc_n821, top_core_EC_mc_n820, top_core_EC_mc_n819,
         top_core_EC_mc_n818, top_core_EC_mc_n817, top_core_EC_mc_n816,
         top_core_EC_mc_n815, top_core_EC_mc_n814, top_core_EC_mc_n813,
         top_core_EC_mc_n812, top_core_EC_mc_n811, top_core_EC_mc_n810,
         top_core_EC_mc_n809, top_core_EC_mc_n808, top_core_EC_mc_n807,
         top_core_EC_mc_n806, top_core_EC_mc_n805, top_core_EC_mc_n804,
         top_core_EC_mc_n803, top_core_EC_mc_n802, top_core_EC_mc_n801,
         top_core_EC_mc_n800, top_core_EC_mc_n799, top_core_EC_mc_n798,
         top_core_EC_mc_n797, top_core_EC_mc_n796, top_core_EC_mc_n795,
         top_core_EC_mc_n794, top_core_EC_mc_n793, top_core_EC_mc_n792,
         top_core_EC_mc_n791, top_core_EC_mc_n790, top_core_EC_mc_n789,
         top_core_EC_mc_n788, top_core_EC_mc_n787, top_core_EC_mc_n786,
         top_core_EC_mc_n785, top_core_EC_mc_n784, top_core_EC_mc_n783,
         top_core_EC_mc_n782, top_core_EC_mc_n781, top_core_EC_mc_n780,
         top_core_EC_mc_n779, top_core_EC_mc_n778, top_core_EC_mc_n777,
         top_core_EC_mc_n776, top_core_EC_mc_n775, top_core_EC_mc_n774,
         top_core_EC_mc_n773, top_core_EC_mc_n772, top_core_EC_mc_n771,
         top_core_EC_mc_n770, top_core_EC_mc_n769, top_core_EC_mc_n768,
         top_core_EC_mc_n767, top_core_EC_mc_n766, top_core_EC_mc_n765,
         top_core_EC_mc_n764, top_core_EC_mc_n763, top_core_EC_mc_n762,
         top_core_EC_mc_n761, top_core_EC_mc_n760, top_core_EC_mc_n759,
         top_core_EC_mc_n758, top_core_EC_mc_n757, top_core_EC_mc_n756,
         top_core_EC_mc_n755, top_core_EC_mc_n754, top_core_EC_mc_n753,
         top_core_EC_mc_n752, top_core_EC_mc_n751, top_core_EC_mc_n750,
         top_core_EC_mc_n749, top_core_EC_mc_n748, top_core_EC_mc_n747,
         top_core_EC_mc_n746, top_core_EC_mc_n745, top_core_EC_mc_n744,
         top_core_EC_mc_n743, top_core_EC_mc_n742, top_core_EC_mc_n741,
         top_core_EC_mc_n740, top_core_EC_mc_n739, top_core_EC_mc_n738,
         top_core_EC_mc_n737, top_core_EC_mc_n736, top_core_EC_mc_n735,
         top_core_EC_mc_n734, top_core_EC_mc_n733, top_core_EC_mc_n732,
         top_core_EC_mc_n731, top_core_EC_mc_n730, top_core_EC_mc_n729,
         top_core_EC_mc_n728, top_core_EC_mc_n727, top_core_EC_mc_n726,
         top_core_EC_mc_n725, top_core_EC_mc_n724, top_core_EC_mc_n723,
         top_core_EC_mc_n722, top_core_EC_mc_n721, top_core_EC_mc_n720,
         top_core_EC_mc_n719, top_core_EC_mc_n718, top_core_EC_mc_n717,
         top_core_EC_mc_n716, top_core_EC_mc_n715, top_core_EC_mc_n714,
         top_core_EC_mc_n713, top_core_EC_mc_n712, top_core_EC_mc_n711,
         top_core_EC_mc_n710, top_core_EC_mc_n709, top_core_EC_mc_n708,
         top_core_EC_mc_n707, top_core_EC_mc_n706, top_core_EC_mc_n705,
         top_core_EC_mc_n704, top_core_EC_mc_n703, top_core_EC_mc_n702,
         top_core_EC_mc_n701, top_core_EC_mc_n700, top_core_EC_mc_n699,
         top_core_EC_mc_n698, top_core_EC_mc_n697, top_core_EC_mc_n696,
         top_core_EC_mc_n695, top_core_EC_mc_n694, top_core_EC_mc_n693,
         top_core_EC_mc_n692, top_core_EC_mc_n691, top_core_EC_mc_n690,
         top_core_EC_mc_n689, top_core_EC_mc_n688, top_core_EC_mc_n687,
         top_core_EC_mc_n686, top_core_EC_mc_n685, top_core_EC_mc_n684,
         top_core_EC_mc_n683, top_core_EC_mc_n682, top_core_EC_mc_n681,
         top_core_EC_mc_n680, top_core_EC_mc_n679, top_core_EC_mc_n678,
         top_core_EC_mc_n677, top_core_EC_mc_n676, top_core_EC_mc_n675,
         top_core_EC_mc_n674, top_core_EC_mc_n673, top_core_EC_mc_n672,
         top_core_EC_mc_n671, top_core_EC_mc_n670, top_core_EC_mc_n669,
         top_core_EC_mc_n668, top_core_EC_mc_n667, top_core_EC_mc_n666,
         top_core_EC_mc_n665, top_core_EC_mc_n664, top_core_EC_mc_n663,
         top_core_EC_mc_n662, top_core_EC_mc_n661, top_core_EC_mc_n660,
         top_core_EC_mc_n659, top_core_EC_mc_n658, top_core_EC_mc_n657,
         top_core_EC_mc_n656, top_core_EC_mc_n655, top_core_EC_mc_n654,
         top_core_EC_mc_n653, top_core_EC_mc_n652, top_core_EC_mc_n651,
         top_core_EC_mc_n650, top_core_EC_mc_n649, top_core_EC_mc_n648,
         top_core_EC_mc_n647, top_core_EC_mc_n646, top_core_EC_mc_n645,
         top_core_EC_mc_n644, top_core_EC_mc_n643, top_core_EC_mc_n642,
         top_core_EC_mc_n641, top_core_EC_mc_n640, top_core_EC_mc_n639,
         top_core_EC_mc_n638, top_core_EC_mc_n637, top_core_EC_mc_n636,
         top_core_EC_mc_n635, top_core_EC_mc_n634, top_core_EC_mc_n633,
         top_core_EC_mc_n632, top_core_EC_mc_n631, top_core_EC_mc_n630,
         top_core_EC_mc_n629, top_core_EC_mc_n628, top_core_EC_mc_n627,
         top_core_EC_mc_n626, top_core_EC_mc_n625, top_core_EC_mc_n624,
         top_core_EC_mc_n623, top_core_EC_mc_n622, top_core_EC_mc_n621,
         top_core_EC_mc_n620, top_core_EC_mc_n619, top_core_EC_mc_n618,
         top_core_EC_mc_n617, top_core_EC_mc_n616, top_core_EC_mc_n615,
         top_core_EC_mc_n614, top_core_EC_mc_n613, top_core_EC_mc_n612,
         top_core_EC_mc_n611, top_core_EC_mc_n610, top_core_EC_mc_n609,
         top_core_EC_mc_n608, top_core_EC_mc_n607, top_core_EC_mc_n606,
         top_core_EC_mc_n605, top_core_EC_mc_n604, top_core_EC_mc_n603,
         top_core_EC_mc_n602, top_core_EC_mc_n601, top_core_EC_mc_n600,
         top_core_EC_mc_n599, top_core_EC_mc_n598, top_core_EC_mc_n597,
         top_core_EC_mc_n596, top_core_EC_mc_n595, top_core_EC_mc_n594,
         top_core_EC_mc_n593, top_core_EC_mc_n592, top_core_EC_mc_n591,
         top_core_EC_mc_n590, top_core_EC_mc_n589, top_core_EC_mc_n588,
         top_core_EC_mc_n587, top_core_EC_mc_n586, top_core_EC_mc_n585,
         top_core_EC_mc_n584, top_core_EC_mc_n583, top_core_EC_mc_n582,
         top_core_EC_mc_n581, top_core_EC_mc_n580, top_core_EC_mc_n579,
         top_core_EC_mc_n578, top_core_EC_mc_n577, top_core_EC_mc_n576,
         top_core_EC_mc_n575, top_core_EC_mc_n574, top_core_EC_mc_n573,
         top_core_EC_mc_n572, top_core_EC_mc_n571, top_core_EC_mc_n570,
         top_core_EC_mc_n569, top_core_EC_mc_n568, top_core_EC_mc_n567,
         top_core_EC_mc_n566, top_core_EC_mc_n565, top_core_EC_mc_n564,
         top_core_EC_mc_n563, top_core_EC_mc_n562, top_core_EC_mc_n561,
         top_core_EC_mc_n560, top_core_EC_mc_n559, top_core_EC_mc_n558,
         top_core_EC_mc_n557, top_core_EC_mc_n556, top_core_EC_mc_n555,
         top_core_EC_mc_n554, top_core_EC_mc_n553, top_core_EC_mc_n552,
         top_core_EC_mc_n551, top_core_EC_mc_n550, top_core_EC_mc_n549,
         top_core_EC_mc_n548, top_core_EC_mc_n547, top_core_EC_mc_n546,
         top_core_EC_mc_n545, top_core_EC_mc_n544, top_core_EC_mc_n543,
         top_core_EC_mc_n542, top_core_EC_mc_n541, top_core_EC_mc_n540,
         top_core_EC_mc_n539, top_core_EC_mc_n538, top_core_EC_mc_n537,
         top_core_EC_mc_n536, top_core_EC_mc_n535, top_core_EC_mc_n534,
         top_core_EC_mc_n533, top_core_EC_mc_n532, top_core_EC_mc_n531,
         top_core_EC_mc_n530, top_core_EC_mc_n529, top_core_EC_mc_n528,
         top_core_EC_mc_n527, top_core_EC_mc_n526, top_core_EC_mc_n525,
         top_core_EC_mc_n524, top_core_EC_mc_n523, top_core_EC_mc_n522,
         top_core_EC_mc_n521, top_core_EC_mc_n520, top_core_EC_mc_n519,
         top_core_EC_mc_n518, top_core_EC_mc_n517, top_core_EC_mc_n516,
         top_core_EC_mc_n515, top_core_EC_mc_n514, top_core_EC_mc_n513,
         top_core_EC_mc_n512, top_core_EC_mc_n511, top_core_EC_mc_n510,
         top_core_EC_mc_n509, top_core_EC_mc_n508, top_core_EC_mc_n507,
         top_core_EC_mc_n506, top_core_EC_mc_n505, top_core_EC_mc_n504,
         top_core_EC_mc_n503, top_core_EC_mc_n502, top_core_EC_mc_n501,
         top_core_EC_mc_n500, top_core_EC_mc_n499, top_core_EC_mc_n498,
         top_core_EC_mc_n497, top_core_EC_mc_n496, top_core_EC_mc_n495,
         top_core_EC_mc_n494, top_core_EC_mc_n493, top_core_EC_mc_n492,
         top_core_EC_mc_n491, top_core_EC_mc_n490, top_core_EC_mc_n489,
         top_core_EC_mc_n488, top_core_EC_mc_n487, top_core_EC_mc_n486,
         top_core_EC_mc_n485, top_core_EC_mc_n484, top_core_EC_mc_n483,
         top_core_EC_mc_n482, top_core_EC_mc_n481, top_core_EC_mc_n480,
         top_core_EC_mc_n479, top_core_EC_mc_n478, top_core_EC_mc_n477,
         top_core_EC_mc_n476, top_core_EC_mc_n475, top_core_EC_mc_n474,
         top_core_EC_mc_n473, top_core_EC_mc_n472, top_core_EC_mc_n471,
         top_core_EC_mc_n470, top_core_EC_mc_n469, top_core_EC_mc_n468,
         top_core_EC_mc_n467, top_core_EC_mc_n466, top_core_EC_mc_n465,
         top_core_EC_mc_n464, top_core_EC_mc_n463, top_core_EC_mc_n462,
         top_core_EC_mc_n461, top_core_EC_mc_n460, top_core_EC_mc_n459,
         top_core_EC_mc_n458, top_core_EC_mc_n457, top_core_EC_mc_n456,
         top_core_EC_mc_n455, top_core_EC_mc_n454, top_core_EC_mc_n453,
         top_core_EC_mc_n452, top_core_EC_mc_n451, top_core_EC_mc_n450,
         top_core_EC_mc_n449, top_core_EC_mc_n448, top_core_EC_mc_n447,
         top_core_EC_mc_n446, top_core_EC_mc_n445, top_core_EC_mc_n444,
         top_core_EC_mc_n443, top_core_EC_mc_n442, top_core_EC_mc_n441,
         top_core_EC_mc_n440, top_core_EC_mc_n439, top_core_EC_mc_n438,
         top_core_EC_mc_n437, top_core_EC_mc_n436, top_core_EC_mc_n435,
         top_core_EC_mc_n434, top_core_EC_mc_n433, top_core_EC_mc_n432,
         top_core_EC_mc_n431, top_core_EC_mc_n430, top_core_EC_mc_n429,
         top_core_EC_mc_n428, top_core_EC_mc_n427, top_core_EC_mc_n426,
         top_core_EC_mc_n425, top_core_EC_mc_n424, top_core_EC_mc_n423,
         top_core_EC_mc_n422, top_core_EC_mc_n421, top_core_EC_mc_n420,
         top_core_EC_mc_n419, top_core_EC_mc_n418, top_core_EC_mc_n417,
         top_core_EC_mc_n416, top_core_EC_mc_n415, top_core_EC_mc_n414,
         top_core_EC_mc_n413, top_core_EC_mc_n412, top_core_EC_mc_n411,
         top_core_EC_mc_n410, top_core_EC_mc_n409, top_core_EC_mc_n408,
         top_core_EC_mc_n407, top_core_EC_mc_n406, top_core_EC_mc_n405,
         top_core_EC_mc_n404, top_core_EC_mc_n403, top_core_EC_mc_n402,
         top_core_EC_mc_n401, top_core_EC_mc_n400, top_core_EC_mc_n399,
         top_core_EC_mc_n398, top_core_EC_mc_n397, top_core_EC_mc_n396,
         top_core_EC_mc_n395, top_core_EC_mc_n394, top_core_EC_mc_n393,
         top_core_EC_mc_n392, top_core_EC_mc_n391, top_core_EC_mc_n390,
         top_core_EC_mc_n389, top_core_EC_mc_n388, top_core_EC_mc_n387,
         top_core_EC_mc_n386, top_core_EC_mc_n385, top_core_EC_mc_n384,
         top_core_EC_mc_n383, top_core_EC_mc_n382, top_core_EC_mc_n381,
         top_core_EC_mc_n380, top_core_EC_mc_n379, top_core_EC_mc_n378,
         top_core_EC_mc_n377, top_core_EC_mc_n376, top_core_EC_mc_n375,
         top_core_EC_mc_n374, top_core_EC_mc_n373, top_core_EC_mc_n372,
         top_core_EC_mc_n371, top_core_EC_mc_n370, top_core_EC_mc_n369,
         top_core_EC_mc_n368, top_core_EC_mc_n367, top_core_EC_mc_n366,
         top_core_EC_mc_n365, top_core_EC_mc_n364, top_core_EC_mc_n363,
         top_core_EC_mc_n362, top_core_EC_mc_n361, top_core_EC_mc_n360,
         top_core_EC_mc_n359, top_core_EC_mc_n358, top_core_EC_mc_n357,
         top_core_EC_mc_n356, top_core_EC_mc_n355, top_core_EC_mc_n354,
         top_core_EC_mc_n353, top_core_EC_mc_n352, top_core_EC_mc_n351,
         top_core_EC_mc_n350, top_core_EC_mc_n349, top_core_EC_mc_n348,
         top_core_EC_mc_n347, top_core_EC_mc_n346, top_core_EC_mc_n345,
         top_core_EC_mc_n344, top_core_EC_mc_n343, top_core_EC_mc_n342,
         top_core_EC_mc_n341, top_core_EC_mc_n340, top_core_EC_mc_n339,
         top_core_EC_mc_n338, top_core_EC_mc_n337, top_core_EC_mc_n336,
         top_core_EC_mc_n335, top_core_EC_mc_n334, top_core_EC_mc_n333,
         top_core_EC_mc_n332, top_core_EC_mc_n331, top_core_EC_mc_n330,
         top_core_EC_mc_n329, top_core_EC_mc_n328, top_core_EC_mc_n327,
         top_core_EC_mc_n326, top_core_EC_mc_n325, top_core_EC_mc_n324,
         top_core_EC_mc_n323, top_core_EC_mc_n322, top_core_EC_mc_n321,
         top_core_EC_mc_n320, top_core_EC_mc_n319, top_core_EC_mc_n318,
         top_core_EC_mc_n317, top_core_EC_mc_n316, top_core_EC_mc_n315,
         top_core_EC_mc_n314, top_core_EC_mc_n313, top_core_EC_mc_n312,
         top_core_EC_mc_n311, top_core_EC_mc_n310, top_core_EC_mc_n309,
         top_core_EC_mc_n308, top_core_EC_mc_n307, top_core_EC_mc_n306,
         top_core_EC_mc_n305, top_core_EC_mc_n304, top_core_EC_mc_n303,
         top_core_EC_mc_n302, top_core_EC_mc_n301, top_core_EC_mc_n300,
         top_core_EC_mc_n299, top_core_EC_mc_n298, top_core_EC_mc_n297,
         top_core_EC_mc_n296, top_core_EC_mc_n295, top_core_EC_mc_n294,
         top_core_EC_mc_n293, top_core_EC_mc_n292, top_core_EC_mc_n291,
         top_core_EC_mc_n290, top_core_EC_mc_n289, top_core_EC_mc_n288,
         top_core_EC_mc_n287, top_core_EC_mc_n286, top_core_EC_mc_n285,
         top_core_EC_mc_n284, top_core_EC_mc_n283, top_core_EC_mc_n282,
         top_core_EC_mc_n281, top_core_EC_mc_n280, top_core_EC_mc_n279,
         top_core_EC_mc_n278, top_core_EC_mc_n277, top_core_EC_mc_n276,
         top_core_EC_mc_n275, top_core_EC_mc_n274, top_core_EC_mc_n273,
         top_core_EC_mc_n272, top_core_EC_mc_n271, top_core_EC_mc_n270,
         top_core_EC_mc_n269, top_core_EC_mc_n268, top_core_EC_mc_n267,
         top_core_EC_mc_n266, top_core_EC_mc_n265, top_core_EC_mc_n264,
         top_core_EC_mc_n263, top_core_EC_mc_n262, top_core_EC_mc_n261,
         top_core_EC_mc_n260, top_core_EC_mc_n259, top_core_EC_mc_n258,
         top_core_EC_mc_n257, top_core_EC_mc_n256, top_core_EC_mc_n255,
         top_core_EC_mc_n254, top_core_EC_mc_n253, top_core_EC_mc_n252,
         top_core_EC_mc_n251, top_core_EC_mc_n250, top_core_EC_mc_n249,
         top_core_EC_mc_n248, top_core_EC_mc_n247, top_core_EC_mc_n246,
         top_core_EC_mc_n245, top_core_EC_mc_n244, top_core_EC_mc_n243,
         top_core_EC_mc_n242, top_core_EC_mc_n241, top_core_EC_mc_n240,
         top_core_EC_mc_n239, top_core_EC_mc_n238, top_core_EC_mc_n237,
         top_core_EC_mc_n236, top_core_EC_mc_n235, top_core_EC_mc_n234,
         top_core_EC_mc_n233, top_core_EC_mc_n232, top_core_EC_mc_n231,
         top_core_EC_mc_n230, top_core_EC_mc_n229, top_core_EC_mc_n228,
         top_core_EC_mc_n227, top_core_EC_mc_n226, top_core_EC_mc_n225,
         top_core_EC_mc_n224, top_core_EC_mc_n223, top_core_EC_mc_n222,
         top_core_EC_mc_n221, top_core_EC_mc_n220, top_core_EC_mc_n219,
         top_core_EC_mc_n218, top_core_EC_mc_n217, top_core_EC_mc_n216,
         top_core_EC_mc_n215, top_core_EC_mc_n214, top_core_EC_mc_n213,
         top_core_EC_mc_n212, top_core_EC_mc_n211, top_core_EC_mc_n210,
         top_core_EC_mc_n209, top_core_EC_mc_n208, top_core_EC_mc_n207,
         top_core_EC_mc_n206, top_core_EC_mc_n205, top_core_EC_mc_n204,
         top_core_EC_mc_n203, top_core_EC_mc_n202, top_core_EC_mc_n201,
         top_core_EC_mc_n200, top_core_EC_mc_n199, top_core_EC_mc_n198,
         top_core_EC_mc_n197, top_core_EC_mc_n196, top_core_EC_mc_n195,
         top_core_EC_mc_n194, top_core_EC_mc_n193, top_core_EC_mc_n192,
         top_core_EC_mc_n191, top_core_EC_mc_n190, top_core_EC_mc_n189,
         top_core_EC_mc_n188, top_core_EC_mc_n187, top_core_EC_mc_n186,
         top_core_EC_mc_n185, top_core_EC_mc_n184, top_core_EC_mc_n183,
         top_core_EC_mc_n182, top_core_EC_mc_n181, top_core_EC_mc_n180,
         top_core_EC_mc_n179, top_core_EC_mc_n178, top_core_EC_mc_n177,
         top_core_EC_mc_n176, top_core_EC_mc_n175, top_core_EC_mc_n174,
         top_core_EC_mc_n173, top_core_EC_mc_n172, top_core_EC_mc_n171,
         top_core_EC_mc_n170, top_core_EC_mc_n169, top_core_EC_mc_n168,
         top_core_EC_mc_n167, top_core_EC_mc_n166, top_core_EC_mc_n165,
         top_core_EC_mc_n164, top_core_EC_mc_n163, top_core_EC_mc_n162,
         top_core_EC_mc_n161, top_core_EC_mc_n160, top_core_EC_mc_n159,
         top_core_EC_mc_n158, top_core_EC_mc_n157, top_core_EC_mc_n156,
         top_core_EC_mc_n155, top_core_EC_mc_n154, top_core_EC_mc_n153,
         top_core_EC_mc_n152, top_core_EC_mc_n151, top_core_EC_mc_n150,
         top_core_EC_mc_n149, top_core_EC_mc_n148, top_core_EC_mc_n147,
         top_core_EC_mc_n146, top_core_EC_mc_n145, top_core_EC_mc_n144,
         top_core_EC_mc_n143, top_core_EC_mc_n142, top_core_EC_mc_n141,
         top_core_EC_mc_n140, top_core_EC_mc_n139, top_core_EC_mc_n138,
         top_core_EC_mc_n137, top_core_EC_mc_n136, top_core_EC_mc_n135,
         top_core_EC_mc_n134, top_core_EC_mc_n133, top_core_EC_mc_n132,
         top_core_EC_mc_n131, top_core_EC_mc_n130, top_core_EC_mc_n129,
         top_core_EC_mc_n128, top_core_EC_mc_n127, top_core_EC_mc_n126,
         top_core_EC_mc_n125, top_core_EC_mc_n124, top_core_EC_mc_n123,
         top_core_EC_mc_n122, top_core_EC_mc_n121, top_core_EC_mc_n120,
         top_core_EC_mc_n119, top_core_EC_mc_n118, top_core_EC_mc_n117,
         top_core_EC_mc_n116, top_core_EC_mc_n115, top_core_EC_mc_n114,
         top_core_EC_mc_n113, top_core_EC_mc_n112, top_core_EC_mc_n111,
         top_core_EC_mc_n110, top_core_EC_mc_n109, top_core_EC_mc_n108,
         top_core_EC_mc_n107, top_core_EC_mc_n106, top_core_EC_mc_n105,
         top_core_EC_mc_n104, top_core_EC_mc_n103, top_core_EC_mc_n102,
         top_core_EC_mc_n101, top_core_EC_mc_n100, top_core_EC_mc_n99,
         top_core_EC_mc_n98, top_core_EC_mc_n97, top_core_EC_mc_n96,
         top_core_EC_mc_n95, top_core_EC_mc_n94, top_core_EC_mc_n93,
         top_core_EC_mc_n92, top_core_EC_mc_n91, top_core_EC_mc_n90,
         top_core_EC_mc_n89, top_core_EC_mc_n88, top_core_EC_mc_n87,
         top_core_EC_mc_n86, top_core_EC_mc_n85, top_core_EC_mc_n84,
         top_core_EC_mc_n83, top_core_EC_mc_n82, top_core_EC_mc_n81,
         top_core_EC_mc_n80, top_core_EC_mc_n79, top_core_EC_mc_n78,
         top_core_EC_mc_n77, top_core_EC_mc_n76, top_core_EC_mc_n75,
         top_core_EC_mc_n74, top_core_EC_mc_n73, top_core_EC_mc_n72,
         top_core_EC_mc_n71, top_core_EC_mc_n70, top_core_EC_mc_n69,
         top_core_EC_mc_n68, top_core_EC_mc_n67, top_core_EC_mc_n66,
         top_core_EC_mc_n65, top_core_EC_mc_n64, top_core_EC_mc_n63,
         top_core_EC_mc_n62, top_core_EC_mc_n61, top_core_EC_mc_n60,
         top_core_EC_mc_n59, top_core_EC_mc_n58, top_core_EC_mc_n57,
         top_core_EC_mc_n56, top_core_EC_mc_n55, top_core_EC_mc_n54,
         top_core_EC_mc_n53, top_core_EC_mc_n52, top_core_EC_mc_n51,
         top_core_EC_mc_n50, top_core_EC_mc_n49, top_core_EC_mc_n48,
         top_core_EC_mc_n47, top_core_EC_mc_n46, top_core_EC_mc_n45,
         top_core_EC_mc_n44, top_core_EC_mc_n43, top_core_EC_mc_n42,
         top_core_EC_mc_n41, top_core_EC_mc_n40, top_core_EC_mc_n39,
         top_core_EC_mc_n38, top_core_EC_mc_n37, top_core_EC_mc_n36,
         top_core_EC_mc_n35, top_core_EC_mc_n34, top_core_EC_mc_n33,
         top_core_EC_mc_n32, top_core_EC_mc_n31, top_core_EC_mc_n30,
         top_core_EC_mc_n29, top_core_EC_mc_n28, top_core_EC_mc_n27,
         top_core_EC_mc_n26, top_core_EC_mc_n25, top_core_EC_mc_n24,
         top_core_EC_mc_n23, top_core_EC_mc_n22, top_core_EC_mc_n21,
         top_core_EC_mc_n20, top_core_EC_mc_n19, top_core_EC_mc_n18,
         top_core_EC_mc_n17, top_core_EC_mc_n16, top_core_EC_mc_n15,
         top_core_EC_mc_n14, top_core_EC_mc_n13, top_core_EC_mc_n12,
         top_core_EC_mc_n11, top_core_EC_mc_n10, top_core_EC_mc_n9,
         top_core_EC_mc_n8, top_core_EC_mc_n7, top_core_EC_mc_n6,
         top_core_EC_mc_n5, top_core_EC_mc_n4, top_core_EC_mc_n3,
         top_core_EC_mc_n2, top_core_EC_mc_mix_in_4_0_,
         top_core_EC_mc_mix_in_4_2_, top_core_EC_mc_mix_in_4_3_,
         top_core_EC_mc_mix_in_4_8_, top_core_EC_mc_mix_in_4_10_,
         top_core_EC_mc_mix_in_4_11_, top_core_EC_mc_mix_in_4_16_,
         top_core_EC_mc_mix_in_4_18_, top_core_EC_mc_mix_in_4_19_,
         top_core_EC_mc_mix_in_4_24_, top_core_EC_mc_mix_in_4_26_,
         top_core_EC_mc_mix_in_4_27_, top_core_EC_mc_mix_in_4_32_,
         top_core_EC_mc_mix_in_4_34_, top_core_EC_mc_mix_in_4_35_,
         top_core_EC_mc_mix_in_4_40_, top_core_EC_mc_mix_in_4_42_,
         top_core_EC_mc_mix_in_4_43_, top_core_EC_mc_mix_in_4_48_,
         top_core_EC_mc_mix_in_4_50_, top_core_EC_mc_mix_in_4_51_,
         top_core_EC_mc_mix_in_4_56_, top_core_EC_mc_mix_in_4_58_,
         top_core_EC_mc_mix_in_4_59_, top_core_EC_mc_mix_in_4_64_,
         top_core_EC_mc_mix_in_4_66_, top_core_EC_mc_mix_in_4_67_,
         top_core_EC_mc_mix_in_4_72_, top_core_EC_mc_mix_in_4_74_,
         top_core_EC_mc_mix_in_4_75_, top_core_EC_mc_mix_in_4_80_,
         top_core_EC_mc_mix_in_4_82_, top_core_EC_mc_mix_in_4_83_,
         top_core_EC_mc_mix_in_4_88_, top_core_EC_mc_mix_in_4_90_,
         top_core_EC_mc_mix_in_4_91_, top_core_EC_mc_mix_in_4_96_,
         top_core_EC_mc_mix_in_4_98_, top_core_EC_mc_mix_in_4_99_,
         top_core_EC_mc_mix_in_4_104_, top_core_EC_mc_mix_in_4_106_,
         top_core_EC_mc_mix_in_4_107_, top_core_EC_mc_mix_in_4_112_,
         top_core_EC_mc_mix_in_4_114_, top_core_EC_mc_mix_in_4_115_,
         top_core_EC_mc_mix_in_4_120_, top_core_EC_mc_mix_in_4_122_,
         top_core_EC_mc_mix_in_4_123_, top_core_EC_mc_mix_in_2_0_,
         top_core_EC_mc_mix_in_2_2_, top_core_EC_mc_mix_in_2_3_,
         top_core_EC_mc_mix_in_2_8_, top_core_EC_mc_mix_in_2_10_,
         top_core_EC_mc_mix_in_2_11_, top_core_EC_mc_mix_in_2_16_,
         top_core_EC_mc_mix_in_2_18_, top_core_EC_mc_mix_in_2_19_,
         top_core_EC_mc_mix_in_2_24_, top_core_EC_mc_mix_in_2_26_,
         top_core_EC_mc_mix_in_2_27_, top_core_EC_mc_mix_in_2_32_,
         top_core_EC_mc_mix_in_2_34_, top_core_EC_mc_mix_in_2_35_,
         top_core_EC_mc_mix_in_2_40_, top_core_EC_mc_mix_in_2_42_,
         top_core_EC_mc_mix_in_2_43_, top_core_EC_mc_mix_in_2_48_,
         top_core_EC_mc_mix_in_2_50_, top_core_EC_mc_mix_in_2_51_,
         top_core_EC_mc_mix_in_2_56_, top_core_EC_mc_mix_in_2_58_,
         top_core_EC_mc_mix_in_2_59_, top_core_EC_mc_mix_in_2_64_,
         top_core_EC_mc_mix_in_2_66_, top_core_EC_mc_mix_in_2_67_,
         top_core_EC_mc_mix_in_2_72_, top_core_EC_mc_mix_in_2_74_,
         top_core_EC_mc_mix_in_2_75_, top_core_EC_mc_mix_in_2_80_,
         top_core_EC_mc_mix_in_2_82_, top_core_EC_mc_mix_in_2_83_,
         top_core_EC_mc_mix_in_2_88_, top_core_EC_mc_mix_in_2_90_,
         top_core_EC_mc_mix_in_2_91_, top_core_EC_mc_mix_in_2_96_,
         top_core_EC_mc_mix_in_2_98_, top_core_EC_mc_mix_in_2_99_,
         top_core_EC_mc_mix_in_2_104_, top_core_EC_mc_mix_in_2_106_,
         top_core_EC_mc_mix_in_2_107_, top_core_EC_mc_mix_in_2_112_,
         top_core_EC_mc_mix_in_2_114_, top_core_EC_mc_mix_in_2_115_,
         top_core_EC_mc_mix_in_2_120_, top_core_EC_mc_mix_in_2_122_,
         top_core_EC_mc_mix_in_2_123_, top_core_KE_sb1_n374,
         top_core_KE_sb1_n373, top_core_KE_sb1_n372, top_core_KE_sb1_n371,
         top_core_KE_sb1_n370, top_core_KE_sb1_n368, top_core_KE_sb1_n367,
         top_core_KE_sb1_n366, top_core_KE_sb1_n365, top_core_KE_sb1_n364,
         top_core_KE_sb1_n363, top_core_KE_sb1_n362, top_core_KE_sb1_n361,
         top_core_KE_sb1_n360, top_core_KE_sb1_n359, top_core_KE_sb1_n358,
         top_core_KE_sb1_n357, top_core_KE_sb1_n356, top_core_KE_sb1_n355,
         top_core_KE_sb1_n354, top_core_KE_sb1_n353, top_core_KE_sb1_n352,
         top_core_KE_sb1_n351, top_core_KE_sb1_n350, top_core_KE_sb1_n349,
         top_core_KE_sb1_n348, top_core_KE_sb1_n347, top_core_KE_sb1_n346,
         top_core_KE_sb1_n345, top_core_KE_sb1_n344, top_core_KE_sb1_n343,
         top_core_KE_sb1_n342, top_core_KE_sb1_n341, top_core_KE_sb1_n340,
         top_core_KE_sb1_n339, top_core_KE_sb1_n338, top_core_KE_sb1_n337,
         top_core_KE_sb1_n336, top_core_KE_sb1_n335, top_core_KE_sb1_n334,
         top_core_KE_sb1_n333, top_core_KE_sb1_n332, top_core_KE_sb1_n331,
         top_core_KE_sb1_n330, top_core_KE_sb1_n329, top_core_KE_sb1_n328,
         top_core_KE_sb1_n327, top_core_KE_sb1_n326, top_core_KE_sb1_n325,
         top_core_KE_sb1_n324, top_core_KE_sb1_n323, top_core_KE_sb1_n322,
         top_core_KE_sb1_n321, top_core_KE_sb1_n320, top_core_KE_sb1_n319,
         top_core_KE_sb1_n318, top_core_KE_sb1_n317, top_core_KE_sb1_n316,
         top_core_KE_sb1_n315, top_core_KE_sb1_n314, top_core_KE_sb1_n313,
         top_core_KE_sb1_n312, top_core_KE_sb1_n311, top_core_KE_sb1_n310,
         top_core_KE_sb1_n309, top_core_KE_sb1_n308, top_core_KE_sb1_n307,
         top_core_KE_sb1_n306, top_core_KE_sb1_n305, top_core_KE_sb1_n304,
         top_core_KE_sb1_n303, top_core_KE_sb1_n302, top_core_KE_sb1_n301,
         top_core_KE_sb1_n300, top_core_KE_sb1_n299, top_core_KE_sb1_n298,
         top_core_KE_sb1_n297, top_core_KE_sb1_n296, top_core_KE_sb1_n295,
         top_core_KE_sb1_n294, top_core_KE_sb1_n293, top_core_KE_sb1_n292,
         top_core_KE_sb1_n291, top_core_KE_sb1_n290, top_core_KE_sb1_n289,
         top_core_KE_sb1_n288, top_core_KE_sb1_n287, top_core_KE_sb1_n286,
         top_core_KE_sb1_n285, top_core_KE_sb1_n284, top_core_KE_sb1_n283,
         top_core_KE_sb1_n282, top_core_KE_sb1_n281, top_core_KE_sb1_n280,
         top_core_KE_sb1_n279, top_core_KE_sb1_n278, top_core_KE_sb1_n277,
         top_core_KE_sb1_n276, top_core_KE_sb1_n275, top_core_KE_sb1_n274,
         top_core_KE_sb1_n273, top_core_KE_sb1_n272, top_core_KE_sb1_n271,
         top_core_KE_sb1_n270, top_core_KE_sb1_n269, top_core_KE_sb1_n268,
         top_core_KE_sb1_n267, top_core_KE_sb1_n266, top_core_KE_sb1_n265,
         top_core_KE_sb1_n264, top_core_KE_sb1_n263, top_core_KE_sb1_n262,
         top_core_KE_sb1_n261, top_core_KE_sb1_n260, top_core_KE_sb1_n259,
         top_core_KE_sb1_n258, top_core_KE_sb1_n257, top_core_KE_sb1_n256,
         top_core_KE_sb1_n255, top_core_KE_sb1_n254, top_core_KE_sb1_n253,
         top_core_KE_sb1_n252, top_core_KE_sb1_n251, top_core_KE_sb1_n250,
         top_core_KE_sb1_n249, top_core_KE_sb1_n247, top_core_KE_sb1_n246,
         top_core_KE_sb1_n245, top_core_KE_sb1_n244, top_core_KE_sb1_n243,
         top_core_KE_sb1_n242, top_core_KE_sb1_n241, top_core_KE_sb1_n240,
         top_core_KE_sb1_n239, top_core_KE_sb1_n238, top_core_KE_sb1_n237,
         top_core_KE_sb1_n236, top_core_KE_sb1_n235, top_core_KE_sb1_n234,
         top_core_KE_sb1_n233, top_core_KE_sb1_n232, top_core_KE_sb1_n231,
         top_core_KE_sb1_n230, top_core_KE_sb1_n229, top_core_KE_sb1_n228,
         top_core_KE_sb1_n227, top_core_KE_sb1_n226, top_core_KE_sb1_n225,
         top_core_KE_sb1_n224, top_core_KE_sb1_n223, top_core_KE_sb1_n222,
         top_core_KE_sb1_n221, top_core_KE_sb1_n220, top_core_KE_sb1_n219,
         top_core_KE_sb1_n218, top_core_KE_sb1_n217, top_core_KE_sb1_n216,
         top_core_KE_sb1_n215, top_core_KE_sb1_n214, top_core_KE_sb1_n213,
         top_core_KE_sb1_n212, top_core_KE_sb1_n211, top_core_KE_sb1_n210,
         top_core_KE_sb1_n209, top_core_KE_sb1_n208, top_core_KE_sb1_n207,
         top_core_KE_sb1_n206, top_core_KE_sb1_n205, top_core_KE_sb1_n204,
         top_core_KE_sb1_n203, top_core_KE_sb1_n202, top_core_KE_sb1_n201,
         top_core_KE_sb1_n200, top_core_KE_sb1_n199, top_core_KE_sb1_n198,
         top_core_KE_sb1_n197, top_core_KE_sb1_n196, top_core_KE_sb1_n195,
         top_core_KE_sb1_n194, top_core_KE_sb1_n193, top_core_KE_sb1_n192,
         top_core_KE_sb1_n191, top_core_KE_sb1_n190, top_core_KE_sb1_n189,
         top_core_KE_sb1_n188, top_core_KE_sb1_n187, top_core_KE_sb1_n186,
         top_core_KE_sb1_n185, top_core_KE_sb1_n184, top_core_KE_sb1_n183,
         top_core_KE_sb1_n182, top_core_KE_sb1_n181, top_core_KE_sb1_n180,
         top_core_KE_sb1_n179, top_core_KE_sb1_n178, top_core_KE_sb1_n177,
         top_core_KE_sb1_n176, top_core_KE_sb1_n175, top_core_KE_sb1_n174,
         top_core_KE_sb1_n173, top_core_KE_sb1_n171, top_core_KE_sb1_n170,
         top_core_KE_sb1_n169, top_core_KE_sb1_n168, top_core_KE_sb1_n167,
         top_core_KE_sb1_n166, top_core_KE_sb1_n165, top_core_KE_sb1_n164,
         top_core_KE_sb1_n163, top_core_KE_sb1_n162, top_core_KE_sb1_n161,
         top_core_KE_sb1_n160, top_core_KE_sb1_n159, top_core_KE_sb1_n158,
         top_core_KE_sb1_n157, top_core_KE_sb1_n156, top_core_KE_sb1_n155,
         top_core_KE_sb1_n154, top_core_KE_sb1_n153, top_core_KE_sb1_n152,
         top_core_KE_sb1_n151, top_core_KE_sb1_n150, top_core_KE_sb1_n149,
         top_core_KE_sb1_n148, top_core_KE_sb1_n147, top_core_KE_sb1_n146,
         top_core_KE_sb1_n145, top_core_KE_sb1_n144, top_core_KE_sb1_n143,
         top_core_KE_sb1_n141, top_core_KE_sb1_n140, top_core_KE_sb1_n139,
         top_core_KE_sb1_n138, top_core_KE_sb1_n137, top_core_KE_sb1_n136,
         top_core_KE_sb1_n134, top_core_KE_sb1_n133, top_core_KE_sb1_n132,
         top_core_KE_sb1_n131, top_core_KE_sb1_n130, top_core_KE_sb1_n129,
         top_core_KE_sb1_n128, top_core_KE_sb1_n127, top_core_KE_sb1_n126,
         top_core_KE_sb1_n125, top_core_KE_sb1_n124, top_core_KE_sb1_n123,
         top_core_KE_sb1_n122, top_core_KE_sb1_n121, top_core_KE_sb1_n120,
         top_core_KE_sb1_n119, top_core_KE_sb1_n118, top_core_KE_sb1_n117,
         top_core_KE_sb1_n116, top_core_KE_sb1_n115, top_core_KE_sb1_n114,
         top_core_KE_sb1_n113, top_core_KE_sb1_n112, top_core_KE_sb1_n111,
         top_core_KE_sb1_n110, top_core_KE_sb1_n109, top_core_KE_sb1_n108,
         top_core_KE_sb1_n107, top_core_KE_sb1_n106, top_core_KE_sb1_n105,
         top_core_KE_sb1_n104, top_core_KE_sb1_n103, top_core_KE_sb1_n102,
         top_core_KE_sb1_n101, top_core_KE_sb1_n100, top_core_KE_sb1_n99,
         top_core_KE_sb1_n98, top_core_KE_sb1_n97, top_core_KE_sb1_n96,
         top_core_KE_sb1_n95, top_core_KE_sb1_n94, top_core_KE_sb1_n93,
         top_core_KE_sb1_n92, top_core_KE_sb1_n91, top_core_KE_sb1_n90,
         top_core_KE_sb1_n89, top_core_KE_sb1_n88, top_core_KE_sb1_n87,
         top_core_KE_sb1_n86, top_core_KE_sb1_n85, top_core_KE_sb1_n84,
         top_core_KE_sb1_n83, top_core_KE_sb1_n82, top_core_KE_sb1_n81,
         top_core_KE_sb1_n80, top_core_KE_sb1_n79, top_core_KE_sb1_n78,
         top_core_KE_sb1_n77, top_core_KE_sb1_n76, top_core_KE_sb1_n75,
         top_core_KE_sb1_n74, top_core_KE_sb1_n73, top_core_KE_sb1_n72,
         top_core_KE_sb1_n71, top_core_KE_sb1_n70, top_core_KE_sb1_n69,
         top_core_KE_sb1_n68, top_core_KE_sb1_n67, top_core_KE_sb1_n66,
         top_core_KE_sb1_n65, top_core_KE_sb1_n64, top_core_KE_sb1_n63,
         top_core_KE_sb1_n62, top_core_KE_sb1_n61, top_core_KE_sb1_n60,
         top_core_KE_sb1_n59, top_core_KE_sb1_n58, top_core_KE_sb1_n57,
         top_core_KE_sb1_n56, top_core_KE_sb1_n55, top_core_KE_sb1_n54,
         top_core_KE_r343_u_div_PartRem_2__2_,
         top_core_KE_r343_u_div_PartRem_2__1_,
         top_core_KE_r343_u_div_PartRem_1__2_,
         top_core_KE_r343_u_div_PartRem_1__1_,
         top_core_KE_r343_u_div_SumTmp_2__1_,
         top_core_KE_r343_u_div_SumTmp_1__1_,
         top_core_KE_r343_u_div_SumTmp_0__1_, top_core_KE_r343_quotient_2_,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n354,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n353,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n352,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n351,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n350,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n349,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n348,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n347,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n346,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n345,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n344,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n343,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n342,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n341,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n340,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n339,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n338,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n337,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n336,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n335,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n334,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n333,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n332,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n331,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n330,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n329,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n328,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n327,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n326,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n325,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n324,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n323,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n322,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n321,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n320,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n319,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n318,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n317,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n316,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n315,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n314,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n313,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n312,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n311,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n310,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n309,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n308,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n307,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n306,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n305,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n304,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n303,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n302,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n301,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n300,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n299,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n298,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n297,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n296,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n295,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n294,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n293,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n292,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n291,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n290,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n289,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n288,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n287,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n286,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n285,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n284,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n283,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n282,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n281,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n280,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n279,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n278,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n277,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n276,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n275,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n274,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n273,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n272,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n271,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n270,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n269,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n268,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n267,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n266,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n265,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n264,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n263,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n262,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n261,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n260,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n259,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n258,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n257,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n256,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n255,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n254,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n253,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n252,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n251,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n250,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n249,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n248,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n247,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n246,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n245,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n244,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n243,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n242,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n241,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n240,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n239,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n238,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n237,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n236,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n235,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n234,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n233,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n232,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n231,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n230,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n229,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n228,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n227,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n226,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n225,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n224,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n223,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n222,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n221,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n220,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n219,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n218,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n217,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n216,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n215,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n214,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n213,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n212,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n211,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n210,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n209,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n208,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n207,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n206,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n205,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n204,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n203,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n202,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n201,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n200,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n199,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n198,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n197,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n196,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n195,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n194,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n193,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n192,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n191,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n190,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n189,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n188,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n187,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n186,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n185,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n184,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n183,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n182,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n181,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n180,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n179,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n178,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n177,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n176,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n175,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n174,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n173,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n172,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n171,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n170,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n169,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n168,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n167,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n166,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n165,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n164,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n163,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n162,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n161,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n160,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n159,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n158,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n157,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n156,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n155,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n154,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n152,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n151,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n150,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n149,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n148,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n147,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n146,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n145,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n144,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n143,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n142,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n141,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n140,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n139,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n138,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n137,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n136,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n135,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n134,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n133,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n132,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n131,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n130,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n129,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n128,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n127,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n126,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n125,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n124,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n123,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n122,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n121,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n120,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n119,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n118,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n117,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n116,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n115,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n114,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n113,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n112,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n111,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n110,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n109,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n108,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n107,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n106,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n105,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n104,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n102,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n101,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n100,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n99,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n98,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n97,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n96,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n95,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n94,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n93,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n92,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n91,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n89,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n88,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n87,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n86,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n85,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n84,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n83,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n82,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n81,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n80,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n79,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n78,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n77,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n76,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n75,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n74,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n73,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n71,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n70,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n69,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n68,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n67,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n66,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n65,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n64,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n63,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n62,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n61,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n60,
         top_core_EC_ss_gen_tbox_0__sboxs_r_n59, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732,
         n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, n743,
         n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754,
         n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
         n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776,
         n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, n787,
         n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798,
         n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809,
         n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
         n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831,
         n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
         n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853,
         n854, n855, n856, n857, n858, n859, n860, n861, n862, n863, n864,
         n865, n866, n867, n868, n869, n870, n871, n872, n873, n874, n875,
         n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
         n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
         n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
         n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
         n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
         n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
         n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
         n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
         n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
         n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
         n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
         n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
         n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
         n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
         n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
         n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
         n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
         n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
         n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
         n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
         n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
         n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
         n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
         n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18879;
  wire   [7:0] n_DIN;
  wire   [6:0] n_ADDR;
  wire   [7:0] n_DOUT;
  wire   [3:0] top_core_Addr;
  wire   [128:0] top_core_Key;
  wire   [2:0] top_core_Nk;
  wire   [255:0] top_core_CipherKey;
  wire   [3:1] top_core_Nr;
  wire   [127:0] top_core_Plain_text;
  wire   [127:0] top_core_Ciphertext;
  wire   [127:0] top_core_EC_ss_in;
  wire   [123:0] top_core_EC_mix_in;
  wire   [127:0] top_core_EC_add_in_r;
  wire   [127:0] top_core_EC_ss_sbox_out_r;
  wire   [127:0] top_core_EC_ss_sbox_out;
  wire   [127:0] top_core_EC_mc_mix_in_8;

  PIW PCLK ( .PAD(CLK), .C(n_CLK) );
  PIW PRSTB ( .PAD(RSTB), .C(n_RSTB) );
  PIW PSTART ( .PAD(START), .C(n_START) );
  PIW PWR ( .PAD(WR), .C(n_WR) );
  PO16W POK ( .I(n_OK), .PAD(OK) );
  CLKINVX8 top_core_KE_U4884 ( .A(n_RSTB), .Y(top_core_KE_n741) );
  JKFFRX4 top_core_KE_round_ctr_reg_reg_0_ ( .J(top_core_KE_n2705), .K(
        top_core_KE_n2719), .CK(n3906), .RN(n_RSTB), .Q(
        top_core_KE_round_ctr_reg_0_), .QN(top_core_KE_n728) );
  DFFX1 top_core_KE_prev_key0_reg_reg_71_ ( .D(top_core_KE_n4720), .CK(n3890), 
        .QN(top_core_KE_n651) );
  DFFX1 top_core_KE_prev_key0_reg_reg_79_ ( .D(top_core_KE_n4712), .CK(n3890), 
        .QN(top_core_KE_n643) );
  DFFX1 top_core_KE_prev_key0_reg_reg_87_ ( .D(top_core_KE_n4704), .CK(n3890), 
        .QN(top_core_KE_n635) );
  DFFX1 top_core_KE_prev_key0_reg_reg_70_ ( .D(top_core_KE_n4721), .CK(n3890), 
        .QN(top_core_KE_n652) );
  DFFX1 top_core_KE_prev_key0_reg_reg_78_ ( .D(top_core_KE_n4713), .CK(n3890), 
        .QN(top_core_KE_n644) );
  DFFX1 top_core_KE_prev_key0_reg_reg_86_ ( .D(top_core_KE_n4705), .CK(n3890), 
        .QN(top_core_KE_n636) );
  DFFX1 top_core_KE_prev_key0_reg_reg_84_ ( .D(top_core_KE_n4707), .CK(n3890), 
        .QN(top_core_KE_n638) );
  DFFX1 top_core_KE_prev_key0_reg_reg_82_ ( .D(top_core_KE_n4709), .CK(n3890), 
        .QN(top_core_KE_n640) );
  DFFX1 top_core_KE_prev_key0_reg_reg_81_ ( .D(top_core_KE_n4710), .CK(n3890), 
        .QN(top_core_KE_n641) );
  DFFX1 top_core_KE_prev_key0_reg_reg_68_ ( .D(top_core_KE_n4723), .CK(n3890), 
        .QN(top_core_KE_n654) );
  DFFX1 top_core_KE_prev_key0_reg_reg_76_ ( .D(top_core_KE_n4715), .CK(n3890), 
        .QN(top_core_KE_n646) );
  DFFX1 top_core_KE_prev_key0_reg_reg_66_ ( .D(top_core_KE_n4725), .CK(n3890), 
        .QN(top_core_KE_n656) );
  DFFX1 top_core_KE_prev_key0_reg_reg_65_ ( .D(top_core_KE_n4726), .CK(n3890), 
        .QN(top_core_KE_n657) );
  DFFX1 top_core_KE_prev_key0_reg_reg_73_ ( .D(top_core_KE_n4718), .CK(n3890), 
        .QN(top_core_KE_n649) );
  DFFX1 top_core_KE_prev_key0_reg_reg_64_ ( .D(top_core_KE_n4727), .CK(n3890), 
        .QN(top_core_KE_n658) );
  DFFX1 top_core_KE_prev_key0_reg_reg_85_ ( .D(top_core_KE_n4706), .CK(n3889), 
        .QN(top_core_KE_n637) );
  DFFX1 top_core_KE_prev_key0_reg_reg_83_ ( .D(top_core_KE_n4708), .CK(n3889), 
        .QN(top_core_KE_n639) );
  DFFX1 top_core_KE_prev_key0_reg_reg_80_ ( .D(top_core_KE_n4711), .CK(n3889), 
        .QN(top_core_KE_n642) );
  DFFX1 top_core_KE_prev_key0_reg_reg_69_ ( .D(top_core_KE_n4722), .CK(n3889), 
        .QN(top_core_KE_n653) );
  DFFX1 top_core_KE_prev_key0_reg_reg_77_ ( .D(top_core_KE_n4714), .CK(n3889), 
        .QN(top_core_KE_n645) );
  DFFX1 top_core_KE_prev_key0_reg_reg_67_ ( .D(top_core_KE_n4724), .CK(n3889), 
        .QN(top_core_KE_n655) );
  DFFX1 top_core_KE_prev_key0_reg_reg_75_ ( .D(top_core_KE_n4716), .CK(n3889), 
        .QN(top_core_KE_n647) );
  DFFX1 top_core_KE_prev_key0_reg_reg_74_ ( .D(top_core_KE_n4717), .CK(n3889), 
        .QN(top_core_KE_n648) );
  DFFX1 top_core_KE_prev_key0_reg_reg_72_ ( .D(top_core_KE_n4719), .CK(n3889), 
        .QN(top_core_KE_n650) );
  DFFHQX1 top_core_KE_Nk0_reg_0_ ( .D(top_core_Nk[0]), .CK(n3695), .Q(
        top_core_KE_Nk0_0_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_31_ ( .D(top_core_KE_n4888), .CK(n3902), .Q(top_core_KE_prev_key1_reg_31_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_94_ ( .D(top_core_KE_n4825), .CK(n3896), .Q(top_core_KE_prev_key1_reg_94_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_30_ ( .D(top_core_KE_n4889), .CK(n3897), .Q(top_core_KE_prev_key1_reg_30_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_84_ ( .D(top_core_KE_n4835), .CK(n3891), .Q(top_core_KE_prev_key1_reg_84_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_20_ ( .D(top_core_KE_n4899), .CK(n3891), .Q(top_core_KE_prev_key1_reg_20_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_92_ ( .D(top_core_KE_n4827), .CK(n3891), .Q(top_core_KE_prev_key1_reg_92_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_28_ ( .D(top_core_KE_n4891), .CK(n3892), .Q(top_core_KE_prev_key1_reg_28_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_83_ ( .D(top_core_KE_n4836), .CK(n3905), .Q(top_core_KE_prev_key1_reg_83_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_19_ ( .D(top_core_KE_n4900), .CK(n3904), .Q(top_core_KE_prev_key1_reg_19_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_91_ ( .D(top_core_KE_n4828), .CK(n3904), .Q(top_core_KE_prev_key1_reg_91_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_27_ ( .D(top_core_KE_n4892), .CK(n3903), .Q(top_core_KE_prev_key1_reg_27_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_18_ ( .D(top_core_KE_n4901), .CK(n3901), .Q(top_core_KE_prev_key1_reg_18_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_26_ ( .D(top_core_KE_n4893), .CK(n3899), .Q(top_core_KE_prev_key1_reg_26_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_22_ ( .D(top_core_KE_n4897), .CK(n3899), .Q(top_core_KE_prev_key1_reg_22_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_86_ ( .D(top_core_KE_n4833), .CK(n3899), .Q(top_core_KE_prev_key1_reg_86_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_78_ ( .D(top_core_KE_n4841), .CK(n3899), .Q(top_core_KE_prev_key1_reg_78_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_14_ ( .D(top_core_KE_n4905), .CK(n3899), .Q(top_core_KE_prev_key1_reg_14_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_68_ ( .D(top_core_KE_n4851), .CK(n3901), .Q(top_core_KE_prev_key1_reg_68_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_4_ ( .D(top_core_KE_n4915), .CK(n3902), 
        .Q(top_core_KE_prev_key1_reg_4_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_76_ ( .D(top_core_KE_n4843), .CK(n3903), .Q(top_core_KE_prev_key1_reg_76_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_12_ ( .D(top_core_KE_n4907), .CK(n3903), .Q(top_core_KE_prev_key1_reg_12_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_67_ ( .D(top_core_KE_n4852), .CK(n3904), .Q(top_core_KE_prev_key1_reg_67_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_3_ ( .D(top_core_KE_n4916), .CK(n3904), 
        .Q(top_core_KE_prev_key1_reg_3_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_75_ ( .D(top_core_KE_n4844), .CK(n3905), .Q(top_core_KE_prev_key1_reg_75_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_11_ ( .D(top_core_KE_n4908), .CK(n3905), .Q(top_core_KE_prev_key1_reg_11_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_2_ ( .D(top_core_KE_n4917), .CK(n3906), 
        .Q(top_core_KE_prev_key1_reg_2_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_10_ ( .D(top_core_KE_n4909), .CK(n3891), .Q(top_core_KE_prev_key1_reg_10_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_6_ ( .D(top_core_KE_n4913), .CK(n3895), 
        .Q(top_core_KE_prev_key1_reg_6_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_70_ ( .D(top_core_KE_n4849), .CK(n3895), .Q(top_core_KE_prev_key1_reg_70_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_95_ ( .D(top_core_KE_n4824), .CK(n3895), .Q(top_core_KE_prev_key1_reg_95_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_87_ ( .D(top_core_KE_n4832), .CK(n3895), .Q(top_core_KE_prev_key1_reg_87_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_23_ ( .D(top_core_KE_n4896), .CK(n3895), .Q(top_core_KE_prev_key1_reg_23_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_15_ ( .D(top_core_KE_n4904), .CK(n3895), .Q(top_core_KE_prev_key1_reg_15_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_79_ ( .D(top_core_KE_n4840), .CK(n3895), .Q(top_core_KE_prev_key1_reg_79_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_71_ ( .D(top_core_KE_n4848), .CK(n3895), .Q(top_core_KE_prev_key1_reg_71_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_7_ ( .D(top_core_KE_n4912), .CK(n3896), 
        .Q(top_core_KE_prev_key1_reg_7_) );
  DFFRHQX1 top_core_EC_Addr_reg_1_ ( .D(top_core_EC_n1293), .CK(n3721), .RN(
        n_RSTB), .Q(top_core_Addr[1]) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_81_ ( .D(top_core_KE_n4838), .CK(n3892), .Q(top_core_KE_prev_key1_reg_81_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_17_ ( .D(top_core_KE_n4902), .CK(n3897), .Q(top_core_KE_prev_key1_reg_17_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_80_ ( .D(top_core_KE_n4839), .CK(n3898), .Q(top_core_KE_prev_key1_reg_80_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_16_ ( .D(top_core_KE_n4903), .CK(n3898), .Q(top_core_KE_prev_key1_reg_16_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_88_ ( .D(top_core_KE_n4831), .CK(n3898), .Q(top_core_KE_prev_key1_reg_88_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_24_ ( .D(top_core_KE_n4895), .CK(n3898), .Q(top_core_KE_prev_key1_reg_24_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_65_ ( .D(top_core_KE_n4854), .CK(n3891), .Q(top_core_KE_prev_key1_reg_65_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_1_ ( .D(top_core_KE_n4918), .CK(n3892), 
        .Q(top_core_KE_prev_key1_reg_1_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_73_ ( .D(top_core_KE_n4846), .CK(n3897), .Q(top_core_KE_prev_key1_reg_73_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_9_ ( .D(top_core_KE_n4910), .CK(n3893), 
        .Q(top_core_KE_prev_key1_reg_9_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_64_ ( .D(top_core_KE_n4855), .CK(n3893), .Q(top_core_KE_prev_key1_reg_64_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_0_ ( .D(top_core_KE_n4919), .CK(n3894), 
        .Q(top_core_KE_prev_key1_reg_0_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_72_ ( .D(top_core_KE_n4847), .CK(n3895), .Q(top_core_KE_prev_key1_reg_72_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_8_ ( .D(top_core_KE_n4911), .CK(n3895), 
        .Q(top_core_KE_prev_key1_reg_8_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_25_ ( .D(top_core_KE_n4894), .CK(n3896), .Q(top_core_KE_prev_key1_reg_25_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_82_ ( .D(top_core_KE_n4837), .CK(n3901), .Q(top_core_KE_prev_key1_reg_82_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_66_ ( .D(top_core_KE_n4853), .CK(n3906), .Q(top_core_KE_prev_key1_reg_66_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_74_ ( .D(top_core_KE_n4845), .CK(n3891), .Q(top_core_KE_prev_key1_reg_74_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_89_ ( .D(top_core_KE_n4830), .CK(n3896), .Q(top_core_KE_prev_key1_reg_89_) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_127_ ( .D(top_core_EC_N276), .CK(n3795), .RN(n_RSTB), .Q(top_core_Ciphertext[7]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_126_ ( .D(top_core_EC_N275), .CK(n3795), .RN(n_RSTB), .Q(top_core_Ciphertext[6]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_125_ ( .D(top_core_EC_N274), .CK(n3795), .RN(n_RSTB), .Q(top_core_Ciphertext[5]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_124_ ( .D(top_core_EC_N273), .CK(n3795), .RN(n_RSTB), .Q(top_core_Ciphertext[4]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_123_ ( .D(top_core_EC_N272), .CK(n3795), .RN(n_RSTB), .Q(top_core_Ciphertext[3]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_122_ ( .D(top_core_EC_N271), .CK(n3795), .RN(n_RSTB), .Q(top_core_Ciphertext[2]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_121_ ( .D(top_core_EC_N270), .CK(n3795), .RN(n_RSTB), .Q(top_core_Ciphertext[1]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_120_ ( .D(top_core_EC_N269), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[0]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_119_ ( .D(top_core_EC_N268), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[15]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_118_ ( .D(top_core_EC_N267), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[14]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_117_ ( .D(top_core_EC_N266), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[13]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_116_ ( .D(top_core_EC_N265), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[12]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_115_ ( .D(top_core_EC_N264), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[11]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_114_ ( .D(top_core_EC_N263), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[10]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_113_ ( .D(top_core_EC_N262), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[9]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_112_ ( .D(top_core_EC_N261), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[8]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_111_ ( .D(top_core_EC_N260), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[23]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_110_ ( .D(top_core_EC_N259), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[22]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_109_ ( .D(top_core_EC_N258), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[21]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_108_ ( .D(top_core_EC_N257), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[20]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_107_ ( .D(top_core_EC_N256), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[19]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_106_ ( .D(top_core_EC_N255), .CK(n3796), .RN(n_RSTB), .Q(top_core_Ciphertext[18]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_105_ ( .D(top_core_EC_N254), .CK(n3797), .RN(n_RSTB), .Q(top_core_Ciphertext[17]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_104_ ( .D(top_core_EC_N253), .CK(n3797), .RN(n_RSTB), .Q(top_core_Ciphertext[16]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_103_ ( .D(top_core_EC_N252), .CK(n3797), .RN(n_RSTB), .Q(top_core_Ciphertext[31]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_102_ ( .D(top_core_EC_N251), .CK(n3797), .RN(n_RSTB), .Q(top_core_Ciphertext[30]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_101_ ( .D(top_core_EC_N250), .CK(n3797), .RN(n_RSTB), .Q(top_core_Ciphertext[29]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_100_ ( .D(top_core_EC_N249), .CK(n3797), .RN(n_RSTB), .Q(top_core_Ciphertext[28]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_99_ ( .D(top_core_EC_N248), .CK(n3797), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[27]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_98_ ( .D(top_core_EC_N247), .CK(n3797), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[26]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_97_ ( .D(top_core_EC_N246), .CK(n3797), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[25]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_96_ ( .D(top_core_EC_N245), .CK(n3797), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[24]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_95_ ( .D(top_core_EC_N244), .CK(n3797), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[39]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_94_ ( .D(top_core_EC_N243), .CK(n3797), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[38]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_93_ ( .D(top_core_EC_N242), .CK(n3797), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[37]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_92_ ( .D(top_core_EC_N241), .CK(n3797), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[36]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_91_ ( .D(top_core_EC_N240), .CK(n3797), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[35]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_90_ ( .D(top_core_EC_N239), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[34]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_89_ ( .D(top_core_EC_N238), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[33]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_88_ ( .D(top_core_EC_N237), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[32]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_87_ ( .D(top_core_EC_N236), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[47]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_86_ ( .D(top_core_EC_N235), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[46]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_85_ ( .D(top_core_EC_N234), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[45]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_84_ ( .D(top_core_EC_N233), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[44]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_83_ ( .D(top_core_EC_N232), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[43]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_82_ ( .D(top_core_EC_N231), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[42]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_81_ ( .D(top_core_EC_N230), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[41]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_80_ ( .D(top_core_EC_N229), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[40]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_79_ ( .D(top_core_EC_N228), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[55]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_78_ ( .D(top_core_EC_N227), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[54]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_77_ ( .D(top_core_EC_N226), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[53]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_76_ ( .D(top_core_EC_N225), .CK(n3798), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[52]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_75_ ( .D(top_core_EC_N224), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[51]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_74_ ( .D(top_core_EC_N223), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[50]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_73_ ( .D(top_core_EC_N222), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[49]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_72_ ( .D(top_core_EC_N221), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[48]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_71_ ( .D(top_core_EC_N220), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[63]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_70_ ( .D(top_core_EC_N219), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[62]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_69_ ( .D(top_core_EC_N218), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[61]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_68_ ( .D(top_core_EC_N217), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[60]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_67_ ( .D(top_core_EC_N216), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[59]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_66_ ( .D(top_core_EC_N215), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[58]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_65_ ( .D(top_core_EC_N214), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[57]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_64_ ( .D(top_core_EC_N213), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[56]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_63_ ( .D(top_core_EC_N212), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[71]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_62_ ( .D(top_core_EC_N211), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[70]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_61_ ( .D(top_core_EC_N210), .CK(n3799), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[69]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_60_ ( .D(top_core_EC_N209), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[68]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_59_ ( .D(top_core_EC_N208), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[67]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_58_ ( .D(top_core_EC_N207), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[66]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_57_ ( .D(top_core_EC_N206), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[65]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_56_ ( .D(top_core_EC_N205), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[64]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_55_ ( .D(top_core_EC_N204), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[79]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_54_ ( .D(top_core_EC_N203), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[78]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_53_ ( .D(top_core_EC_N202), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[77]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_52_ ( .D(top_core_EC_N201), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[76]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_51_ ( .D(top_core_EC_N200), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[75]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_50_ ( .D(top_core_EC_N199), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[74]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_49_ ( .D(top_core_EC_N198), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[73]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_48_ ( .D(top_core_EC_N197), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[72]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_47_ ( .D(top_core_EC_N196), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[87]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_46_ ( .D(top_core_EC_N195), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[86]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_45_ ( .D(top_core_EC_N194), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[85]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_44_ ( .D(top_core_EC_N193), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[84]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_43_ ( .D(top_core_EC_N192), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[83]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_42_ ( .D(top_core_EC_N191), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[82]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_41_ ( .D(top_core_EC_N190), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[81]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_40_ ( .D(top_core_EC_N189), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[80]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_39_ ( .D(top_core_EC_N188), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[95]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_38_ ( .D(top_core_EC_N187), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[94]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_37_ ( .D(top_core_EC_N186), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[93]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_36_ ( .D(top_core_EC_N185), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[92]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_35_ ( .D(top_core_EC_N184), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[91]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_34_ ( .D(top_core_EC_N183), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[90]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_33_ ( .D(top_core_EC_N182), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[89]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_32_ ( .D(top_core_EC_N181), .CK(n3801), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[88]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_31_ ( .D(top_core_EC_N180), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[103]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_30_ ( .D(top_core_EC_N179), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[102]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_29_ ( .D(top_core_EC_N178), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[101]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_28_ ( .D(top_core_EC_N177), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[100]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_27_ ( .D(top_core_EC_N176), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[99]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_26_ ( .D(top_core_EC_N175), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[98]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_25_ ( .D(top_core_EC_N174), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[97]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_24_ ( .D(top_core_EC_N173), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[96]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_23_ ( .D(top_core_EC_N172), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[111]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_22_ ( .D(top_core_EC_N171), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[110]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_21_ ( .D(top_core_EC_N170), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[109]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_20_ ( .D(top_core_EC_N169), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[108]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_19_ ( .D(top_core_EC_N168), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[107]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_18_ ( .D(top_core_EC_N167), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[106]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_17_ ( .D(top_core_EC_N166), .CK(n3802), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[105]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_16_ ( .D(top_core_EC_N165), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[104]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_15_ ( .D(top_core_EC_N164), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[119]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_14_ ( .D(top_core_EC_N163), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[118]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_13_ ( .D(top_core_EC_N162), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[117]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_12_ ( .D(top_core_EC_N161), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[116]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_11_ ( .D(top_core_EC_N160), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[115]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_10_ ( .D(top_core_EC_N159), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[114]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_9_ ( .D(top_core_EC_N158), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[113]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_8_ ( .D(top_core_EC_N157), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[112]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_7_ ( .D(top_core_EC_N156), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[127]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_6_ ( .D(top_core_EC_N155), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[126]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_5_ ( .D(top_core_EC_N154), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[125]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_4_ ( .D(top_core_EC_N153), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[124]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_3_ ( .D(top_core_EC_N152), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[123]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_2_ ( .D(top_core_EC_N151), .CK(n3803), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[122]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_1_ ( .D(top_core_EC_N150), .CK(n3804), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[121]) );
  DFFRHQX1 top_core_EC_Ciphertext_r_reg_0_ ( .D(top_core_EC_N149), .CK(n3804), 
        .RN(n_RSTB), .Q(top_core_Ciphertext[120]) );
  DFFHQX1 top_core_KE_CipherKey0_reg_192_ ( .D(top_core_CipherKey[192]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_192_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_193_ ( .D(top_core_CipherKey[193]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_193_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_194_ ( .D(top_core_CipherKey[194]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_194_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_195_ ( .D(top_core_CipherKey[195]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_195_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_196_ ( .D(top_core_CipherKey[196]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_196_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_197_ ( .D(top_core_CipherKey[197]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_197_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_198_ ( .D(top_core_CipherKey[198]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_198_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_199_ ( .D(top_core_CipherKey[199]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_199_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_200_ ( .D(top_core_CipherKey[200]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_200_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_201_ ( .D(top_core_CipherKey[201]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_201_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_202_ ( .D(top_core_CipherKey[202]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_202_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_203_ ( .D(top_core_CipherKey[203]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_203_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_204_ ( .D(top_core_CipherKey[204]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_204_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_205_ ( .D(top_core_CipherKey[205]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_205_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_206_ ( .D(top_core_CipherKey[206]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_206_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_207_ ( .D(top_core_CipherKey[207]), .CK(
        n3699), .Q(top_core_KE_CipherKey0_207_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_208_ ( .D(top_core_CipherKey[208]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_208_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_209_ ( .D(top_core_CipherKey[209]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_209_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_210_ ( .D(top_core_CipherKey[210]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_210_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_211_ ( .D(top_core_CipherKey[211]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_211_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_212_ ( .D(top_core_CipherKey[212]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_212_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_213_ ( .D(top_core_CipherKey[213]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_213_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_214_ ( .D(top_core_CipherKey[214]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_214_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_215_ ( .D(top_core_CipherKey[215]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_215_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_216_ ( .D(top_core_CipherKey[216]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_216_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_217_ ( .D(top_core_CipherKey[217]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_217_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_218_ ( .D(top_core_CipherKey[218]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_218_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_219_ ( .D(top_core_CipherKey[219]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_219_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_220_ ( .D(top_core_CipherKey[220]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_220_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_221_ ( .D(top_core_CipherKey[221]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_221_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_222_ ( .D(top_core_CipherKey[222]), .CK(
        n3698), .Q(top_core_KE_CipherKey0_222_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_223_ ( .D(top_core_CipherKey[223]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_223_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_224_ ( .D(top_core_CipherKey[224]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_224_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_225_ ( .D(top_core_CipherKey[225]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_225_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_226_ ( .D(top_core_CipherKey[226]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_226_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_227_ ( .D(top_core_CipherKey[227]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_227_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_228_ ( .D(top_core_CipherKey[228]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_228_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_229_ ( .D(top_core_CipherKey[229]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_229_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_230_ ( .D(top_core_CipherKey[230]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_230_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_231_ ( .D(top_core_CipherKey[231]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_231_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_232_ ( .D(top_core_CipherKey[232]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_232_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_233_ ( .D(top_core_CipherKey[233]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_233_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_234_ ( .D(top_core_CipherKey[234]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_234_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_235_ ( .D(top_core_CipherKey[235]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_235_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_236_ ( .D(top_core_CipherKey[236]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_236_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_237_ ( .D(top_core_CipherKey[237]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_237_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_238_ ( .D(top_core_CipherKey[238]), .CK(
        n3697), .Q(top_core_KE_CipherKey0_238_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_239_ ( .D(top_core_CipherKey[239]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_239_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_240_ ( .D(top_core_CipherKey[240]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_240_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_241_ ( .D(top_core_CipherKey[241]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_241_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_242_ ( .D(top_core_CipherKey[242]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_242_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_243_ ( .D(top_core_CipherKey[243]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_243_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_244_ ( .D(top_core_CipherKey[244]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_244_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_245_ ( .D(top_core_CipherKey[245]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_245_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_246_ ( .D(top_core_CipherKey[246]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_246_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_247_ ( .D(top_core_CipherKey[247]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_247_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_248_ ( .D(top_core_CipherKey[248]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_248_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_249_ ( .D(top_core_CipherKey[249]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_249_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_250_ ( .D(top_core_CipherKey[250]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_250_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_251_ ( .D(top_core_CipherKey[251]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_251_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_252_ ( .D(top_core_CipherKey[252]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_252_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_253_ ( .D(top_core_CipherKey[253]), .CK(
        n3696), .Q(top_core_KE_CipherKey0_253_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_254_ ( .D(top_core_CipherKey[254]), .CK(
        n3695), .Q(top_core_KE_CipherKey0_254_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_255_ ( .D(top_core_CipherKey[255]), .CK(
        n3695), .Q(top_core_KE_CipherKey0_255_) );
  DFFRHQX1 top_core_io_Nr_reg_1_ ( .D(top_core_io_N125), .CK(n3806), .RN(
        n_RSTB), .Q(top_core_Nr[1]) );
  DFFRHQX1 top_core_io_Nr_reg_2_ ( .D(top_core_io_N126), .CK(n3775), .RN(
        n_RSTB), .Q(top_core_Nr[2]) );
  DFFRHQX1 top_core_io_Nr_reg_3_ ( .D(top_core_io_N127), .CK(n3769), .RN(
        n_RSTB), .Q(top_core_Nr[3]) );
  DFFRHQX1 top_core_io_op_reg ( .D(top_core_io_N515), .CK(n3795), .RN(n_RSTB), 
        .Q(top_core_op) );
  DFFRHQX1 top_core_EC_round_result_r_reg_57_ ( .D(top_core_EC_n1233), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_57_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_56_ ( .D(top_core_EC_n1234), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_56_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_55_ ( .D(top_core_EC_n1235), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_55_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_54_ ( .D(top_core_EC_n1236), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_54_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_53_ ( .D(top_core_EC_n1237), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_53_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_52_ ( .D(top_core_EC_n1238), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_52_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_51_ ( .D(top_core_EC_n1239), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_51_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_50_ ( .D(top_core_EC_n1240), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_50_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_49_ ( .D(top_core_EC_n1241), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_49_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_48_ ( .D(top_core_EC_n1242), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_48_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_47_ ( .D(top_core_EC_n1243), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_47_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_46_ ( .D(top_core_EC_n1244), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_46_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_45_ ( .D(top_core_EC_n1245), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_45_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_44_ ( .D(top_core_EC_n1246), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_44_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_43_ ( .D(top_core_EC_n1247), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_43_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_42_ ( .D(top_core_EC_n1248), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_42_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_41_ ( .D(top_core_EC_n1249), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_41_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_40_ ( .D(top_core_EC_n1250), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_40_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_39_ ( .D(top_core_EC_n1251), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_39_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_38_ ( .D(top_core_EC_n1252), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_38_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_37_ ( .D(top_core_EC_n1253), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_37_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_36_ ( .D(top_core_EC_n1254), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_36_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_35_ ( .D(top_core_EC_n1255), .CK(
        n3793), .RN(n_RSTB), .Q(top_core_EC_round_result_r_35_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_34_ ( .D(top_core_EC_n1256), .CK(
        n3794), .RN(n_RSTB), .Q(top_core_EC_round_result_r_34_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_33_ ( .D(top_core_EC_n1257), .CK(
        n3794), .RN(n_RSTB), .Q(top_core_EC_round_result_r_33_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_32_ ( .D(top_core_EC_n1258), .CK(
        n3794), .RN(n_RSTB), .Q(top_core_EC_round_result_r_32_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_31_ ( .D(top_core_EC_n1259), .CK(
        n3794), .RN(n_RSTB), .Q(top_core_EC_round_result_r_31_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_30_ ( .D(top_core_EC_n1260), .CK(
        n3794), .RN(n_RSTB), .Q(top_core_EC_round_result_r_30_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_29_ ( .D(top_core_EC_n1261), .CK(
        n3794), .RN(n_RSTB), .Q(top_core_EC_round_result_r_29_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_28_ ( .D(top_core_EC_n1262), .CK(
        n3732), .RN(n_RSTB), .Q(top_core_EC_round_result_r_28_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_27_ ( .D(top_core_EC_n1263), .CK(
        n3725), .RN(n_RSTB), .Q(top_core_EC_round_result_r_27_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_26_ ( .D(top_core_EC_n1264), .CK(
        n3719), .RN(n_RSTB), .Q(top_core_EC_round_result_r_26_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_25_ ( .D(top_core_EC_n1265), .CK(
        n3719), .RN(n_RSTB), .Q(top_core_EC_round_result_r_25_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_24_ ( .D(top_core_EC_n1266), .CK(
        n3719), .RN(n_RSTB), .Q(top_core_EC_round_result_r_24_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_23_ ( .D(top_core_EC_n1267), .CK(
        n3719), .RN(n_RSTB), .Q(top_core_EC_round_result_r_23_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_22_ ( .D(top_core_EC_n1268), .CK(
        n3719), .RN(n_RSTB), .Q(top_core_EC_round_result_r_22_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_21_ ( .D(top_core_EC_n1269), .CK(
        n3719), .RN(n_RSTB), .Q(top_core_EC_round_result_r_21_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_20_ ( .D(top_core_EC_n1270), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_20_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_19_ ( .D(top_core_EC_n1271), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_19_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_18_ ( .D(top_core_EC_n1272), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_18_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_17_ ( .D(top_core_EC_n1273), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_17_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_16_ ( .D(top_core_EC_n1274), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_16_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_15_ ( .D(top_core_EC_n1275), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_15_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_14_ ( .D(top_core_EC_n1276), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_14_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_13_ ( .D(top_core_EC_n1277), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_13_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_12_ ( .D(top_core_EC_n1278), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_12_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_11_ ( .D(top_core_EC_n1279), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_11_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_10_ ( .D(top_core_EC_n1280), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_10_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_9_ ( .D(top_core_EC_n1281), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_9_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_8_ ( .D(top_core_EC_n1282), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_8_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_7_ ( .D(top_core_EC_n1283), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_7_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_6_ ( .D(top_core_EC_n1284), .CK(
        n3720), .RN(n_RSTB), .Q(top_core_EC_round_result_r_6_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_5_ ( .D(top_core_EC_n1285), .CK(
        n3721), .RN(n_RSTB), .Q(top_core_EC_round_result_r_5_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_4_ ( .D(top_core_EC_n1286), .CK(
        n3721), .RN(n_RSTB), .Q(top_core_EC_round_result_r_4_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_3_ ( .D(top_core_EC_n1287), .CK(
        n3721), .RN(n_RSTB), .Q(top_core_EC_round_result_r_3_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_2_ ( .D(top_core_EC_n1288), .CK(
        n3721), .RN(n_RSTB), .Q(top_core_EC_round_result_r_2_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_1_ ( .D(top_core_EC_n1289), .CK(
        n3721), .RN(n_RSTB), .Q(top_core_EC_round_result_r_1_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_0_ ( .D(top_core_EC_n1290), .CK(
        n3721), .RN(n_RSTB), .Q(top_core_EC_round_result_r_0_) );
  DFFRHQX1 top_core_EC_Addr_reg_3_ ( .D(top_core_EC_n1291), .CK(n3721), .RN(
        n_RSTB), .Q(top_core_Addr[3]) );
  DFFRHQX1 top_core_EC_Addr_reg_2_ ( .D(top_core_EC_n1292), .CK(n3721), .RN(
        n_RSTB), .Q(top_core_Addr[2]) );
  DFFRHQX1 top_core_KE_round_ctr_reg_reg_3_ ( .D(top_core_KE_n4929), .CK(n3837), .RN(n_RSTB), .Q(top_core_KE_round_ctr_reg_3_) );
  DFFRHQX1 top_core_KE_round_ctr_reg_reg_2_ ( .D(top_core_KE_n4930), .CK(n3837), .RN(n_RSTB), .Q(top_core_KE_round_ctr_reg_2_) );
  DFFRHQX1 top_core_KE_round_ctr_reg_reg_1_ ( .D(top_core_KE_n4931), .CK(n3837), .RN(n_RSTB), .Q(top_core_KE_round_ctr_reg_1_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_63_ ( .D(top_core_KE_n4728), .CK(n3902), .Q(top_core_KE_prev_key0_reg_63_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_119_ ( .D(top_core_KE_n4673), .CK(
        n3891), .Q(top_core_KE_prev_key0_reg_119_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_118_ ( .D(top_core_KE_n4674), .CK(
        n3896), .Q(top_core_KE_prev_key0_reg_118_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_117_ ( .D(top_core_KE_n4675), .CK(
        n3894), .Q(top_core_KE_prev_key0_reg_117_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_116_ ( .D(top_core_KE_n4676), .CK(
        n3892), .Q(top_core_KE_prev_key0_reg_116_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_115_ ( .D(top_core_KE_n4677), .CK(
        n3904), .Q(top_core_KE_prev_key0_reg_115_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_114_ ( .D(top_core_KE_n4678), .CK(
        n3901), .Q(top_core_KE_prev_key0_reg_114_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_113_ ( .D(top_core_KE_n4679), .CK(
        n3901), .Q(top_core_KE_prev_key0_reg_113_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_112_ ( .D(top_core_KE_n4680), .CK(
        n3898), .Q(top_core_KE_prev_key0_reg_112_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_63_ ( .D(top_core_CipherKey[63]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_63_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_85_ ( .D(top_core_KE_n4834), .CK(n3895), .Q(top_core_KE_prev_key1_reg_85_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_69_ ( .D(top_core_KE_n4850), .CK(n3900), .Q(top_core_KE_prev_key1_reg_69_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_77_ ( .D(top_core_KE_n4842), .CK(n3901), .Q(top_core_KE_prev_key1_reg_77_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_0_ ( .D(top_core_CipherKey[0]), .CK(n3695), .Q(top_core_KE_CipherKey0_0_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_1_ ( .D(top_core_CipherKey[1]), .CK(n3695), .Q(top_core_KE_CipherKey0_1_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_2_ ( .D(top_core_CipherKey[2]), .CK(n3695), .Q(top_core_KE_CipherKey0_2_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_3_ ( .D(top_core_CipherKey[3]), .CK(n3695), .Q(top_core_KE_CipherKey0_3_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_4_ ( .D(top_core_CipherKey[4]), .CK(n3695), .Q(top_core_KE_CipherKey0_4_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_5_ ( .D(top_core_CipherKey[5]), .CK(n3695), .Q(top_core_KE_CipherKey0_5_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_6_ ( .D(top_core_CipherKey[6]), .CK(n3695), .Q(top_core_KE_CipherKey0_6_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_7_ ( .D(top_core_CipherKey[7]), .CK(n3695), .Q(top_core_KE_CipherKey0_7_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_8_ ( .D(top_core_CipherKey[8]), .CK(n3695), .Q(top_core_KE_CipherKey0_8_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_9_ ( .D(top_core_CipherKey[9]), .CK(n3695), .Q(top_core_KE_CipherKey0_9_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_10_ ( .D(top_core_CipherKey[10]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_10_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_11_ ( .D(top_core_CipherKey[11]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_11_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_12_ ( .D(top_core_CipherKey[12]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_12_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_13_ ( .D(top_core_CipherKey[13]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_13_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_14_ ( .D(top_core_CipherKey[14]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_14_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_15_ ( .D(top_core_CipherKey[15]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_15_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_16_ ( .D(top_core_CipherKey[16]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_16_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_17_ ( .D(top_core_CipherKey[17]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_17_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_18_ ( .D(top_core_CipherKey[18]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_18_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_19_ ( .D(top_core_CipherKey[19]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_19_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_20_ ( .D(top_core_CipherKey[20]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_20_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_21_ ( .D(top_core_CipherKey[21]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_21_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_22_ ( .D(top_core_CipherKey[22]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_22_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_23_ ( .D(top_core_CipherKey[23]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_23_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_24_ ( .D(top_core_CipherKey[24]), .CK(
        n3694), .Q(top_core_KE_CipherKey0_24_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_25_ ( .D(top_core_CipherKey[25]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_25_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_26_ ( .D(top_core_CipherKey[26]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_26_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_27_ ( .D(top_core_CipherKey[27]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_27_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_28_ ( .D(top_core_CipherKey[28]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_28_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_29_ ( .D(top_core_CipherKey[29]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_29_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_30_ ( .D(top_core_CipherKey[30]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_30_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_31_ ( .D(top_core_CipherKey[31]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_31_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_32_ ( .D(top_core_CipherKey[32]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_32_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_33_ ( .D(top_core_CipherKey[33]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_33_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_34_ ( .D(top_core_CipherKey[34]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_34_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_35_ ( .D(top_core_CipherKey[35]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_35_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_36_ ( .D(top_core_CipherKey[36]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_36_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_37_ ( .D(top_core_CipherKey[37]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_37_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_38_ ( .D(top_core_CipherKey[38]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_38_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_39_ ( .D(top_core_CipherKey[39]), .CK(
        n3693), .Q(top_core_KE_CipherKey0_39_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_40_ ( .D(top_core_CipherKey[40]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_40_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_41_ ( .D(top_core_CipherKey[41]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_41_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_42_ ( .D(top_core_CipherKey[42]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_42_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_43_ ( .D(top_core_CipherKey[43]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_43_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_44_ ( .D(top_core_CipherKey[44]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_44_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_45_ ( .D(top_core_CipherKey[45]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_45_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_46_ ( .D(top_core_CipherKey[46]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_46_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_47_ ( .D(top_core_CipherKey[47]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_47_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_48_ ( .D(top_core_CipherKey[48]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_48_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_49_ ( .D(top_core_CipherKey[49]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_49_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_50_ ( .D(top_core_CipherKey[50]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_50_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_51_ ( .D(top_core_CipherKey[51]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_51_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_52_ ( .D(top_core_CipherKey[52]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_52_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_53_ ( .D(top_core_CipherKey[53]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_53_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_54_ ( .D(top_core_CipherKey[54]), .CK(
        n3692), .Q(top_core_KE_CipherKey0_54_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_55_ ( .D(top_core_CipherKey[55]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_55_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_56_ ( .D(top_core_CipherKey[56]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_56_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_57_ ( .D(top_core_CipherKey[57]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_57_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_58_ ( .D(top_core_CipherKey[58]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_58_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_59_ ( .D(top_core_CipherKey[59]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_59_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_60_ ( .D(top_core_CipherKey[60]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_60_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_61_ ( .D(top_core_CipherKey[61]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_61_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_62_ ( .D(top_core_CipherKey[62]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_62_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_39_ ( .D(top_core_KE_n4880), .CK(n3899), .Q(top_core_KE_prev_key1_reg_39_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_47_ ( .D(top_core_KE_n4872), .CK(n3898), .Q(top_core_KE_prev_key1_reg_47_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_55_ ( .D(top_core_KE_n4864), .CK(n3897), .Q(top_core_KE_prev_key1_reg_55_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_38_ ( .D(top_core_KE_n4881), .CK(n3903), .Q(top_core_KE_prev_key1_reg_38_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_46_ ( .D(top_core_KE_n4873), .CK(n3905), .Q(top_core_KE_prev_key1_reg_46_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_54_ ( .D(top_core_KE_n4865), .CK(n3893), .Q(top_core_KE_prev_key1_reg_54_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_53_ ( .D(top_core_KE_n4866), .CK(n3896), .Q(top_core_KE_prev_key1_reg_53_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_52_ ( .D(top_core_KE_n4867), .CK(n3893), .Q(top_core_KE_prev_key1_reg_52_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_51_ ( .D(top_core_KE_n4868), .CK(n3905), .Q(top_core_KE_prev_key1_reg_51_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_50_ ( .D(top_core_KE_n4869), .CK(n3902), .Q(top_core_KE_prev_key1_reg_50_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_49_ ( .D(top_core_KE_n4870), .CK(n3897), .Q(top_core_KE_prev_key1_reg_49_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_48_ ( .D(top_core_KE_n4871), .CK(n3897), .Q(top_core_KE_prev_key1_reg_48_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_37_ ( .D(top_core_KE_n4882), .CK(n3899), .Q(top_core_KE_prev_key1_reg_37_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_45_ ( .D(top_core_KE_n4874), .CK(n3900), .Q(top_core_KE_prev_key1_reg_45_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_36_ ( .D(top_core_KE_n4883), .CK(n3901), .Q(top_core_KE_prev_key1_reg_36_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_44_ ( .D(top_core_KE_n4875), .CK(n3902), .Q(top_core_KE_prev_key1_reg_44_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_35_ ( .D(top_core_KE_n4884), .CK(n3903), .Q(top_core_KE_prev_key1_reg_35_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_43_ ( .D(top_core_KE_n4876), .CK(n3904), .Q(top_core_KE_prev_key1_reg_43_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_34_ ( .D(top_core_KE_n4885), .CK(n3905), .Q(top_core_KE_prev_key1_reg_34_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_42_ ( .D(top_core_KE_n4877), .CK(n3906), .Q(top_core_KE_prev_key1_reg_42_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_33_ ( .D(top_core_KE_n4886), .CK(n3891), .Q(top_core_KE_prev_key1_reg_33_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_41_ ( .D(top_core_KE_n4878), .CK(n3892), .Q(top_core_KE_prev_key1_reg_41_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_32_ ( .D(top_core_KE_n4887), .CK(n3893), .Q(top_core_KE_prev_key1_reg_32_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_40_ ( .D(top_core_KE_n4879), .CK(n3894), .Q(top_core_KE_prev_key1_reg_40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__0_ ( .D(top_core_KE_n4664), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__1_ ( .D(top_core_KE_n4663), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__2_ ( .D(top_core_KE_n4662), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__3_ ( .D(top_core_KE_n4661), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__4_ ( .D(top_core_KE_n4660), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__5_ ( .D(top_core_KE_n4659), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__6_ ( .D(top_core_KE_n4658), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__7_ ( .D(top_core_KE_n4657), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__8_ ( .D(top_core_KE_n4656), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__9_ ( .D(top_core_KE_n4655), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__10_ ( .D(top_core_KE_n4654), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__11_ ( .D(top_core_KE_n4653), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__12_ ( .D(top_core_KE_n4652), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__13_ ( .D(top_core_KE_n4651), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__14_ ( .D(top_core_KE_n4650), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__15_ ( .D(top_core_KE_n4649), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__16_ ( .D(top_core_KE_n4648), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__17_ ( .D(top_core_KE_n4647), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__18_ ( .D(top_core_KE_n4646), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__19_ ( .D(top_core_KE_n4645), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__20_ ( .D(top_core_KE_n4644), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__21_ ( .D(top_core_KE_n4643), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__22_ ( .D(top_core_KE_n4642), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__23_ ( .D(top_core_KE_n4641), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__24_ ( .D(top_core_KE_n4640), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__25_ ( .D(top_core_KE_n4639), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__26_ ( .D(top_core_KE_n4638), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__27_ ( .D(top_core_KE_n4637), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__28_ ( .D(top_core_KE_n4636), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__29_ ( .D(top_core_KE_n4635), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__30_ ( .D(top_core_KE_n4634), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__31_ ( .D(top_core_KE_n4633), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__32_ ( .D(top_core_KE_n4632), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__33_ ( .D(top_core_KE_n4631), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__34_ ( .D(top_core_KE_n4630), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__35_ ( .D(top_core_KE_n4629), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__36_ ( .D(top_core_KE_n4628), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__37_ ( .D(top_core_KE_n4627), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__38_ ( .D(top_core_KE_n4626), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__39_ ( .D(top_core_KE_n4625), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__40_ ( .D(top_core_KE_n4624), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__41_ ( .D(top_core_KE_n4623), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__42_ ( .D(top_core_KE_n4622), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__43_ ( .D(top_core_KE_n4621), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__44_ ( .D(top_core_KE_n4620), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__45_ ( .D(top_core_KE_n4619), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__46_ ( .D(top_core_KE_n4618), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__47_ ( .D(top_core_KE_n4617), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__48_ ( .D(top_core_KE_n4616), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__49_ ( .D(top_core_KE_n4615), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__50_ ( .D(top_core_KE_n4614), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__51_ ( .D(top_core_KE_n4613), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__52_ ( .D(top_core_KE_n4612), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__53_ ( .D(top_core_KE_n4611), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__54_ ( .D(top_core_KE_n4610), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__55_ ( .D(top_core_KE_n4609), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__56_ ( .D(top_core_KE_n4608), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__57_ ( .D(top_core_KE_n4607), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__58_ ( .D(top_core_KE_n4606), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__59_ ( .D(top_core_KE_n4605), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__60_ ( .D(top_core_KE_n4604), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__61_ ( .D(top_core_KE_n4603), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__62_ ( .D(top_core_KE_n4602), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__63_ ( .D(top_core_KE_n4601), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__88_ ( .D(top_core_KE_n4576), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__89_ ( .D(top_core_KE_n4575), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__90_ ( .D(top_core_KE_n4574), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__91_ ( .D(top_core_KE_n4573), .CK(n3889), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__92_ ( .D(top_core_KE_n4572), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__93_ ( .D(top_core_KE_n4571), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__94_ ( .D(top_core_KE_n4570), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__95_ ( .D(top_core_KE_n4569), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__96_ ( .D(top_core_KE_n4568), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__97_ ( .D(top_core_KE_n4567), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__98_ ( .D(top_core_KE_n4566), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__99_ ( .D(top_core_KE_n4565), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__100_ ( .D(top_core_KE_n4564), .CK(n3877), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__101_ ( .D(top_core_KE_n4563), .CK(n3878), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__102_ ( .D(top_core_KE_n4562), .CK(n3879), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__103_ ( .D(top_core_KE_n4561), .CK(n3880), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__104_ ( .D(top_core_KE_n4560), .CK(n3881), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__105_ ( .D(top_core_KE_n4559), .CK(n3882), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__106_ ( .D(top_core_KE_n4558), .CK(n3883), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__107_ ( .D(top_core_KE_n4557), .CK(n3817), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__108_ ( .D(top_core_KE_n4556), .CK(n3818), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__109_ ( .D(top_core_KE_n4555), .CK(n3819), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__110_ ( .D(top_core_KE_n4554), .CK(n3820), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__111_ ( .D(top_core_KE_n4553), .CK(n3821), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__120_ ( .D(top_core_KE_n4544), .CK(n3821), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__121_ ( .D(top_core_KE_n4543), .CK(n3822), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__122_ ( .D(top_core_KE_n4542), .CK(n3823), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__123_ ( .D(top_core_KE_n4541), .CK(n3824), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__124_ ( .D(top_core_KE_n4540), .CK(n3825), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__125_ ( .D(top_core_KE_n4539), .CK(n3826), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__126_ ( .D(top_core_KE_n4538), .CK(n3827), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__71_ ( .D(top_core_KE_n4593), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__79_ ( .D(top_core_KE_n4585), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__119_ ( .D(top_core_KE_n4545), .CK(n3809), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__87_ ( .D(top_core_KE_n4577), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__127_ ( .D(top_core_KE_n4537), .CK(n3810), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__70_ ( .D(top_core_KE_n4594), .CK(n3811), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__78_ ( .D(top_core_KE_n4586), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__118_ ( .D(top_core_KE_n4546), .CK(n3813), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__86_ ( .D(top_core_KE_n4578), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__117_ ( .D(top_core_KE_n4547), .CK(n3815), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__85_ ( .D(top_core_KE_n4579), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__116_ ( .D(top_core_KE_n4548), .CK(n3817), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__84_ ( .D(top_core_KE_n4580), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__115_ ( .D(top_core_KE_n4549), .CK(n3839), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__83_ ( .D(top_core_KE_n4581), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__114_ ( .D(top_core_KE_n4550), .CK(n3841), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__82_ ( .D(top_core_KE_n4582), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__113_ ( .D(top_core_KE_n4551), .CK(n3842), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__81_ ( .D(top_core_KE_n4583), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__112_ ( .D(top_core_KE_n4552), .CK(n3844), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__80_ ( .D(top_core_KE_n4584), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__69_ ( .D(top_core_KE_n4595), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__77_ ( .D(top_core_KE_n4587), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__68_ ( .D(top_core_KE_n4596), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__76_ ( .D(top_core_KE_n4588), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__67_ ( .D(top_core_KE_n4597), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__75_ ( .D(top_core_KE_n4589), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__66_ ( .D(top_core_KE_n4598), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__74_ ( .D(top_core_KE_n4590), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__65_ ( .D(top_core_KE_n4599), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__73_ ( .D(top_core_KE_n4591), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__64_ ( .D(top_core_KE_n4600), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__72_ ( .D(top_core_KE_n4592), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_14__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_14__128_ ( .D(top_core_KE_n4536), .CK(n3836), .RN(n_RSTB), .Q(top_core_KE_key_mem_14__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__0_ ( .D(top_core_KE_n4535), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__1_ ( .D(top_core_KE_n4534), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__2_ ( .D(top_core_KE_n4533), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__3_ ( .D(top_core_KE_n4532), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__4_ ( .D(top_core_KE_n4531), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__5_ ( .D(top_core_KE_n4530), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__6_ ( .D(top_core_KE_n4529), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__7_ ( .D(top_core_KE_n4528), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__8_ ( .D(top_core_KE_n4527), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__9_ ( .D(top_core_KE_n4526), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__10_ ( .D(top_core_KE_n4525), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__11_ ( .D(top_core_KE_n4524), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__12_ ( .D(top_core_KE_n4523), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__13_ ( .D(top_core_KE_n4522), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__14_ ( .D(top_core_KE_n4521), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__15_ ( .D(top_core_KE_n4520), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__16_ ( .D(top_core_KE_n4519), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__17_ ( .D(top_core_KE_n4518), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__18_ ( .D(top_core_KE_n4517), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__19_ ( .D(top_core_KE_n4516), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__20_ ( .D(top_core_KE_n4515), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__21_ ( .D(top_core_KE_n4514), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__22_ ( .D(top_core_KE_n4513), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__23_ ( .D(top_core_KE_n4512), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__24_ ( .D(top_core_KE_n4511), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__25_ ( .D(top_core_KE_n4510), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__26_ ( .D(top_core_KE_n4509), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__27_ ( .D(top_core_KE_n4508), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__28_ ( .D(top_core_KE_n4507), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__29_ ( .D(top_core_KE_n4506), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__30_ ( .D(top_core_KE_n4505), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__31_ ( .D(top_core_KE_n4504), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__32_ ( .D(top_core_KE_n4503), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__33_ ( .D(top_core_KE_n4502), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__34_ ( .D(top_core_KE_n4501), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__35_ ( .D(top_core_KE_n4500), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__36_ ( .D(top_core_KE_n4499), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__37_ ( .D(top_core_KE_n4498), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__38_ ( .D(top_core_KE_n4497), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__39_ ( .D(top_core_KE_n4496), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__40_ ( .D(top_core_KE_n4495), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__41_ ( .D(top_core_KE_n4494), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__42_ ( .D(top_core_KE_n4493), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__43_ ( .D(top_core_KE_n4492), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__44_ ( .D(top_core_KE_n4491), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__45_ ( .D(top_core_KE_n4490), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__46_ ( .D(top_core_KE_n4489), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__47_ ( .D(top_core_KE_n4488), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__48_ ( .D(top_core_KE_n4487), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__49_ ( .D(top_core_KE_n4486), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__50_ ( .D(top_core_KE_n4485), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__51_ ( .D(top_core_KE_n4484), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__52_ ( .D(top_core_KE_n4483), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__53_ ( .D(top_core_KE_n4482), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__54_ ( .D(top_core_KE_n4481), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__55_ ( .D(top_core_KE_n4480), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__56_ ( .D(top_core_KE_n4479), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__57_ ( .D(top_core_KE_n4478), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__58_ ( .D(top_core_KE_n4477), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__59_ ( .D(top_core_KE_n4476), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__60_ ( .D(top_core_KE_n4475), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__61_ ( .D(top_core_KE_n4474), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__62_ ( .D(top_core_KE_n4473), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__63_ ( .D(top_core_KE_n4472), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__88_ ( .D(top_core_KE_n4447), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__89_ ( .D(top_core_KE_n4446), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__90_ ( .D(top_core_KE_n4445), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__91_ ( .D(top_core_KE_n4444), .CK(n3889), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__92_ ( .D(top_core_KE_n4443), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__93_ ( .D(top_core_KE_n4442), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__94_ ( .D(top_core_KE_n4441), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__95_ ( .D(top_core_KE_n4440), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__96_ ( .D(top_core_KE_n4439), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__97_ ( .D(top_core_KE_n4438), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__98_ ( .D(top_core_KE_n4437), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__99_ ( .D(top_core_KE_n4436), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__100_ ( .D(top_core_KE_n4435), .CK(n3878), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__101_ ( .D(top_core_KE_n4434), .CK(n3878), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__102_ ( .D(top_core_KE_n4433), .CK(n3879), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__103_ ( .D(top_core_KE_n4432), .CK(n3880), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__104_ ( .D(top_core_KE_n4431), .CK(n3881), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__105_ ( .D(top_core_KE_n4430), .CK(n3882), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__106_ ( .D(top_core_KE_n4429), .CK(n3883), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__107_ ( .D(top_core_KE_n4428), .CK(n3817), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__108_ ( .D(top_core_KE_n4427), .CK(n3818), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__109_ ( .D(top_core_KE_n4426), .CK(n3819), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__110_ ( .D(top_core_KE_n4425), .CK(n3820), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__111_ ( .D(top_core_KE_n4424), .CK(n3821), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__120_ ( .D(top_core_KE_n4415), .CK(n3822), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__121_ ( .D(top_core_KE_n4414), .CK(n3822), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__122_ ( .D(top_core_KE_n4413), .CK(n3823), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__123_ ( .D(top_core_KE_n4412), .CK(n3824), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__124_ ( .D(top_core_KE_n4411), .CK(n3825), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__125_ ( .D(top_core_KE_n4410), .CK(n3826), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__126_ ( .D(top_core_KE_n4409), .CK(n3827), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__71_ ( .D(top_core_KE_n4464), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__79_ ( .D(top_core_KE_n4456), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__119_ ( .D(top_core_KE_n4416), .CK(n3809), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__87_ ( .D(top_core_KE_n4448), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__127_ ( .D(top_core_KE_n4408), .CK(n3811), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__70_ ( .D(top_core_KE_n4465), .CK(n3811), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__78_ ( .D(top_core_KE_n4457), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__118_ ( .D(top_core_KE_n4417), .CK(n3813), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__86_ ( .D(top_core_KE_n4449), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__117_ ( .D(top_core_KE_n4418), .CK(n3815), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__85_ ( .D(top_core_KE_n4450), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__116_ ( .D(top_core_KE_n4419), .CK(n3842), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__84_ ( .D(top_core_KE_n4451), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__115_ ( .D(top_core_KE_n4420), .CK(n3839), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__83_ ( .D(top_core_KE_n4452), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__114_ ( .D(top_core_KE_n4421), .CK(n3841), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__82_ ( .D(top_core_KE_n4453), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__113_ ( .D(top_core_KE_n4422), .CK(n3843), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__81_ ( .D(top_core_KE_n4454), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__112_ ( .D(top_core_KE_n4423), .CK(n3844), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__80_ ( .D(top_core_KE_n4455), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__69_ ( .D(top_core_KE_n4466), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__77_ ( .D(top_core_KE_n4458), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__68_ ( .D(top_core_KE_n4467), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__76_ ( .D(top_core_KE_n4459), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__67_ ( .D(top_core_KE_n4468), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__75_ ( .D(top_core_KE_n4460), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__66_ ( .D(top_core_KE_n4469), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__74_ ( .D(top_core_KE_n4461), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__65_ ( .D(top_core_KE_n4470), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__73_ ( .D(top_core_KE_n4462), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__64_ ( .D(top_core_KE_n4471), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__72_ ( .D(top_core_KE_n4463), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_13__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_13__128_ ( .D(top_core_KE_n4407), .CK(n3836), .RN(n_RSTB), .Q(top_core_KE_key_mem_13__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__0_ ( .D(top_core_KE_n4019), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__1_ ( .D(top_core_KE_n4018), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__2_ ( .D(top_core_KE_n4017), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__3_ ( .D(top_core_KE_n4016), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__4_ ( .D(top_core_KE_n4015), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__5_ ( .D(top_core_KE_n4014), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__6_ ( .D(top_core_KE_n4013), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__7_ ( .D(top_core_KE_n4012), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__8_ ( .D(top_core_KE_n4011), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__9_ ( .D(top_core_KE_n4010), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__10_ ( .D(top_core_KE_n4009), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__11_ ( .D(top_core_KE_n4008), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__12_ ( .D(top_core_KE_n4007), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__13_ ( .D(top_core_KE_n4006), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__14_ ( .D(top_core_KE_n4005), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__15_ ( .D(top_core_KE_n4004), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__16_ ( .D(top_core_KE_n4003), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__17_ ( .D(top_core_KE_n4002), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__18_ ( .D(top_core_KE_n4001), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__19_ ( .D(top_core_KE_n4000), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__20_ ( .D(top_core_KE_n3999), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__21_ ( .D(top_core_KE_n3998), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__22_ ( .D(top_core_KE_n3997), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__23_ ( .D(top_core_KE_n3996), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__24_ ( .D(top_core_KE_n3995), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__25_ ( .D(top_core_KE_n3994), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__26_ ( .D(top_core_KE_n3993), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__27_ ( .D(top_core_KE_n3992), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__28_ ( .D(top_core_KE_n3991), .CK(n3723), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__29_ ( .D(top_core_KE_n3990), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__30_ ( .D(top_core_KE_n3989), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__31_ ( .D(top_core_KE_n3988), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__32_ ( .D(top_core_KE_n3987), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__33_ ( .D(top_core_KE_n3986), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__34_ ( .D(top_core_KE_n3985), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__35_ ( .D(top_core_KE_n3984), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__36_ ( .D(top_core_KE_n3983), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__37_ ( .D(top_core_KE_n3982), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__38_ ( .D(top_core_KE_n3981), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__39_ ( .D(top_core_KE_n3980), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__40_ ( .D(top_core_KE_n3979), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__41_ ( .D(top_core_KE_n3978), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__42_ ( .D(top_core_KE_n3977), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__43_ ( .D(top_core_KE_n3976), .CK(n3724), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__44_ ( .D(top_core_KE_n3975), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__45_ ( .D(top_core_KE_n3974), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__46_ ( .D(top_core_KE_n3973), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__47_ ( .D(top_core_KE_n3972), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__48_ ( .D(top_core_KE_n3971), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__49_ ( .D(top_core_KE_n3970), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__50_ ( .D(top_core_KE_n3969), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__51_ ( .D(top_core_KE_n3968), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__52_ ( .D(top_core_KE_n3967), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__53_ ( .D(top_core_KE_n3966), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__54_ ( .D(top_core_KE_n3965), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__55_ ( .D(top_core_KE_n3964), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__56_ ( .D(top_core_KE_n3963), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__57_ ( .D(top_core_KE_n3962), .CK(n3725), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__58_ ( .D(top_core_KE_n3961), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__59_ ( .D(top_core_KE_n3960), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__60_ ( .D(top_core_KE_n3959), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__61_ ( .D(top_core_KE_n3958), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__62_ ( .D(top_core_KE_n3957), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__63_ ( .D(top_core_KE_n3956), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__64_ ( .D(top_core_KE_n3955), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__65_ ( .D(top_core_KE_n3954), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__66_ ( .D(top_core_KE_n3953), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__67_ ( .D(top_core_KE_n3952), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__68_ ( .D(top_core_KE_n3951), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__69_ ( .D(top_core_KE_n3950), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__70_ ( .D(top_core_KE_n3949), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__71_ ( .D(top_core_KE_n3948), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__72_ ( .D(top_core_KE_n3947), .CK(n3726), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__73_ ( .D(top_core_KE_n3946), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__74_ ( .D(top_core_KE_n3945), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__75_ ( .D(top_core_KE_n3944), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__76_ ( .D(top_core_KE_n3943), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__77_ ( .D(top_core_KE_n3942), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__78_ ( .D(top_core_KE_n3941), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__79_ ( .D(top_core_KE_n3940), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__80_ ( .D(top_core_KE_n3939), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__81_ ( .D(top_core_KE_n3938), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__82_ ( .D(top_core_KE_n3937), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__83_ ( .D(top_core_KE_n3936), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__84_ ( .D(top_core_KE_n3935), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__85_ ( .D(top_core_KE_n3934), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__86_ ( .D(top_core_KE_n3933), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__87_ ( .D(top_core_KE_n3932), .CK(n3727), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__88_ ( .D(top_core_KE_n3931), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__89_ ( .D(top_core_KE_n3930), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__90_ ( .D(top_core_KE_n3929), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__91_ ( .D(top_core_KE_n3928), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__92_ ( .D(top_core_KE_n3927), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__93_ ( .D(top_core_KE_n3926), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__94_ ( .D(top_core_KE_n3925), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__95_ ( .D(top_core_KE_n3924), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__96_ ( .D(top_core_KE_n3923), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__97_ ( .D(top_core_KE_n3922), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__98_ ( .D(top_core_KE_n3921), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__99_ ( .D(top_core_KE_n3920), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__100_ ( .D(top_core_KE_n3919), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__101_ ( .D(top_core_KE_n3918), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__102_ ( .D(top_core_KE_n3917), .CK(n3728), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__103_ ( .D(top_core_KE_n3916), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__104_ ( .D(top_core_KE_n3915), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__105_ ( .D(top_core_KE_n3914), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__106_ ( .D(top_core_KE_n3913), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__107_ ( .D(top_core_KE_n3912), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__108_ ( .D(top_core_KE_n3911), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__109_ ( .D(top_core_KE_n3910), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__110_ ( .D(top_core_KE_n3909), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__111_ ( .D(top_core_KE_n3908), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__112_ ( .D(top_core_KE_n3907), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__113_ ( .D(top_core_KE_n3906), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__114_ ( .D(top_core_KE_n3905), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__115_ ( .D(top_core_KE_n3904), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__116_ ( .D(top_core_KE_n3903), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__117_ ( .D(top_core_KE_n3902), .CK(n3729), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__118_ ( .D(top_core_KE_n3901), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__119_ ( .D(top_core_KE_n3900), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__120_ ( .D(top_core_KE_n3899), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__121_ ( .D(top_core_KE_n3898), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__122_ ( .D(top_core_KE_n3897), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__123_ ( .D(top_core_KE_n3896), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__124_ ( .D(top_core_KE_n3895), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__125_ ( .D(top_core_KE_n3894), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__126_ ( .D(top_core_KE_n3893), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__127_ ( .D(top_core_KE_n3892), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_9__128_ ( .D(top_core_KE_n3891), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_9__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__0_ ( .D(top_core_KE_n3503), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__0_ ( .D(top_core_KE_n2987), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__1_ ( .D(top_core_KE_n3502), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__1_ ( .D(top_core_KE_n2986), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__2_ ( .D(top_core_KE_n3501), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__2_ ( .D(top_core_KE_n2985), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__3_ ( .D(top_core_KE_n3500), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__3_ ( .D(top_core_KE_n2984), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__4_ ( .D(top_core_KE_n3499), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__4_ ( .D(top_core_KE_n2983), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__5_ ( .D(top_core_KE_n3498), .CK(n3719), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__5_ ( .D(top_core_KE_n2982), .CK(n3719), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__6_ ( .D(top_core_KE_n3497), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__6_ ( .D(top_core_KE_n2981), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__7_ ( .D(top_core_KE_n3496), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__7_ ( .D(top_core_KE_n2980), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__8_ ( .D(top_core_KE_n3495), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__8_ ( .D(top_core_KE_n2979), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__9_ ( .D(top_core_KE_n3494), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__9_ ( .D(top_core_KE_n2978), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__10_ ( .D(top_core_KE_n3493), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__10_ ( .D(top_core_KE_n2977), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__11_ ( .D(top_core_KE_n3492), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__11_ ( .D(top_core_KE_n2976), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__12_ ( .D(top_core_KE_n3491), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__12_ ( .D(top_core_KE_n2975), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__13_ ( .D(top_core_KE_n3490), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__13_ ( .D(top_core_KE_n2974), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__14_ ( .D(top_core_KE_n3489), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__14_ ( .D(top_core_KE_n2973), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__15_ ( .D(top_core_KE_n3488), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__15_ ( .D(top_core_KE_n2972), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__16_ ( .D(top_core_KE_n3487), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__16_ ( .D(top_core_KE_n2971), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__17_ ( .D(top_core_KE_n3486), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__17_ ( .D(top_core_KE_n2970), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__18_ ( .D(top_core_KE_n3485), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__18_ ( .D(top_core_KE_n2969), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__19_ ( .D(top_core_KE_n3484), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__19_ ( .D(top_core_KE_n2968), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__20_ ( .D(top_core_KE_n3483), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__20_ ( .D(top_core_KE_n2967), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__21_ ( .D(top_core_KE_n3482), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__21_ ( .D(top_core_KE_n2966), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__22_ ( .D(top_core_KE_n3481), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__22_ ( .D(top_core_KE_n2965), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__23_ ( .D(top_core_KE_n3480), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__23_ ( .D(top_core_KE_n2964), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__24_ ( .D(top_core_KE_n3479), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__24_ ( .D(top_core_KE_n2963), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__25_ ( .D(top_core_KE_n3478), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__25_ ( .D(top_core_KE_n2962), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__26_ ( .D(top_core_KE_n3477), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__26_ ( .D(top_core_KE_n2961), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__27_ ( .D(top_core_KE_n3476), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__27_ ( .D(top_core_KE_n2960), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__28_ ( .D(top_core_KE_n3475), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__28_ ( .D(top_core_KE_n2959), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__29_ ( .D(top_core_KE_n3474), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__29_ ( .D(top_core_KE_n2958), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__30_ ( .D(top_core_KE_n3473), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__30_ ( .D(top_core_KE_n2957), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__31_ ( .D(top_core_KE_n3472), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__31_ ( .D(top_core_KE_n2956), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__32_ ( .D(top_core_KE_n3471), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__32_ ( .D(top_core_KE_n2955), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__33_ ( .D(top_core_KE_n3470), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__33_ ( .D(top_core_KE_n2954), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__34_ ( .D(top_core_KE_n3469), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__34_ ( .D(top_core_KE_n2953), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__35_ ( .D(top_core_KE_n3468), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__35_ ( .D(top_core_KE_n2952), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__36_ ( .D(top_core_KE_n3467), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__36_ ( .D(top_core_KE_n2951), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__37_ ( .D(top_core_KE_n3466), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__37_ ( .D(top_core_KE_n2950), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__38_ ( .D(top_core_KE_n3465), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__38_ ( .D(top_core_KE_n2949), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__39_ ( .D(top_core_KE_n3464), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__39_ ( .D(top_core_KE_n2948), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__40_ ( .D(top_core_KE_n3463), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__40_ ( .D(top_core_KE_n2947), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__41_ ( .D(top_core_KE_n3462), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__41_ ( .D(top_core_KE_n2946), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__42_ ( .D(top_core_KE_n3461), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__42_ ( .D(top_core_KE_n2945), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__43_ ( .D(top_core_KE_n3460), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__43_ ( .D(top_core_KE_n2944), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__44_ ( .D(top_core_KE_n3459), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__44_ ( .D(top_core_KE_n2943), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__45_ ( .D(top_core_KE_n3458), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__45_ ( .D(top_core_KE_n2942), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__46_ ( .D(top_core_KE_n3457), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__46_ ( .D(top_core_KE_n2941), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__47_ ( .D(top_core_KE_n3456), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__47_ ( .D(top_core_KE_n2940), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__48_ ( .D(top_core_KE_n3455), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__48_ ( .D(top_core_KE_n2939), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__49_ ( .D(top_core_KE_n3454), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__49_ ( .D(top_core_KE_n2938), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__50_ ( .D(top_core_KE_n3453), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__50_ ( .D(top_core_KE_n2937), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__51_ ( .D(top_core_KE_n3452), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__51_ ( .D(top_core_KE_n2936), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__52_ ( .D(top_core_KE_n3451), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__52_ ( .D(top_core_KE_n2935), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__53_ ( .D(top_core_KE_n3450), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__53_ ( .D(top_core_KE_n2934), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__54_ ( .D(top_core_KE_n3449), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__54_ ( .D(top_core_KE_n2933), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__55_ ( .D(top_core_KE_n3448), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__55_ ( .D(top_core_KE_n2932), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__56_ ( .D(top_core_KE_n3447), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__56_ ( .D(top_core_KE_n2931), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__57_ ( .D(top_core_KE_n3446), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__57_ ( .D(top_core_KE_n2930), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__58_ ( .D(top_core_KE_n3445), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__58_ ( .D(top_core_KE_n2929), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__59_ ( .D(top_core_KE_n3444), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__59_ ( .D(top_core_KE_n2928), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__60_ ( .D(top_core_KE_n3443), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__60_ ( .D(top_core_KE_n2927), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__61_ ( .D(top_core_KE_n3442), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__61_ ( .D(top_core_KE_n2926), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__62_ ( .D(top_core_KE_n3441), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__62_ ( .D(top_core_KE_n2925), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__63_ ( .D(top_core_KE_n3440), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__63_ ( .D(top_core_KE_n2924), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__88_ ( .D(top_core_KE_n3415), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__88_ ( .D(top_core_KE_n2899), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__89_ ( .D(top_core_KE_n3414), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__89_ ( .D(top_core_KE_n2898), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__90_ ( .D(top_core_KE_n3413), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__90_ ( .D(top_core_KE_n2897), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__91_ ( .D(top_core_KE_n3412), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__91_ ( .D(top_core_KE_n2896), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__92_ ( .D(top_core_KE_n3411), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__92_ ( .D(top_core_KE_n2895), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__93_ ( .D(top_core_KE_n3410), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__93_ ( .D(top_core_KE_n2894), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__94_ ( .D(top_core_KE_n3409), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__94_ ( .D(top_core_KE_n2893), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__95_ ( .D(top_core_KE_n3408), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__95_ ( .D(top_core_KE_n2892), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__96_ ( .D(top_core_KE_n3407), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__96_ ( .D(top_core_KE_n2891), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__97_ ( .D(top_core_KE_n3406), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__97_ ( .D(top_core_KE_n2890), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__98_ ( .D(top_core_KE_n3405), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__98_ ( .D(top_core_KE_n2889), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__99_ ( .D(top_core_KE_n3404), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__99_ ( .D(top_core_KE_n2888), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__100_ ( .D(top_core_KE_n3403), .CK(n3878), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__100_ ( .D(top_core_KE_n2887), .CK(n3878), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__101_ ( .D(top_core_KE_n3402), .CK(n3879), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__101_ ( .D(top_core_KE_n2886), .CK(n3879), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__102_ ( .D(top_core_KE_n3401), .CK(n3880), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__102_ ( .D(top_core_KE_n2885), .CK(n3880), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__103_ ( .D(top_core_KE_n3400), .CK(n3881), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__103_ ( .D(top_core_KE_n2884), .CK(n3881), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__104_ ( .D(top_core_KE_n3399), .CK(n3881), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__104_ ( .D(top_core_KE_n2883), .CK(n3882), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__105_ ( .D(top_core_KE_n3398), .CK(n3882), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__105_ ( .D(top_core_KE_n2882), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__106_ ( .D(top_core_KE_n3397), .CK(n3817), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__106_ ( .D(top_core_KE_n2881), .CK(n3817), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__107_ ( .D(top_core_KE_n3396), .CK(n3818), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__107_ ( .D(top_core_KE_n2880), .CK(n3818), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__108_ ( .D(top_core_KE_n3395), .CK(n3818), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__108_ ( .D(top_core_KE_n2879), .CK(n3819), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__109_ ( .D(top_core_KE_n3394), .CK(n3819), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__109_ ( .D(top_core_KE_n2878), .CK(n3820), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__110_ ( .D(top_core_KE_n3393), .CK(n3820), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__110_ ( .D(top_core_KE_n2877), .CK(n3820), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__111_ ( .D(top_core_KE_n3392), .CK(n3821), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__111_ ( .D(top_core_KE_n2876), .CK(n3821), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__120_ ( .D(top_core_KE_n3383), .CK(n3822), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__120_ ( .D(top_core_KE_n2867), .CK(n3822), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__121_ ( .D(top_core_KE_n3382), .CK(n3823), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__121_ ( .D(top_core_KE_n2866), .CK(n3823), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__122_ ( .D(top_core_KE_n3381), .CK(n3824), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__122_ ( .D(top_core_KE_n2865), .CK(n3824), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__123_ ( .D(top_core_KE_n3380), .CK(n3825), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__123_ ( .D(top_core_KE_n2864), .CK(n3825), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__124_ ( .D(top_core_KE_n3379), .CK(n3825), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__124_ ( .D(top_core_KE_n2863), .CK(n3826), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__125_ ( .D(top_core_KE_n3378), .CK(n3826), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__125_ ( .D(top_core_KE_n2862), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__126_ ( .D(top_core_KE_n3377), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__126_ ( .D(top_core_KE_n2861), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__71_ ( .D(top_core_KE_n3432), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__71_ ( .D(top_core_KE_n2916), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__79_ ( .D(top_core_KE_n3424), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__79_ ( .D(top_core_KE_n2908), .CK(n3809), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__119_ ( .D(top_core_KE_n3384), .CK(n3809), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__119_ ( .D(top_core_KE_n2868), .CK(n3809), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__87_ ( .D(top_core_KE_n3416), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__87_ ( .D(top_core_KE_n2900), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__127_ ( .D(top_core_KE_n3376), .CK(n3811), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__127_ ( .D(top_core_KE_n2860), .CK(n3811), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__70_ ( .D(top_core_KE_n3433), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__70_ ( .D(top_core_KE_n2917), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__78_ ( .D(top_core_KE_n3425), .CK(n3813), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__78_ ( .D(top_core_KE_n2909), .CK(n3813), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__118_ ( .D(top_core_KE_n3385), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__118_ ( .D(top_core_KE_n2869), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__86_ ( .D(top_core_KE_n3417), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__86_ ( .D(top_core_KE_n2901), .CK(n3815), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__117_ ( .D(top_core_KE_n3386), .CK(n3815), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__117_ ( .D(top_core_KE_n2870), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__85_ ( .D(top_core_KE_n3418), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__85_ ( .D(top_core_KE_n2902), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__116_ ( .D(top_core_KE_n3387), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__116_ ( .D(top_core_KE_n2871), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__84_ ( .D(top_core_KE_n3419), .CK(n3839), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__84_ ( .D(top_core_KE_n2903), .CK(n3839), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__115_ ( .D(top_core_KE_n3388), .CK(n3839), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__115_ ( .D(top_core_KE_n2872), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__83_ ( .D(top_core_KE_n3420), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__83_ ( .D(top_core_KE_n2904), .CK(n3841), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__114_ ( .D(top_core_KE_n3389), .CK(n3841), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__114_ ( .D(top_core_KE_n2873), .CK(n3841), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__82_ ( .D(top_core_KE_n3421), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__82_ ( .D(top_core_KE_n2905), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__113_ ( .D(top_core_KE_n3390), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__113_ ( .D(top_core_KE_n2874), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__81_ ( .D(top_core_KE_n3422), .CK(n3844), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__81_ ( .D(top_core_KE_n2906), .CK(n3844), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__112_ ( .D(top_core_KE_n3391), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__112_ ( .D(top_core_KE_n2875), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__80_ ( .D(top_core_KE_n3423), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__80_ ( .D(top_core_KE_n2907), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__69_ ( .D(top_core_KE_n3434), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__69_ ( .D(top_core_KE_n2918), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__77_ ( .D(top_core_KE_n3426), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__77_ ( .D(top_core_KE_n2910), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__68_ ( .D(top_core_KE_n3435), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__68_ ( .D(top_core_KE_n2919), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__76_ ( .D(top_core_KE_n3427), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__76_ ( .D(top_core_KE_n2911), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__67_ ( .D(top_core_KE_n3436), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__67_ ( .D(top_core_KE_n2920), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__75_ ( .D(top_core_KE_n3428), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__75_ ( .D(top_core_KE_n2912), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__66_ ( .D(top_core_KE_n3437), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__66_ ( .D(top_core_KE_n2921), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__74_ ( .D(top_core_KE_n3429), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__74_ ( .D(top_core_KE_n2913), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__65_ ( .D(top_core_KE_n3438), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__65_ ( .D(top_core_KE_n2922), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__73_ ( .D(top_core_KE_n3430), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__73_ ( .D(top_core_KE_n2914), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__64_ ( .D(top_core_KE_n3439), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__64_ ( .D(top_core_KE_n2923), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__72_ ( .D(top_core_KE_n3431), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__72_ ( .D(top_core_KE_n2915), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_1__128_ ( .D(top_core_KE_n2859), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_1__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_5__128_ ( .D(top_core_KE_n3375), .CK(n3837), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_5__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__0_ ( .D(top_core_KE_n4277), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__0_ ( .D(top_core_KE_n3761), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__0_ ( .D(top_core_KE_n3245), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__1_ ( .D(top_core_KE_n4276), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__1_ ( .D(top_core_KE_n3760), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__1_ ( .D(top_core_KE_n3244), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__2_ ( .D(top_core_KE_n4275), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__2_ ( .D(top_core_KE_n3759), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__2_ ( .D(top_core_KE_n3243), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__3_ ( .D(top_core_KE_n4274), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__3_ ( .D(top_core_KE_n3758), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__3_ ( .D(top_core_KE_n3242), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__4_ ( .D(top_core_KE_n4273), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__4_ ( .D(top_core_KE_n3757), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__4_ ( .D(top_core_KE_n3241), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__5_ ( .D(top_core_KE_n4272), .CK(n3719), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__5_ ( .D(top_core_KE_n3756), .CK(n3719), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__5_ ( .D(top_core_KE_n3240), .CK(n3719), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__6_ ( .D(top_core_KE_n4271), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__6_ ( .D(top_core_KE_n3755), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__6_ ( .D(top_core_KE_n3239), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__7_ ( .D(top_core_KE_n4270), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__7_ ( .D(top_core_KE_n3754), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__7_ ( .D(top_core_KE_n3238), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__8_ ( .D(top_core_KE_n4269), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__8_ ( .D(top_core_KE_n3753), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__8_ ( .D(top_core_KE_n3237), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__9_ ( .D(top_core_KE_n4268), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__9_ ( .D(top_core_KE_n3752), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__9_ ( .D(top_core_KE_n3236), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__10_ ( .D(top_core_KE_n4267), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__10_ ( .D(top_core_KE_n3751), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__10_ ( .D(top_core_KE_n3235), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__11_ ( .D(top_core_KE_n4266), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__11_ ( .D(top_core_KE_n3750), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__11_ ( .D(top_core_KE_n3234), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__12_ ( .D(top_core_KE_n4265), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__12_ ( .D(top_core_KE_n3749), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__12_ ( .D(top_core_KE_n3233), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__13_ ( .D(top_core_KE_n4264), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__13_ ( .D(top_core_KE_n3748), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__13_ ( .D(top_core_KE_n3232), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__14_ ( .D(top_core_KE_n4263), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__14_ ( .D(top_core_KE_n3747), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__14_ ( .D(top_core_KE_n3231), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__15_ ( .D(top_core_KE_n4262), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__15_ ( .D(top_core_KE_n3746), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__15_ ( .D(top_core_KE_n3230), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__16_ ( .D(top_core_KE_n4261), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__16_ ( .D(top_core_KE_n3745), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__16_ ( .D(top_core_KE_n3229), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__17_ ( .D(top_core_KE_n4260), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__17_ ( .D(top_core_KE_n3744), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__17_ ( .D(top_core_KE_n3228), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__18_ ( .D(top_core_KE_n4259), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__18_ ( .D(top_core_KE_n3743), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__18_ ( .D(top_core_KE_n3227), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__19_ ( .D(top_core_KE_n4258), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__19_ ( .D(top_core_KE_n3742), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__19_ ( .D(top_core_KE_n3226), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__20_ ( .D(top_core_KE_n4257), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__20_ ( .D(top_core_KE_n3741), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__20_ ( .D(top_core_KE_n3225), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__21_ ( .D(top_core_KE_n4256), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__21_ ( .D(top_core_KE_n3740), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__21_ ( .D(top_core_KE_n3224), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__22_ ( .D(top_core_KE_n4255), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__22_ ( .D(top_core_KE_n3739), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__22_ ( .D(top_core_KE_n3223), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__23_ ( .D(top_core_KE_n4254), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__23_ ( .D(top_core_KE_n3738), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__23_ ( .D(top_core_KE_n3222), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__24_ ( .D(top_core_KE_n4253), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__24_ ( .D(top_core_KE_n3737), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__24_ ( .D(top_core_KE_n3221), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__25_ ( .D(top_core_KE_n4252), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__25_ ( .D(top_core_KE_n3736), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__25_ ( .D(top_core_KE_n3220), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__26_ ( .D(top_core_KE_n4251), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__26_ ( .D(top_core_KE_n3735), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__26_ ( .D(top_core_KE_n3219), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__27_ ( .D(top_core_KE_n4250), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__27_ ( .D(top_core_KE_n3734), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__27_ ( .D(top_core_KE_n3218), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__28_ ( .D(top_core_KE_n4249), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__28_ ( .D(top_core_KE_n3733), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__28_ ( .D(top_core_KE_n3217), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__29_ ( .D(top_core_KE_n4248), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__29_ ( .D(top_core_KE_n3732), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__29_ ( .D(top_core_KE_n3216), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__30_ ( .D(top_core_KE_n4247), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__30_ ( .D(top_core_KE_n3731), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__30_ ( .D(top_core_KE_n3215), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__31_ ( .D(top_core_KE_n4246), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__31_ ( .D(top_core_KE_n3730), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__31_ ( .D(top_core_KE_n3214), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__32_ ( .D(top_core_KE_n4245), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__32_ ( .D(top_core_KE_n3729), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__32_ ( .D(top_core_KE_n3213), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__33_ ( .D(top_core_KE_n4244), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__33_ ( .D(top_core_KE_n3728), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__33_ ( .D(top_core_KE_n3212), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__34_ ( .D(top_core_KE_n4243), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__34_ ( .D(top_core_KE_n3727), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__34_ ( .D(top_core_KE_n3211), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__35_ ( .D(top_core_KE_n4242), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__35_ ( .D(top_core_KE_n3726), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__35_ ( .D(top_core_KE_n3210), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__36_ ( .D(top_core_KE_n4241), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__36_ ( .D(top_core_KE_n3725), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__36_ ( .D(top_core_KE_n3209), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__37_ ( .D(top_core_KE_n4240), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__37_ ( .D(top_core_KE_n3724), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__37_ ( .D(top_core_KE_n3208), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__38_ ( .D(top_core_KE_n4239), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__38_ ( .D(top_core_KE_n3723), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__38_ ( .D(top_core_KE_n3207), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__39_ ( .D(top_core_KE_n4238), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__39_ ( .D(top_core_KE_n3722), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__39_ ( .D(top_core_KE_n3206), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__40_ ( .D(top_core_KE_n4237), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__40_ ( .D(top_core_KE_n3721), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__40_ ( .D(top_core_KE_n3205), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__41_ ( .D(top_core_KE_n4236), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__41_ ( .D(top_core_KE_n3720), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__41_ ( .D(top_core_KE_n3204), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__42_ ( .D(top_core_KE_n4235), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__42_ ( .D(top_core_KE_n3719), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__42_ ( .D(top_core_KE_n3203), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__43_ ( .D(top_core_KE_n4234), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__43_ ( .D(top_core_KE_n3718), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__43_ ( .D(top_core_KE_n3202), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__44_ ( .D(top_core_KE_n4233), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__44_ ( .D(top_core_KE_n3717), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__44_ ( .D(top_core_KE_n3201), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__45_ ( .D(top_core_KE_n4232), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__45_ ( .D(top_core_KE_n3716), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__45_ ( .D(top_core_KE_n3200), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__46_ ( .D(top_core_KE_n4231), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__46_ ( .D(top_core_KE_n3715), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__46_ ( .D(top_core_KE_n3199), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__47_ ( .D(top_core_KE_n4230), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__47_ ( .D(top_core_KE_n3714), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__47_ ( .D(top_core_KE_n3198), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__48_ ( .D(top_core_KE_n4229), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__48_ ( .D(top_core_KE_n3713), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__48_ ( .D(top_core_KE_n3197), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__49_ ( .D(top_core_KE_n4228), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__49_ ( .D(top_core_KE_n3712), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__49_ ( .D(top_core_KE_n3196), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__50_ ( .D(top_core_KE_n4227), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__50_ ( .D(top_core_KE_n3711), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__50_ ( .D(top_core_KE_n3195), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__51_ ( .D(top_core_KE_n4226), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__51_ ( .D(top_core_KE_n3710), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__51_ ( .D(top_core_KE_n3194), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__52_ ( .D(top_core_KE_n4225), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__52_ ( .D(top_core_KE_n3709), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__52_ ( .D(top_core_KE_n3193), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__53_ ( .D(top_core_KE_n4224), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__53_ ( .D(top_core_KE_n3708), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__53_ ( .D(top_core_KE_n3192), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__54_ ( .D(top_core_KE_n4223), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__54_ ( .D(top_core_KE_n3707), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__54_ ( .D(top_core_KE_n3191), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__55_ ( .D(top_core_KE_n4222), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__55_ ( .D(top_core_KE_n3706), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__55_ ( .D(top_core_KE_n3190), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__56_ ( .D(top_core_KE_n4221), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__56_ ( .D(top_core_KE_n3705), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__56_ ( .D(top_core_KE_n3189), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__57_ ( .D(top_core_KE_n4220), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__57_ ( .D(top_core_KE_n3704), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__57_ ( .D(top_core_KE_n3188), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__58_ ( .D(top_core_KE_n4219), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__58_ ( .D(top_core_KE_n3703), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__58_ ( .D(top_core_KE_n3187), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__59_ ( .D(top_core_KE_n4218), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__59_ ( .D(top_core_KE_n3702), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__59_ ( .D(top_core_KE_n3186), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__60_ ( .D(top_core_KE_n4217), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__60_ ( .D(top_core_KE_n3701), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__60_ ( .D(top_core_KE_n3185), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__61_ ( .D(top_core_KE_n4216), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__61_ ( .D(top_core_KE_n3700), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__61_ ( .D(top_core_KE_n3184), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__62_ ( .D(top_core_KE_n4215), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__62_ ( .D(top_core_KE_n3699), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__62_ ( .D(top_core_KE_n3183), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__63_ ( .D(top_core_KE_n4214), .CK(n3889), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__63_ ( .D(top_core_KE_n3698), .CK(n3889), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__63_ ( .D(top_core_KE_n3182), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__88_ ( .D(top_core_KE_n4189), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__88_ ( .D(top_core_KE_n3673), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__88_ ( .D(top_core_KE_n3157), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__89_ ( .D(top_core_KE_n4188), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__89_ ( .D(top_core_KE_n3672), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__89_ ( .D(top_core_KE_n3156), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__90_ ( .D(top_core_KE_n4187), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__90_ ( .D(top_core_KE_n3671), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__90_ ( .D(top_core_KE_n3155), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__91_ ( .D(top_core_KE_n4186), .CK(n3889), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__91_ ( .D(top_core_KE_n3670), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__91_ ( .D(top_core_KE_n3154), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__92_ ( .D(top_core_KE_n4185), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__92_ ( .D(top_core_KE_n3669), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__92_ ( .D(top_core_KE_n3153), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__93_ ( .D(top_core_KE_n4184), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__93_ ( .D(top_core_KE_n3668), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__93_ ( .D(top_core_KE_n3152), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__94_ ( .D(top_core_KE_n4183), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__94_ ( .D(top_core_KE_n3667), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__94_ ( .D(top_core_KE_n3151), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__95_ ( .D(top_core_KE_n4182), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__95_ ( .D(top_core_KE_n3666), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__95_ ( .D(top_core_KE_n3150), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__96_ ( .D(top_core_KE_n4181), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__96_ ( .D(top_core_KE_n3665), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__96_ ( .D(top_core_KE_n3149), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__97_ ( .D(top_core_KE_n4180), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__97_ ( .D(top_core_KE_n3664), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__97_ ( .D(top_core_KE_n3148), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__98_ ( .D(top_core_KE_n4179), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__98_ ( .D(top_core_KE_n3663), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__98_ ( .D(top_core_KE_n3147), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__99_ ( .D(top_core_KE_n4178), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__99_ ( .D(top_core_KE_n3662), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__99_ ( .D(top_core_KE_n3146), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__100_ ( .D(top_core_KE_n4177), .CK(n3878), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__100_ ( .D(top_core_KE_n3661), .CK(n3878), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__100_ ( .D(top_core_KE_n3145), .CK(n3878), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__101_ ( .D(top_core_KE_n4176), .CK(n3879), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__101_ ( .D(top_core_KE_n3660), .CK(n3879), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__101_ ( .D(top_core_KE_n3144), .CK(n3879), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__102_ ( .D(top_core_KE_n4175), .CK(n3879), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__102_ ( .D(top_core_KE_n3659), .CK(n3880), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__102_ ( .D(top_core_KE_n3143), .CK(n3880), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__103_ ( .D(top_core_KE_n4174), .CK(n3880), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__103_ ( .D(top_core_KE_n3658), .CK(n3880), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__103_ ( .D(top_core_KE_n3142), .CK(n3881), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__104_ ( .D(top_core_KE_n4173), .CK(n3881), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__104_ ( .D(top_core_KE_n3657), .CK(n3881), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__104_ ( .D(top_core_KE_n3141), .CK(n3882), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__105_ ( .D(top_core_KE_n4172), .CK(n3882), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__105_ ( .D(top_core_KE_n3656), .CK(n3882), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__105_ ( .D(top_core_KE_n3140), .CK(n3882), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__106_ ( .D(top_core_KE_n4171), .CK(n3883), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__106_ ( .D(top_core_KE_n3655), .CK(n3822), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__106_ ( .D(top_core_KE_n3139), .CK(n3817), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__107_ ( .D(top_core_KE_n4170), .CK(n3817), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__107_ ( .D(top_core_KE_n3654), .CK(n3817), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__107_ ( .D(top_core_KE_n3138), .CK(n3818), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__108_ ( .D(top_core_KE_n4169), .CK(n3818), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__108_ ( .D(top_core_KE_n3653), .CK(n3818), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__108_ ( .D(top_core_KE_n3137), .CK(n3819), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__109_ ( .D(top_core_KE_n4168), .CK(n3819), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__109_ ( .D(top_core_KE_n3652), .CK(n3819), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__109_ ( .D(top_core_KE_n3136), .CK(n3819), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__110_ ( .D(top_core_KE_n4167), .CK(n3820), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__110_ ( .D(top_core_KE_n3651), .CK(n3820), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__110_ ( .D(top_core_KE_n3135), .CK(n3820), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__111_ ( .D(top_core_KE_n4166), .CK(n3821), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__111_ ( .D(top_core_KE_n3650), .CK(n3821), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__111_ ( .D(top_core_KE_n3134), .CK(n3821), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__120_ ( .D(top_core_KE_n4157), .CK(n3822), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__120_ ( .D(top_core_KE_n3641), .CK(n3822), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__120_ ( .D(top_core_KE_n3125), .CK(n3822), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__121_ ( .D(top_core_KE_n4156), .CK(n3823), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__121_ ( .D(top_core_KE_n3640), .CK(n3823), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__121_ ( .D(top_core_KE_n3124), .CK(n3823), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__122_ ( .D(top_core_KE_n4155), .CK(n3823), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__122_ ( .D(top_core_KE_n3639), .CK(n3824), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__122_ ( .D(top_core_KE_n3123), .CK(n3824), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__123_ ( .D(top_core_KE_n4154), .CK(n3824), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__123_ ( .D(top_core_KE_n3638), .CK(n3824), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__123_ ( .D(top_core_KE_n3122), .CK(n3825), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__124_ ( .D(top_core_KE_n4153), .CK(n3825), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__124_ ( .D(top_core_KE_n3637), .CK(n3825), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__124_ ( .D(top_core_KE_n3121), .CK(n3826), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__125_ ( .D(top_core_KE_n4152), .CK(n3826), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__125_ ( .D(top_core_KE_n3636), .CK(n3826), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__125_ ( .D(top_core_KE_n3120), .CK(n3826), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__126_ ( .D(top_core_KE_n4151), .CK(n3811), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__126_ ( .D(top_core_KE_n3635), .CK(n3806), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__126_ ( .D(top_core_KE_n3119), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__71_ ( .D(top_core_KE_n4206), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__71_ ( .D(top_core_KE_n3690), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__71_ ( .D(top_core_KE_n3174), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__79_ ( .D(top_core_KE_n4198), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__79_ ( .D(top_core_KE_n3682), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__79_ ( .D(top_core_KE_n3166), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__119_ ( .D(top_core_KE_n4158), .CK(n3809), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__119_ ( .D(top_core_KE_n3642), .CK(n3809), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__119_ ( .D(top_core_KE_n3126), .CK(n3809), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__87_ ( .D(top_core_KE_n4190), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__87_ ( .D(top_core_KE_n3674), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__87_ ( .D(top_core_KE_n3158), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__127_ ( .D(top_core_KE_n4150), .CK(n3811), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__127_ ( .D(top_core_KE_n3634), .CK(n3811), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__127_ ( .D(top_core_KE_n3118), .CK(n3811), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__70_ ( .D(top_core_KE_n4207), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__70_ ( .D(top_core_KE_n3691), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__70_ ( .D(top_core_KE_n3175), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__78_ ( .D(top_core_KE_n4199), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__78_ ( .D(top_core_KE_n3683), .CK(n3813), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__78_ ( .D(top_core_KE_n3167), .CK(n3813), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__118_ ( .D(top_core_KE_n4159), .CK(n3813), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__118_ ( .D(top_core_KE_n3643), .CK(n3813), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__118_ ( .D(top_core_KE_n3127), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__86_ ( .D(top_core_KE_n4191), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__86_ ( .D(top_core_KE_n3675), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__86_ ( .D(top_core_KE_n3159), .CK(n3815), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__117_ ( .D(top_core_KE_n4160), .CK(n3815), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__117_ ( .D(top_core_KE_n3644), .CK(n3815), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__117_ ( .D(top_core_KE_n3128), .CK(n3815), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__85_ ( .D(top_core_KE_n4192), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__85_ ( .D(top_core_KE_n3676), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__85_ ( .D(top_core_KE_n3160), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__116_ ( .D(top_core_KE_n4161), .CK(n3837), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__116_ ( .D(top_core_KE_n3645), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__116_ ( .D(top_core_KE_n3129), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__84_ ( .D(top_core_KE_n4193), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__84_ ( .D(top_core_KE_n3677), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__84_ ( .D(top_core_KE_n3161), .CK(n3839), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__115_ ( .D(top_core_KE_n4162), .CK(n3839), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__115_ ( .D(top_core_KE_n3646), .CK(n3839), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__115_ ( .D(top_core_KE_n3130), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__83_ ( .D(top_core_KE_n4194), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__83_ ( .D(top_core_KE_n3678), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__83_ ( .D(top_core_KE_n3162), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__114_ ( .D(top_core_KE_n4163), .CK(n3841), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__114_ ( .D(top_core_KE_n3647), .CK(n3841), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__114_ ( .D(top_core_KE_n3131), .CK(n3841), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__82_ ( .D(top_core_KE_n4195), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__82_ ( .D(top_core_KE_n3679), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__82_ ( .D(top_core_KE_n3163), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__113_ ( .D(top_core_KE_n4164), .CK(n3843), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__113_ ( .D(top_core_KE_n3648), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__113_ ( .D(top_core_KE_n3132), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__81_ ( .D(top_core_KE_n4196), .CK(n3844), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__81_ ( .D(top_core_KE_n3680), .CK(n3844), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__81_ ( .D(top_core_KE_n3164), .CK(n3844), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__112_ ( .D(top_core_KE_n4165), .CK(n3844), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__112_ ( .D(top_core_KE_n3649), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__112_ ( .D(top_core_KE_n3133), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__80_ ( .D(top_core_KE_n4197), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__80_ ( .D(top_core_KE_n3681), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__80_ ( .D(top_core_KE_n3165), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__69_ ( .D(top_core_KE_n4208), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__69_ ( .D(top_core_KE_n3692), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__69_ ( .D(top_core_KE_n3176), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__77_ ( .D(top_core_KE_n4200), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__77_ ( .D(top_core_KE_n3684), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__77_ ( .D(top_core_KE_n3168), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__68_ ( .D(top_core_KE_n4209), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__68_ ( .D(top_core_KE_n3693), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__68_ ( .D(top_core_KE_n3177), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__76_ ( .D(top_core_KE_n4201), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__76_ ( .D(top_core_KE_n3685), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__76_ ( .D(top_core_KE_n3169), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__67_ ( .D(top_core_KE_n4210), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__67_ ( .D(top_core_KE_n3694), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__67_ ( .D(top_core_KE_n3178), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__75_ ( .D(top_core_KE_n4202), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__75_ ( .D(top_core_KE_n3686), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__75_ ( .D(top_core_KE_n3170), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__66_ ( .D(top_core_KE_n4211), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__66_ ( .D(top_core_KE_n3695), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__66_ ( .D(top_core_KE_n3179), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__74_ ( .D(top_core_KE_n4203), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__74_ ( .D(top_core_KE_n3687), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__74_ ( .D(top_core_KE_n3171), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__65_ ( .D(top_core_KE_n4212), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__65_ ( .D(top_core_KE_n3696), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__65_ ( .D(top_core_KE_n3180), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__73_ ( .D(top_core_KE_n4204), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__73_ ( .D(top_core_KE_n3688), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__73_ ( .D(top_core_KE_n3172), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__64_ ( .D(top_core_KE_n4213), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__64_ ( .D(top_core_KE_n3697), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__64_ ( .D(top_core_KE_n3181), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__72_ ( .D(top_core_KE_n4205), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_11__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__72_ ( .D(top_core_KE_n3689), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__72_ ( .D(top_core_KE_n3173), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_11__128_ ( .D(top_core_KE_n4149), .CK(n3837), .RN(n_RSTB), .Q(top_core_KE_key_mem_11__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_7__128_ ( .D(top_core_KE_n3633), .CK(n3837), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_7__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_3__128_ ( .D(top_core_KE_n3117), .CK(n3837), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_3__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__0_ ( .D(top_core_KE_n3890), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__1_ ( .D(top_core_KE_n3889), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__2_ ( .D(top_core_KE_n3888), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__3_ ( .D(top_core_KE_n3887), .CK(n3730), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__4_ ( .D(top_core_KE_n3886), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__5_ ( .D(top_core_KE_n3885), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__6_ ( .D(top_core_KE_n3884), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__7_ ( .D(top_core_KE_n3883), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__8_ ( .D(top_core_KE_n3882), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__9_ ( .D(top_core_KE_n3881), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__10_ ( .D(top_core_KE_n3880), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__11_ ( .D(top_core_KE_n3879), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__12_ ( .D(top_core_KE_n3878), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__13_ ( .D(top_core_KE_n3877), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__14_ ( .D(top_core_KE_n3876), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__15_ ( .D(top_core_KE_n3875), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__16_ ( .D(top_core_KE_n3874), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__17_ ( .D(top_core_KE_n3873), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__18_ ( .D(top_core_KE_n3872), .CK(n3731), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__19_ ( .D(top_core_KE_n3871), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__20_ ( .D(top_core_KE_n3870), .CK(n3955), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__21_ ( .D(top_core_KE_n3869), .CK(n3956), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__22_ ( .D(top_core_KE_n3868), .CK(n3953), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__23_ ( .D(top_core_KE_n3867), .CK(n3949), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__24_ ( .D(top_core_KE_n3866), .CK(n3948), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__25_ ( .D(top_core_KE_n3865), .CK(n3952), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__26_ ( .D(top_core_KE_n3864), .CK(
        top_core_clk_slow), .RN(n_RSTB), .Q(top_core_KE_key_mem_8__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__27_ ( .D(top_core_KE_n3863), .CK(n3906), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__28_ ( .D(top_core_KE_n3862), .CK(n3960), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__29_ ( .D(top_core_KE_n3861), .CK(n3722), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__30_ ( .D(top_core_KE_n3860), .CK(n3951), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__31_ ( .D(top_core_KE_n3859), .CK(n3906), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__32_ ( .D(top_core_KE_n3858), .CK(n3906), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__33_ ( .D(top_core_KE_n3857), .CK(n3950), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__34_ ( .D(top_core_KE_n3856), .CK(n3954), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__35_ ( .D(top_core_KE_n3855), .CK(n3959), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__36_ ( .D(top_core_KE_n3854), .CK(n3958), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__37_ ( .D(top_core_KE_n3853), .CK(n3952), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__38_ ( .D(top_core_KE_n3852), .CK(n3957), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__39_ ( .D(top_core_KE_n3851), .CK(n3952), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__40_ ( .D(top_core_KE_n3850), .CK(n3951), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__41_ ( .D(top_core_KE_n3849), .CK(n3950), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__42_ ( .D(top_core_KE_n3848), .CK(n3954), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__43_ ( .D(top_core_KE_n3847), .CK(n3959), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__44_ ( .D(top_core_KE_n3846), .CK(n3958), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__45_ ( .D(top_core_KE_n3845), .CK(n3960), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__46_ ( .D(top_core_KE_n3844), .CK(n3957), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__47_ ( .D(top_core_KE_n3843), .CK(n3952), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__48_ ( .D(top_core_KE_n3842), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__49_ ( .D(top_core_KE_n3841), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__50_ ( .D(top_core_KE_n3840), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__51_ ( .D(top_core_KE_n3839), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__52_ ( .D(top_core_KE_n3838), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__53_ ( .D(top_core_KE_n3837), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__54_ ( .D(top_core_KE_n3836), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__55_ ( .D(top_core_KE_n3835), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__56_ ( .D(top_core_KE_n3834), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__57_ ( .D(top_core_KE_n3833), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__58_ ( .D(top_core_KE_n3832), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__59_ ( .D(top_core_KE_n3831), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__60_ ( .D(top_core_KE_n3830), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__61_ ( .D(top_core_KE_n3829), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__62_ ( .D(top_core_KE_n3828), .CK(n3709), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__63_ ( .D(top_core_KE_n3827), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__64_ ( .D(top_core_KE_n3826), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__65_ ( .D(top_core_KE_n3825), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__66_ ( .D(top_core_KE_n3824), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__67_ ( .D(top_core_KE_n3823), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__68_ ( .D(top_core_KE_n3822), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__69_ ( .D(top_core_KE_n3821), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__70_ ( .D(top_core_KE_n3820), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__71_ ( .D(top_core_KE_n3819), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__72_ ( .D(top_core_KE_n3818), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__73_ ( .D(top_core_KE_n3817), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__74_ ( .D(top_core_KE_n3816), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__75_ ( .D(top_core_KE_n3815), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__76_ ( .D(top_core_KE_n3814), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__77_ ( .D(top_core_KE_n3813), .CK(n3710), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__78_ ( .D(top_core_KE_n3812), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__79_ ( .D(top_core_KE_n3811), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__80_ ( .D(top_core_KE_n3810), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__81_ ( .D(top_core_KE_n3809), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__82_ ( .D(top_core_KE_n3808), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__83_ ( .D(top_core_KE_n3807), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__84_ ( .D(top_core_KE_n3806), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__85_ ( .D(top_core_KE_n3805), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__86_ ( .D(top_core_KE_n3804), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__87_ ( .D(top_core_KE_n3803), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__88_ ( .D(top_core_KE_n3802), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__89_ ( .D(top_core_KE_n3801), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__90_ ( .D(top_core_KE_n3800), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__91_ ( .D(top_core_KE_n3799), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__92_ ( .D(top_core_KE_n3798), .CK(n3711), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__93_ ( .D(top_core_KE_n3797), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__94_ ( .D(top_core_KE_n3796), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__95_ ( .D(top_core_KE_n3795), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__96_ ( .D(top_core_KE_n3794), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__97_ ( .D(top_core_KE_n3793), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__98_ ( .D(top_core_KE_n3792), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__99_ ( .D(top_core_KE_n3791), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__100_ ( .D(top_core_KE_n3790), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__101_ ( .D(top_core_KE_n3789), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__102_ ( .D(top_core_KE_n3788), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__103_ ( .D(top_core_KE_n3787), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__104_ ( .D(top_core_KE_n3786), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__105_ ( .D(top_core_KE_n3785), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__106_ ( .D(top_core_KE_n3784), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__107_ ( .D(top_core_KE_n3783), .CK(n3712), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__108_ ( .D(top_core_KE_n3782), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__109_ ( .D(top_core_KE_n3781), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__110_ ( .D(top_core_KE_n3780), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__111_ ( .D(top_core_KE_n3779), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__112_ ( .D(top_core_KE_n3778), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__113_ ( .D(top_core_KE_n3777), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__114_ ( .D(top_core_KE_n3776), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__115_ ( .D(top_core_KE_n3775), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__116_ ( .D(top_core_KE_n3774), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__117_ ( .D(top_core_KE_n3773), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__118_ ( .D(top_core_KE_n3772), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__119_ ( .D(top_core_KE_n3771), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__120_ ( .D(top_core_KE_n3770), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__121_ ( .D(top_core_KE_n3769), .CK(n3713), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__122_ ( .D(top_core_KE_n3768), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__123_ ( .D(top_core_KE_n3767), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__124_ ( .D(top_core_KE_n3766), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__125_ ( .D(top_core_KE_n3765), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__126_ ( .D(top_core_KE_n3764), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__127_ ( .D(top_core_KE_n3763), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_8__128_ ( .D(top_core_KE_n3762), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_8__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__0_ ( .D(top_core_KE_n3374), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__0_ ( .D(top_core_KE_n2858), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__1_ ( .D(top_core_KE_n3373), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__1_ ( .D(top_core_KE_n2857), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__2_ ( .D(top_core_KE_n3372), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__2_ ( .D(top_core_KE_n2856), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__3_ ( .D(top_core_KE_n3371), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__3_ ( .D(top_core_KE_n2855), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__4_ ( .D(top_core_KE_n3370), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__4_ ( .D(top_core_KE_n2854), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__5_ ( .D(top_core_KE_n3369), .CK(n3719), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__5_ ( .D(top_core_KE_n2853), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__6_ ( .D(top_core_KE_n3368), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__6_ ( .D(top_core_KE_n2852), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__7_ ( .D(top_core_KE_n3367), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__7_ ( .D(top_core_KE_n2851), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__8_ ( .D(top_core_KE_n3366), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__8_ ( .D(top_core_KE_n2850), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__9_ ( .D(top_core_KE_n3365), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__9_ ( .D(top_core_KE_n2849), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__10_ ( .D(top_core_KE_n3364), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__10_ ( .D(top_core_KE_n2848), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__11_ ( .D(top_core_KE_n3363), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__11_ ( .D(top_core_KE_n2847), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__12_ ( .D(top_core_KE_n3362), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__12_ ( .D(top_core_KE_n2846), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__13_ ( .D(top_core_KE_n3361), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__13_ ( .D(top_core_KE_n2845), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__14_ ( .D(top_core_KE_n3360), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__14_ ( .D(top_core_KE_n2844), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__15_ ( .D(top_core_KE_n3359), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__15_ ( .D(top_core_KE_n2843), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__16_ ( .D(top_core_KE_n3358), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__16_ ( .D(top_core_KE_n2842), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__17_ ( .D(top_core_KE_n3357), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__17_ ( .D(top_core_KE_n2841), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__18_ ( .D(top_core_KE_n3356), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__18_ ( .D(top_core_KE_n2840), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__19_ ( .D(top_core_KE_n3355), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__19_ ( .D(top_core_KE_n2839), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__20_ ( .D(top_core_KE_n3354), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__20_ ( .D(top_core_KE_n2838), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__21_ ( .D(top_core_KE_n3353), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__21_ ( .D(top_core_KE_n2837), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__22_ ( .D(top_core_KE_n3352), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__22_ ( .D(top_core_KE_n2836), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__23_ ( .D(top_core_KE_n3351), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__23_ ( .D(top_core_KE_n2835), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__24_ ( .D(top_core_KE_n3350), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__24_ ( .D(top_core_KE_n2834), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__25_ ( .D(top_core_KE_n3349), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__25_ ( .D(top_core_KE_n2833), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__26_ ( .D(top_core_KE_n3348), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__26_ ( .D(top_core_KE_n2832), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__27_ ( .D(top_core_KE_n3347), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__27_ ( .D(top_core_KE_n2831), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__28_ ( .D(top_core_KE_n3346), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__28_ ( .D(top_core_KE_n2830), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__29_ ( .D(top_core_KE_n3345), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__29_ ( .D(top_core_KE_n2829), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__30_ ( .D(top_core_KE_n3344), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__30_ ( .D(top_core_KE_n2828), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__31_ ( .D(top_core_KE_n3343), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__31_ ( .D(top_core_KE_n2827), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__32_ ( .D(top_core_KE_n3342), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__32_ ( .D(top_core_KE_n2826), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__33_ ( .D(top_core_KE_n3341), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__33_ ( .D(top_core_KE_n2825), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__34_ ( .D(top_core_KE_n3340), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__34_ ( .D(top_core_KE_n2824), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__35_ ( .D(top_core_KE_n3339), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__35_ ( .D(top_core_KE_n2823), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__36_ ( .D(top_core_KE_n3338), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__36_ ( .D(top_core_KE_n2822), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__37_ ( .D(top_core_KE_n3337), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__37_ ( .D(top_core_KE_n2821), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__38_ ( .D(top_core_KE_n3336), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__38_ ( .D(top_core_KE_n2820), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__39_ ( .D(top_core_KE_n3335), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__39_ ( .D(top_core_KE_n2819), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__40_ ( .D(top_core_KE_n3334), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__40_ ( .D(top_core_KE_n2818), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__41_ ( .D(top_core_KE_n3333), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__41_ ( .D(top_core_KE_n2817), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__42_ ( .D(top_core_KE_n3332), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__42_ ( .D(top_core_KE_n2816), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__43_ ( .D(top_core_KE_n3331), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__43_ ( .D(top_core_KE_n2815), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__44_ ( .D(top_core_KE_n3330), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__44_ ( .D(top_core_KE_n2814), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__45_ ( .D(top_core_KE_n3329), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__45_ ( .D(top_core_KE_n2813), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__46_ ( .D(top_core_KE_n3328), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__46_ ( .D(top_core_KE_n2812), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__47_ ( .D(top_core_KE_n3327), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__47_ ( .D(top_core_KE_n2811), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__48_ ( .D(top_core_KE_n3326), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__48_ ( .D(top_core_KE_n2810), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__49_ ( .D(top_core_KE_n3325), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__49_ ( .D(top_core_KE_n2809), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__50_ ( .D(top_core_KE_n3324), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__50_ ( .D(top_core_KE_n2808), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__51_ ( .D(top_core_KE_n3323), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__51_ ( .D(top_core_KE_n2807), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__52_ ( .D(top_core_KE_n3322), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__52_ ( .D(top_core_KE_n2806), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__53_ ( .D(top_core_KE_n3321), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__53_ ( .D(top_core_KE_n2805), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__54_ ( .D(top_core_KE_n3320), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__54_ ( .D(top_core_KE_n2804), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__55_ ( .D(top_core_KE_n3319), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__55_ ( .D(top_core_KE_n2803), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__56_ ( .D(top_core_KE_n3318), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__56_ ( .D(top_core_KE_n2802), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__57_ ( .D(top_core_KE_n3317), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__57_ ( .D(top_core_KE_n2801), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__58_ ( .D(top_core_KE_n3316), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__58_ ( .D(top_core_KE_n2800), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__59_ ( .D(top_core_KE_n3315), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__59_ ( .D(top_core_KE_n2799), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__60_ ( .D(top_core_KE_n3314), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__60_ ( .D(top_core_KE_n2798), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__61_ ( .D(top_core_KE_n3313), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__61_ ( .D(top_core_KE_n2797), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__62_ ( .D(top_core_KE_n3312), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__62_ ( .D(top_core_KE_n2796), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__63_ ( .D(top_core_KE_n3311), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__63_ ( .D(top_core_KE_n2795), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__88_ ( .D(top_core_KE_n3286), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__88_ ( .D(top_core_KE_n2770), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__89_ ( .D(top_core_KE_n3285), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__89_ ( .D(top_core_KE_n2769), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__90_ ( .D(top_core_KE_n3284), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__90_ ( .D(top_core_KE_n2768), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__91_ ( .D(top_core_KE_n3283), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__91_ ( .D(top_core_KE_n2767), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__92_ ( .D(top_core_KE_n3282), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__92_ ( .D(top_core_KE_n2766), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__93_ ( .D(top_core_KE_n3281), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__93_ ( .D(top_core_KE_n2765), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__94_ ( .D(top_core_KE_n3280), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__94_ ( .D(top_core_KE_n2764), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__95_ ( .D(top_core_KE_n3279), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__95_ ( .D(top_core_KE_n2763), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__96_ ( .D(top_core_KE_n3278), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__96_ ( .D(top_core_KE_n2762), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__97_ ( .D(top_core_KE_n3277), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__97_ ( .D(top_core_KE_n2761), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__98_ ( .D(top_core_KE_n3276), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__98_ ( .D(top_core_KE_n2760), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__99_ ( .D(top_core_KE_n3275), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__99_ ( .D(top_core_KE_n2759), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__100_ ( .D(top_core_KE_n3274), .CK(n3878), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__100_ ( .D(top_core_KE_n2758), .CK(n3878), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__101_ ( .D(top_core_KE_n3273), .CK(n3879), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__101_ ( .D(top_core_KE_n2757), .CK(n3879), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__102_ ( .D(top_core_KE_n3272), .CK(n3880), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__102_ ( .D(top_core_KE_n2756), .CK(n3880), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__103_ ( .D(top_core_KE_n3271), .CK(n3881), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__103_ ( .D(top_core_KE_n2755), .CK(n3881), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__104_ ( .D(top_core_KE_n3270), .CK(n3881), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__104_ ( .D(top_core_KE_n2754), .CK(n3882), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__105_ ( .D(top_core_KE_n3269), .CK(n3882), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__105_ ( .D(top_core_KE_n2753), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__106_ ( .D(top_core_KE_n3268), .CK(n3817), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__106_ ( .D(top_core_KE_n2752), .CK(n3817), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__107_ ( .D(top_core_KE_n3267), .CK(n3818), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__107_ ( .D(top_core_KE_n2751), .CK(n3818), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__108_ ( .D(top_core_KE_n3266), .CK(n3819), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__108_ ( .D(top_core_KE_n2750), .CK(n3819), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__109_ ( .D(top_core_KE_n3265), .CK(n3819), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__109_ ( .D(top_core_KE_n2749), .CK(n3820), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__110_ ( .D(top_core_KE_n3264), .CK(n3820), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__110_ ( .D(top_core_KE_n2748), .CK(n3821), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__111_ ( .D(top_core_KE_n3263), .CK(n3821), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__111_ ( .D(top_core_KE_n2747), .CK(n3821), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__120_ ( .D(top_core_KE_n3254), .CK(n3822), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__120_ ( .D(top_core_KE_n2738), .CK(n3822), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__121_ ( .D(top_core_KE_n3253), .CK(n3823), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__121_ ( .D(top_core_KE_n2737), .CK(n3823), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__122_ ( .D(top_core_KE_n3252), .CK(n3824), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__122_ ( .D(top_core_KE_n2736), .CK(n3824), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__123_ ( .D(top_core_KE_n3251), .CK(n3825), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__123_ ( .D(top_core_KE_n2735), .CK(n3825), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__124_ ( .D(top_core_KE_n3250), .CK(n3826), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__124_ ( .D(top_core_KE_n2734), .CK(n3826), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__125_ ( .D(top_core_KE_n3249), .CK(n3826), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__125_ ( .D(top_core_KE_n2733), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__126_ ( .D(top_core_KE_n3248), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__126_ ( .D(top_core_KE_n2732), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__71_ ( .D(top_core_KE_n3303), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__71_ ( .D(top_core_KE_n2787), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__79_ ( .D(top_core_KE_n3295), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__79_ ( .D(top_core_KE_n2779), .CK(n3809), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__119_ ( .D(top_core_KE_n3255), .CK(n3809), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__119_ ( .D(top_core_KE_n2739), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__87_ ( .D(top_core_KE_n3287), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__87_ ( .D(top_core_KE_n2771), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__127_ ( .D(top_core_KE_n3247), .CK(n3811), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__127_ ( .D(top_core_KE_n2731), .CK(n3811), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__70_ ( .D(top_core_KE_n3304), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__70_ ( .D(top_core_KE_n2788), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__78_ ( .D(top_core_KE_n3296), .CK(n3813), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__78_ ( .D(top_core_KE_n2780), .CK(n3813), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__118_ ( .D(top_core_KE_n3256), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__118_ ( .D(top_core_KE_n2740), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__86_ ( .D(top_core_KE_n3288), .CK(n3815), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__86_ ( .D(top_core_KE_n2772), .CK(n3815), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__117_ ( .D(top_core_KE_n3257), .CK(n3815), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__117_ ( .D(top_core_KE_n2741), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__85_ ( .D(top_core_KE_n3289), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__85_ ( .D(top_core_KE_n2773), .CK(n3817), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__116_ ( .D(top_core_KE_n3258), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__116_ ( .D(top_core_KE_n2742), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__84_ ( .D(top_core_KE_n3290), .CK(n3839), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__84_ ( .D(top_core_KE_n2774), .CK(n3839), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__115_ ( .D(top_core_KE_n3259), .CK(n3839), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__115_ ( .D(top_core_KE_n2743), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__83_ ( .D(top_core_KE_n3291), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__83_ ( .D(top_core_KE_n2775), .CK(n3841), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__114_ ( .D(top_core_KE_n3260), .CK(n3841), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__114_ ( .D(top_core_KE_n2744), .CK(n3841), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__82_ ( .D(top_core_KE_n3292), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__82_ ( .D(top_core_KE_n2776), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__113_ ( .D(top_core_KE_n3261), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__113_ ( .D(top_core_KE_n2745), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__81_ ( .D(top_core_KE_n3293), .CK(n3844), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__81_ ( .D(top_core_KE_n2777), .CK(n3844), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__112_ ( .D(top_core_KE_n3262), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__112_ ( .D(top_core_KE_n2746), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__80_ ( .D(top_core_KE_n3294), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__80_ ( .D(top_core_KE_n2778), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__69_ ( .D(top_core_KE_n3305), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__69_ ( .D(top_core_KE_n2789), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__77_ ( .D(top_core_KE_n3297), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__77_ ( .D(top_core_KE_n2781), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__68_ ( .D(top_core_KE_n3306), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__68_ ( .D(top_core_KE_n2790), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__76_ ( .D(top_core_KE_n3298), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__76_ ( .D(top_core_KE_n2782), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__67_ ( .D(top_core_KE_n3307), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__67_ ( .D(top_core_KE_n2791), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__75_ ( .D(top_core_KE_n3299), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__75_ ( .D(top_core_KE_n2783), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__66_ ( .D(top_core_KE_n3308), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__66_ ( .D(top_core_KE_n2792), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__74_ ( .D(top_core_KE_n3300), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__74_ ( .D(top_core_KE_n2784), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__65_ ( .D(top_core_KE_n3309), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__65_ ( .D(top_core_KE_n2793), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__73_ ( .D(top_core_KE_n3301), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__73_ ( .D(top_core_KE_n2785), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__64_ ( .D(top_core_KE_n3310), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__64_ ( .D(top_core_KE_n2794), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__72_ ( .D(top_core_KE_n3302), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__72_ ( .D(top_core_KE_n2786), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_4__128_ ( .D(top_core_KE_n3246), .CK(n3837), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_4__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_0__128_ ( .D(top_core_KE_n2730), .CK(n3837), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_0__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__0_ ( .D(top_core_KE_n4148), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__0_ ( .D(top_core_KE_n3632), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__0_ ( .D(top_core_KE_n3116), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__1_ ( .D(top_core_KE_n4147), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__1_ ( .D(top_core_KE_n3631), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__1_ ( .D(top_core_KE_n3115), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__2_ ( .D(top_core_KE_n4146), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__2_ ( .D(top_core_KE_n3630), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__2_ ( .D(top_core_KE_n3114), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__3_ ( .D(top_core_KE_n4145), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__3_ ( .D(top_core_KE_n3629), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__3_ ( .D(top_core_KE_n3113), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__4_ ( .D(top_core_KE_n4144), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__4_ ( .D(top_core_KE_n3628), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__4_ ( .D(top_core_KE_n3112), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__5_ ( .D(top_core_KE_n4143), .CK(n3719), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__5_ ( .D(top_core_KE_n3627), .CK(n3719), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__5_ ( .D(top_core_KE_n3111), .CK(n3719), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__6_ ( .D(top_core_KE_n4142), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__6_ ( .D(top_core_KE_n3626), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__6_ ( .D(top_core_KE_n3110), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__7_ ( .D(top_core_KE_n4141), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__7_ ( .D(top_core_KE_n3625), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__7_ ( .D(top_core_KE_n3109), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__8_ ( .D(top_core_KE_n4140), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__8_ ( .D(top_core_KE_n3624), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__8_ ( .D(top_core_KE_n3108), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__9_ ( .D(top_core_KE_n4139), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__9_ ( .D(top_core_KE_n3623), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__9_ ( .D(top_core_KE_n3107), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__10_ ( .D(top_core_KE_n4138), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__10_ ( .D(top_core_KE_n3622), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__10_ ( .D(top_core_KE_n3106), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__11_ ( .D(top_core_KE_n4137), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__11_ ( .D(top_core_KE_n3621), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__11_ ( .D(top_core_KE_n3105), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__12_ ( .D(top_core_KE_n4136), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__12_ ( .D(top_core_KE_n3620), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__12_ ( .D(top_core_KE_n3104), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__13_ ( .D(top_core_KE_n4135), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__13_ ( .D(top_core_KE_n3619), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__13_ ( .D(top_core_KE_n3103), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__14_ ( .D(top_core_KE_n4134), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__14_ ( .D(top_core_KE_n3618), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__14_ ( .D(top_core_KE_n3102), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__15_ ( .D(top_core_KE_n4133), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__15_ ( .D(top_core_KE_n3617), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__15_ ( .D(top_core_KE_n3101), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__16_ ( .D(top_core_KE_n4132), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__16_ ( .D(top_core_KE_n3616), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__16_ ( .D(top_core_KE_n3100), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__17_ ( .D(top_core_KE_n4131), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__17_ ( .D(top_core_KE_n3615), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__17_ ( .D(top_core_KE_n3099), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__18_ ( .D(top_core_KE_n4130), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__18_ ( .D(top_core_KE_n3614), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__18_ ( .D(top_core_KE_n3098), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__19_ ( .D(top_core_KE_n4129), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__19_ ( .D(top_core_KE_n3613), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__19_ ( .D(top_core_KE_n3097), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__20_ ( .D(top_core_KE_n4128), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__20_ ( .D(top_core_KE_n3612), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__20_ ( .D(top_core_KE_n3096), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__21_ ( .D(top_core_KE_n4127), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__21_ ( .D(top_core_KE_n3611), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__21_ ( .D(top_core_KE_n3095), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__22_ ( .D(top_core_KE_n4126), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__22_ ( .D(top_core_KE_n3610), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__22_ ( .D(top_core_KE_n3094), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__23_ ( .D(top_core_KE_n4125), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__23_ ( .D(top_core_KE_n3609), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__23_ ( .D(top_core_KE_n3093), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__24_ ( .D(top_core_KE_n4124), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__24_ ( .D(top_core_KE_n3608), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__24_ ( .D(top_core_KE_n3092), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__25_ ( .D(top_core_KE_n4123), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__25_ ( .D(top_core_KE_n3607), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__25_ ( .D(top_core_KE_n3091), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__26_ ( .D(top_core_KE_n4122), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__26_ ( .D(top_core_KE_n3606), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__26_ ( .D(top_core_KE_n3090), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__27_ ( .D(top_core_KE_n4121), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__27_ ( .D(top_core_KE_n3605), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__27_ ( .D(top_core_KE_n3089), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__28_ ( .D(top_core_KE_n4120), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__28_ ( .D(top_core_KE_n3604), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__28_ ( .D(top_core_KE_n3088), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__29_ ( .D(top_core_KE_n4119), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__29_ ( .D(top_core_KE_n3603), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__29_ ( .D(top_core_KE_n3087), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__30_ ( .D(top_core_KE_n4118), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__30_ ( .D(top_core_KE_n3602), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__30_ ( .D(top_core_KE_n3086), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__31_ ( .D(top_core_KE_n4117), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__31_ ( .D(top_core_KE_n3601), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__31_ ( .D(top_core_KE_n3085), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__32_ ( .D(top_core_KE_n4116), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__32_ ( .D(top_core_KE_n3600), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__32_ ( .D(top_core_KE_n3084), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__33_ ( .D(top_core_KE_n4115), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__33_ ( .D(top_core_KE_n3599), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__33_ ( .D(top_core_KE_n3083), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__34_ ( .D(top_core_KE_n4114), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__34_ ( .D(top_core_KE_n3598), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__34_ ( .D(top_core_KE_n3082), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__35_ ( .D(top_core_KE_n4113), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__35_ ( .D(top_core_KE_n3597), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__35_ ( .D(top_core_KE_n3081), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__36_ ( .D(top_core_KE_n4112), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__36_ ( .D(top_core_KE_n3596), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__36_ ( .D(top_core_KE_n3080), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__37_ ( .D(top_core_KE_n4111), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__37_ ( .D(top_core_KE_n3595), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__37_ ( .D(top_core_KE_n3079), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__38_ ( .D(top_core_KE_n4110), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__38_ ( .D(top_core_KE_n3594), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__38_ ( .D(top_core_KE_n3078), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__39_ ( .D(top_core_KE_n4109), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__39_ ( .D(top_core_KE_n3593), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__39_ ( .D(top_core_KE_n3077), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__40_ ( .D(top_core_KE_n4108), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__40_ ( .D(top_core_KE_n3592), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__40_ ( .D(top_core_KE_n3076), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__41_ ( .D(top_core_KE_n4107), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__41_ ( .D(top_core_KE_n3591), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__41_ ( .D(top_core_KE_n3075), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__42_ ( .D(top_core_KE_n4106), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__42_ ( .D(top_core_KE_n3590), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__42_ ( .D(top_core_KE_n3074), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__43_ ( .D(top_core_KE_n4105), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__43_ ( .D(top_core_KE_n3589), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__43_ ( .D(top_core_KE_n3073), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__44_ ( .D(top_core_KE_n4104), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__44_ ( .D(top_core_KE_n3588), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__44_ ( .D(top_core_KE_n3072), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__45_ ( .D(top_core_KE_n4103), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__45_ ( .D(top_core_KE_n3587), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__45_ ( .D(top_core_KE_n3071), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__46_ ( .D(top_core_KE_n4102), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__46_ ( .D(top_core_KE_n3586), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__46_ ( .D(top_core_KE_n3070), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__47_ ( .D(top_core_KE_n4101), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__47_ ( .D(top_core_KE_n3585), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__47_ ( .D(top_core_KE_n3069), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__48_ ( .D(top_core_KE_n4100), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__48_ ( .D(top_core_KE_n3584), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__48_ ( .D(top_core_KE_n3068), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__49_ ( .D(top_core_KE_n4099), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__49_ ( .D(top_core_KE_n3583), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__49_ ( .D(top_core_KE_n3067), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__50_ ( .D(top_core_KE_n4098), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__50_ ( .D(top_core_KE_n3582), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__50_ ( .D(top_core_KE_n3066), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__51_ ( .D(top_core_KE_n4097), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__51_ ( .D(top_core_KE_n3581), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__51_ ( .D(top_core_KE_n3065), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__52_ ( .D(top_core_KE_n4096), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__52_ ( .D(top_core_KE_n3580), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__52_ ( .D(top_core_KE_n3064), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__53_ ( .D(top_core_KE_n4095), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__53_ ( .D(top_core_KE_n3579), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__53_ ( .D(top_core_KE_n3063), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__54_ ( .D(top_core_KE_n4094), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__54_ ( .D(top_core_KE_n3578), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__54_ ( .D(top_core_KE_n3062), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__55_ ( .D(top_core_KE_n4093), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__55_ ( .D(top_core_KE_n3577), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__55_ ( .D(top_core_KE_n3061), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__56_ ( .D(top_core_KE_n4092), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__56_ ( .D(top_core_KE_n3576), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__56_ ( .D(top_core_KE_n3060), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__57_ ( .D(top_core_KE_n4091), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__57_ ( .D(top_core_KE_n3575), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__57_ ( .D(top_core_KE_n3059), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__58_ ( .D(top_core_KE_n4090), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__58_ ( .D(top_core_KE_n3574), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__58_ ( .D(top_core_KE_n3058), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__59_ ( .D(top_core_KE_n4089), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__59_ ( .D(top_core_KE_n3573), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__59_ ( .D(top_core_KE_n3057), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__60_ ( .D(top_core_KE_n4088), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__60_ ( .D(top_core_KE_n3572), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__60_ ( .D(top_core_KE_n3056), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__61_ ( .D(top_core_KE_n4087), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__61_ ( .D(top_core_KE_n3571), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__61_ ( .D(top_core_KE_n3055), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__62_ ( .D(top_core_KE_n4086), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__62_ ( .D(top_core_KE_n3570), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__62_ ( .D(top_core_KE_n3054), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__63_ ( .D(top_core_KE_n4085), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__63_ ( .D(top_core_KE_n3569), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__63_ ( .D(top_core_KE_n3053), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__88_ ( .D(top_core_KE_n4060), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__88_ ( .D(top_core_KE_n3544), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__88_ ( .D(top_core_KE_n3028), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__89_ ( .D(top_core_KE_n4059), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__89_ ( .D(top_core_KE_n3543), .CK(n3885), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__89_ ( .D(top_core_KE_n3027), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__90_ ( .D(top_core_KE_n4058), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__90_ ( .D(top_core_KE_n3542), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__90_ ( .D(top_core_KE_n3026), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__91_ ( .D(top_core_KE_n4057), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__91_ ( .D(top_core_KE_n3541), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__91_ ( .D(top_core_KE_n3025), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__92_ ( .D(top_core_KE_n4056), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__92_ ( .D(top_core_KE_n3540), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__92_ ( .D(top_core_KE_n3024), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__93_ ( .D(top_core_KE_n4055), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__93_ ( .D(top_core_KE_n3539), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__93_ ( .D(top_core_KE_n3023), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__94_ ( .D(top_core_KE_n4054), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__94_ ( .D(top_core_KE_n3538), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__94_ ( .D(top_core_KE_n3022), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__95_ ( .D(top_core_KE_n4053), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__95_ ( .D(top_core_KE_n3537), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__95_ ( .D(top_core_KE_n3021), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__96_ ( .D(top_core_KE_n4052), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__96_ ( .D(top_core_KE_n3536), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__96_ ( .D(top_core_KE_n3020), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__97_ ( .D(top_core_KE_n4051), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__97_ ( .D(top_core_KE_n3535), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__97_ ( .D(top_core_KE_n3019), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__98_ ( .D(top_core_KE_n4050), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__98_ ( .D(top_core_KE_n3534), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__98_ ( .D(top_core_KE_n3018), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__99_ ( .D(top_core_KE_n4049), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__99_ ( .D(top_core_KE_n3533), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__99_ ( .D(top_core_KE_n3017), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__100_ ( .D(top_core_KE_n4048), .CK(n3878), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__100_ ( .D(top_core_KE_n3532), .CK(n3878), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__100_ ( .D(top_core_KE_n3016), .CK(n3878), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__101_ ( .D(top_core_KE_n4047), .CK(n3879), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__101_ ( .D(top_core_KE_n3531), .CK(n3879), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__101_ ( .D(top_core_KE_n3015), .CK(n3879), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__102_ ( .D(top_core_KE_n4046), .CK(n3879), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__102_ ( .D(top_core_KE_n3530), .CK(n3880), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__102_ ( .D(top_core_KE_n3014), .CK(n3880), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__103_ ( .D(top_core_KE_n4045), .CK(n3880), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__103_ ( .D(top_core_KE_n3529), .CK(n3880), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__103_ ( .D(top_core_KE_n3013), .CK(n3881), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__104_ ( .D(top_core_KE_n4044), .CK(n3881), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__104_ ( .D(top_core_KE_n3528), .CK(n3881), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__104_ ( .D(top_core_KE_n3012), .CK(n3882), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__105_ ( .D(top_core_KE_n4043), .CK(n3882), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__105_ ( .D(top_core_KE_n3527), .CK(n3882), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__105_ ( .D(top_core_KE_n3011), .CK(n3882), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__106_ ( .D(top_core_KE_n4042), .CK(n3827), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__106_ ( .D(top_core_KE_n3526), .CK(n3817), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__106_ ( .D(top_core_KE_n3010), .CK(n3817), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__107_ ( .D(top_core_KE_n4041), .CK(n3817), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__107_ ( .D(top_core_KE_n3525), .CK(n3818), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__107_ ( .D(top_core_KE_n3009), .CK(n3818), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__108_ ( .D(top_core_KE_n4040), .CK(n3818), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__108_ ( .D(top_core_KE_n3524), .CK(n3818), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__108_ ( .D(top_core_KE_n3008), .CK(n3819), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__109_ ( .D(top_core_KE_n4039), .CK(n3819), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__109_ ( .D(top_core_KE_n3523), .CK(n3819), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__109_ ( .D(top_core_KE_n3007), .CK(n3820), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__110_ ( .D(top_core_KE_n4038), .CK(n3820), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__110_ ( .D(top_core_KE_n3522), .CK(n3820), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__110_ ( .D(top_core_KE_n3006), .CK(n3820), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__111_ ( .D(top_core_KE_n4037), .CK(n3821), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__111_ ( .D(top_core_KE_n3521), .CK(n3821), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__111_ ( .D(top_core_KE_n3005), .CK(n3821), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__120_ ( .D(top_core_KE_n4028), .CK(n3822), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__120_ ( .D(top_core_KE_n3512), .CK(n3822), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__120_ ( .D(top_core_KE_n2996), .CK(n3822), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__121_ ( .D(top_core_KE_n4027), .CK(n3823), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__121_ ( .D(top_core_KE_n3511), .CK(n3823), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__121_ ( .D(top_core_KE_n2995), .CK(n3823), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__122_ ( .D(top_core_KE_n4026), .CK(n3824), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__122_ ( .D(top_core_KE_n3510), .CK(n3824), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__122_ ( .D(top_core_KE_n2994), .CK(n3824), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__123_ ( .D(top_core_KE_n4025), .CK(n3824), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__123_ ( .D(top_core_KE_n3509), .CK(n3825), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__123_ ( .D(top_core_KE_n2993), .CK(n3825), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__124_ ( .D(top_core_KE_n4024), .CK(n3825), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__124_ ( .D(top_core_KE_n3508), .CK(n3825), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__124_ ( .D(top_core_KE_n2992), .CK(n3826), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__125_ ( .D(top_core_KE_n4023), .CK(n3826), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__125_ ( .D(top_core_KE_n3507), .CK(n3826), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__125_ ( .D(top_core_KE_n2991), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__126_ ( .D(top_core_KE_n4022), .CK(n3806), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__126_ ( .D(top_core_KE_n3506), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__126_ ( .D(top_core_KE_n2990), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__71_ ( .D(top_core_KE_n4077), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__71_ ( .D(top_core_KE_n3561), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__71_ ( .D(top_core_KE_n3045), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__79_ ( .D(top_core_KE_n4069), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__79_ ( .D(top_core_KE_n3553), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__79_ ( .D(top_core_KE_n3037), .CK(n3809), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__119_ ( .D(top_core_KE_n4029), .CK(n3809), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__119_ ( .D(top_core_KE_n3513), .CK(n3809), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__119_ ( .D(top_core_KE_n2997), .CK(n3809), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__87_ ( .D(top_core_KE_n4061), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__87_ ( .D(top_core_KE_n3545), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__87_ ( .D(top_core_KE_n3029), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__127_ ( .D(top_core_KE_n4021), .CK(n3811), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__127_ ( .D(top_core_KE_n3505), .CK(n3811), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__127_ ( .D(top_core_KE_n2989), .CK(n3811), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__70_ ( .D(top_core_KE_n4078), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__70_ ( .D(top_core_KE_n3562), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__70_ ( .D(top_core_KE_n3046), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__78_ ( .D(top_core_KE_n4070), .CK(n3813), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__78_ ( .D(top_core_KE_n3554), .CK(n3813), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__78_ ( .D(top_core_KE_n3038), .CK(n3813), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__118_ ( .D(top_core_KE_n4030), .CK(n3813), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__118_ ( .D(top_core_KE_n3514), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__118_ ( .D(top_core_KE_n2998), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__86_ ( .D(top_core_KE_n4062), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__86_ ( .D(top_core_KE_n3546), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__86_ ( .D(top_core_KE_n3030), .CK(n3815), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__117_ ( .D(top_core_KE_n4031), .CK(n3815), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__117_ ( .D(top_core_KE_n3515), .CK(n3815), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__117_ ( .D(top_core_KE_n2999), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__85_ ( .D(top_core_KE_n4063), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__85_ ( .D(top_core_KE_n3547), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__85_ ( .D(top_core_KE_n3031), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__116_ ( .D(top_core_KE_n4032), .CK(n3837), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__116_ ( .D(top_core_KE_n3516), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__116_ ( .D(top_core_KE_n3000), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__84_ ( .D(top_core_KE_n4064), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__84_ ( .D(top_core_KE_n3548), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__84_ ( .D(top_core_KE_n3032), .CK(n3839), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__115_ ( .D(top_core_KE_n4033), .CK(n3839), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__115_ ( .D(top_core_KE_n3517), .CK(n3839), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__115_ ( .D(top_core_KE_n3001), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__83_ ( .D(top_core_KE_n4065), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__83_ ( .D(top_core_KE_n3549), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__83_ ( .D(top_core_KE_n3033), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__114_ ( .D(top_core_KE_n4034), .CK(n3841), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__114_ ( .D(top_core_KE_n3518), .CK(n3841), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__114_ ( .D(top_core_KE_n3002), .CK(n3841), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__82_ ( .D(top_core_KE_n4066), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__82_ ( .D(top_core_KE_n3550), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__82_ ( .D(top_core_KE_n3034), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__113_ ( .D(top_core_KE_n4035), .CK(n3843), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__113_ ( .D(top_core_KE_n3519), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__113_ ( .D(top_core_KE_n3003), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__81_ ( .D(top_core_KE_n4067), .CK(n3844), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__81_ ( .D(top_core_KE_n3551), .CK(n3844), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__81_ ( .D(top_core_KE_n3035), .CK(n3844), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__112_ ( .D(top_core_KE_n4036), .CK(n3844), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__112_ ( .D(top_core_KE_n3520), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__112_ ( .D(top_core_KE_n3004), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__80_ ( .D(top_core_KE_n4068), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__80_ ( .D(top_core_KE_n3552), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__80_ ( .D(top_core_KE_n3036), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__69_ ( .D(top_core_KE_n4079), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__69_ ( .D(top_core_KE_n3563), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__69_ ( .D(top_core_KE_n3047), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__77_ ( .D(top_core_KE_n4071), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__77_ ( .D(top_core_KE_n3555), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__77_ ( .D(top_core_KE_n3039), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__68_ ( .D(top_core_KE_n4080), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__68_ ( .D(top_core_KE_n3564), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__68_ ( .D(top_core_KE_n3048), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__76_ ( .D(top_core_KE_n4072), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__76_ ( .D(top_core_KE_n3556), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__76_ ( .D(top_core_KE_n3040), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__67_ ( .D(top_core_KE_n4081), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__67_ ( .D(top_core_KE_n3565), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__67_ ( .D(top_core_KE_n3049), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__75_ ( .D(top_core_KE_n4073), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__75_ ( .D(top_core_KE_n3557), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__75_ ( .D(top_core_KE_n3041), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__66_ ( .D(top_core_KE_n4082), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__66_ ( .D(top_core_KE_n3566), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__66_ ( .D(top_core_KE_n3050), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__74_ ( .D(top_core_KE_n4074), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__74_ ( .D(top_core_KE_n3558), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__74_ ( .D(top_core_KE_n3042), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__65_ ( .D(top_core_KE_n4083), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__65_ ( .D(top_core_KE_n3567), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__65_ ( .D(top_core_KE_n3051), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__73_ ( .D(top_core_KE_n4075), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__73_ ( .D(top_core_KE_n3559), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__73_ ( .D(top_core_KE_n3043), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__64_ ( .D(top_core_KE_n4084), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__64_ ( .D(top_core_KE_n3568), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__64_ ( .D(top_core_KE_n3052), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__72_ ( .D(top_core_KE_n4076), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_10__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__72_ ( .D(top_core_KE_n3560), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__72_ ( .D(top_core_KE_n3044), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_10__128_ ( .D(top_core_KE_n4020), .CK(n3837), .RN(n_RSTB), .Q(top_core_KE_key_mem_10__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_6__128_ ( .D(top_core_KE_n3504), .CK(n3837), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_6__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_2__128_ ( .D(top_core_KE_n2988), .CK(n3837), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_2__128_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__0_ ( .D(top_core_KE_n4406), .CK(n3714), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__0_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__1_ ( .D(top_core_KE_n4405), .CK(n3715), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__1_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__2_ ( .D(top_core_KE_n4404), .CK(n3716), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__2_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__3_ ( .D(top_core_KE_n4403), .CK(n3717), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__3_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__4_ ( .D(top_core_KE_n4402), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__4_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__5_ ( .D(top_core_KE_n4401), .CK(n3718), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__5_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__6_ ( .D(top_core_KE_n4400), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__6_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__7_ ( .D(top_core_KE_n4399), .CK(n3745), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__7_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__8_ ( .D(top_core_KE_n4398), .CK(n3746), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__8_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__9_ ( .D(top_core_KE_n4397), .CK(n3747), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__9_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__10_ ( .D(top_core_KE_n4396), .CK(n3748), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__10_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__11_ ( .D(top_core_KE_n4395), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__11_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__12_ ( .D(top_core_KE_n4394), .CK(n3749), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__12_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__13_ ( .D(top_core_KE_n4393), .CK(n3750), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__13_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__14_ ( .D(top_core_KE_n4392), .CK(n3751), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__14_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__15_ ( .D(top_core_KE_n4391), .CK(n3752), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__15_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__16_ ( .D(top_core_KE_n4390), .CK(n3753), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__16_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__17_ ( .D(top_core_KE_n4389), .CK(n3754), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__17_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__18_ ( .D(top_core_KE_n4388), .CK(n3755), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__18_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__19_ ( .D(top_core_KE_n4387), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__19_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__20_ ( .D(top_core_KE_n4386), .CK(n3756), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__20_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__21_ ( .D(top_core_KE_n4385), .CK(n3732), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__21_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__22_ ( .D(top_core_KE_n4384), .CK(n3733), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__22_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__23_ ( .D(top_core_KE_n4383), .CK(n3734), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__23_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__24_ ( .D(top_core_KE_n4382), .CK(n3735), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__24_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__25_ ( .D(top_core_KE_n4381), .CK(n3736), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__25_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__26_ ( .D(top_core_KE_n4380), .CK(n3737), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__26_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__27_ ( .D(top_core_KE_n4379), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__27_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__28_ ( .D(top_core_KE_n4378), .CK(n3738), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__28_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__29_ ( .D(top_core_KE_n4377), .CK(n3739), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__29_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__30_ ( .D(top_core_KE_n4376), .CK(n3740), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__30_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__31_ ( .D(top_core_KE_n4375), .CK(n3741), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__31_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__32_ ( .D(top_core_KE_n4374), .CK(n3742), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__32_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__33_ ( .D(top_core_KE_n4373), .CK(n3743), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__33_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__34_ ( .D(top_core_KE_n4372), .CK(n3744), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__34_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__35_ ( .D(top_core_KE_n4371), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__35_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__36_ ( .D(top_core_KE_n4370), .CK(n3860), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__36_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__37_ ( .D(top_core_KE_n4369), .CK(n3861), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__37_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__38_ ( .D(top_core_KE_n4368), .CK(n3862), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__38_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__39_ ( .D(top_core_KE_n4367), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__39_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__40_ ( .D(top_core_KE_n4366), .CK(n3863), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__40_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__41_ ( .D(top_core_KE_n4365), .CK(n3864), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__41_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__42_ ( .D(top_core_KE_n4364), .CK(n3865), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__42_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__43_ ( .D(top_core_KE_n4363), .CK(n3866), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__43_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__44_ ( .D(top_core_KE_n4362), .CK(n3867), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__44_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__45_ ( .D(top_core_KE_n4361), .CK(n3868), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__45_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__46_ ( .D(top_core_KE_n4360), .CK(n3869), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__46_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__47_ ( .D(top_core_KE_n4359), .CK(n3870), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__47_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__48_ ( .D(top_core_KE_n4358), .CK(n3848), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__48_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__49_ ( .D(top_core_KE_n4357), .CK(n3849), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__49_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__50_ ( .D(top_core_KE_n4356), .CK(n3850), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__50_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__51_ ( .D(top_core_KE_n4355), .CK(n3851), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__51_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__52_ ( .D(top_core_KE_n4354), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__52_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__53_ ( .D(top_core_KE_n4353), .CK(n3852), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__53_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__54_ ( .D(top_core_KE_n4352), .CK(n3853), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__54_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__55_ ( .D(top_core_KE_n4351), .CK(n3854), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__55_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__56_ ( .D(top_core_KE_n4350), .CK(n3855), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__56_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__57_ ( .D(top_core_KE_n4349), .CK(n3856), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__57_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__58_ ( .D(top_core_KE_n4348), .CK(n3857), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__58_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__59_ ( .D(top_core_KE_n4347), .CK(n3858), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__59_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__60_ ( .D(top_core_KE_n4346), .CK(n3859), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__60_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__61_ ( .D(top_core_KE_n4345), .CK(n3887), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__61_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__62_ ( .D(top_core_KE_n4344), .CK(n3883), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__62_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__63_ ( .D(top_core_KE_n4343), .CK(n3889), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__63_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__88_ ( .D(top_core_KE_n4318), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__88_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__89_ ( .D(top_core_KE_n4317), .CK(n3884), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__89_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__90_ ( .D(top_core_KE_n4316), .CK(n3886), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__90_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__91_ ( .D(top_core_KE_n4315), .CK(n3888), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__91_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__92_ ( .D(top_core_KE_n4314), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__92_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__93_ ( .D(top_core_KE_n4313), .CK(n3871), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__93_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__94_ ( .D(top_core_KE_n4312), .CK(n3872), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__94_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__95_ ( .D(top_core_KE_n4311), .CK(n3873), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__95_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__96_ ( .D(top_core_KE_n4310), .CK(n3874), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__96_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__97_ ( .D(top_core_KE_n4309), .CK(n3875), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__97_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__98_ ( .D(top_core_KE_n4308), .CK(n3876), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__98_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__99_ ( .D(top_core_KE_n4307), .CK(n3877), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__99_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__100_ ( .D(top_core_KE_n4306), .CK(n3878), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__100_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__101_ ( .D(top_core_KE_n4305), .CK(n3878), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__101_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__102_ ( .D(top_core_KE_n4304), .CK(n3879), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__102_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__103_ ( .D(top_core_KE_n4303), .CK(n3880), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__103_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__104_ ( .D(top_core_KE_n4302), .CK(n3881), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__104_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__105_ ( .D(top_core_KE_n4301), .CK(n3882), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__105_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__106_ ( .D(top_core_KE_n4300), .CK(n3883), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__106_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__107_ ( .D(top_core_KE_n4299), .CK(n3817), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__107_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__108_ ( .D(top_core_KE_n4298), .CK(n3818), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__108_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__109_ ( .D(top_core_KE_n4297), .CK(n3819), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__109_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__110_ ( .D(top_core_KE_n4296), .CK(n3820), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__110_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__111_ ( .D(top_core_KE_n4295), .CK(n3821), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__111_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__120_ ( .D(top_core_KE_n4286), .CK(n3822), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__120_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__121_ ( .D(top_core_KE_n4285), .CK(n3823), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__121_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__122_ ( .D(top_core_KE_n4284), .CK(n3823), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__122_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__123_ ( .D(top_core_KE_n4283), .CK(n3824), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__123_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__124_ ( .D(top_core_KE_n4282), .CK(n3825), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__124_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__125_ ( .D(top_core_KE_n4281), .CK(n3826), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__125_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__126_ ( .D(top_core_KE_n4280), .CK(n3827), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__126_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__71_ ( .D(top_core_KE_n4335), .CK(n3807), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__71_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__79_ ( .D(top_core_KE_n4327), .CK(n3808), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__79_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__119_ ( .D(top_core_KE_n4287), .CK(n3809), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__119_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__87_ ( .D(top_core_KE_n4319), .CK(n3810), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__87_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__127_ ( .D(top_core_KE_n4279), .CK(n3811), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__127_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__70_ ( .D(top_core_KE_n4336), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__70_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__78_ ( .D(top_core_KE_n4328), .CK(n3812), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__78_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__118_ ( .D(top_core_KE_n4288), .CK(n3813), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__118_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__86_ ( .D(top_core_KE_n4320), .CK(n3814), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__86_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__117_ ( .D(top_core_KE_n4289), .CK(n3815), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__117_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__85_ ( .D(top_core_KE_n4321), .CK(n3816), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__85_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__116_ ( .D(top_core_KE_n4290), .CK(n3837), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__116_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__84_ ( .D(top_core_KE_n4322), .CK(n3838), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__84_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__115_ ( .D(top_core_KE_n4291), .CK(n3839), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__115_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__83_ ( .D(top_core_KE_n4323), .CK(n3840), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__83_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__114_ ( .D(top_core_KE_n4292), .CK(n3841), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__114_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__82_ ( .D(top_core_KE_n4324), .CK(n3842), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__82_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__113_ ( .D(top_core_KE_n4293), .CK(n3843), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__113_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__81_ ( .D(top_core_KE_n4325), .CK(n3843), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__81_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__112_ ( .D(top_core_KE_n4294), .CK(n3844), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__112_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__80_ ( .D(top_core_KE_n4326), .CK(n3845), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__80_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__69_ ( .D(top_core_KE_n4337), .CK(n3846), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__69_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__77_ ( .D(top_core_KE_n4329), .CK(n3847), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__77_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__68_ ( .D(top_core_KE_n4338), .CK(n3827), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__68_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__76_ ( .D(top_core_KE_n4330), .CK(n3828), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__76_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__67_ ( .D(top_core_KE_n4339), .CK(n3829), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__67_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__75_ ( .D(top_core_KE_n4331), .CK(n3830), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__75_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__66_ ( .D(top_core_KE_n4340), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__66_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__74_ ( .D(top_core_KE_n4332), .CK(n3831), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__74_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__65_ ( .D(top_core_KE_n4341), .CK(n3832), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__65_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__73_ ( .D(top_core_KE_n4333), .CK(n3833), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__73_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__64_ ( .D(top_core_KE_n4342), .CK(n3834), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__64_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__72_ ( .D(top_core_KE_n4334), .CK(n3835), 
        .RN(n_RSTB), .Q(top_core_KE_key_mem_12__72_) );
  DFFRHQX1 top_core_KE_key_mem_reg_12__128_ ( .D(top_core_KE_n4278), .CK(n3836), .RN(n_RSTB), .Q(top_core_KE_key_mem_12__128_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_63_ ( .D(top_core_KE_n4856), .CK(n3902), .Q(top_core_KE_prev_key1_reg_63_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_127_ ( .D(top_core_KE_n4665), .CK(
        n3902), .Q(top_core_KE_prev_key0_reg_127_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_39_ ( .D(top_core_KE_n4752), .CK(n3899), .Q(top_core_KE_prev_key0_reg_39_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_95_ ( .D(top_core_KE_n4696), .CK(n3902), .Q(top_core_KE_prev_key0_reg_95_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_38_ ( .D(top_core_KE_n4753), .CK(n3903), .Q(top_core_KE_prev_key0_reg_38_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_94_ ( .D(top_core_KE_n4697), .CK(n3896), .Q(top_core_KE_prev_key0_reg_94_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_93_ ( .D(top_core_KE_n4698), .CK(n3894), .Q(top_core_KE_prev_key0_reg_93_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_92_ ( .D(top_core_KE_n4699), .CK(n3891), .Q(top_core_KE_prev_key0_reg_92_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_91_ ( .D(top_core_KE_n4700), .CK(n3904), .Q(top_core_KE_prev_key0_reg_91_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_90_ ( .D(top_core_KE_n4701), .CK(n3900), .Q(top_core_KE_prev_key0_reg_90_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_88_ ( .D(top_core_KE_n4703), .CK(n3898), .Q(top_core_KE_prev_key0_reg_88_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_37_ ( .D(top_core_KE_n4754), .CK(n3899), .Q(top_core_KE_prev_key0_reg_37_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_36_ ( .D(top_core_KE_n4755), .CK(n3901), .Q(top_core_KE_prev_key0_reg_36_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_35_ ( .D(top_core_KE_n4756), .CK(n3903), .Q(top_core_KE_prev_key0_reg_35_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_41_ ( .D(top_core_KE_n4750), .CK(n3892), .Q(top_core_KE_prev_key0_reg_41_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_40_ ( .D(top_core_KE_n4751), .CK(n3894), .Q(top_core_KE_prev_key0_reg_40_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_89_ ( .D(top_core_KE_n4702), .CK(n3896), .Q(top_core_KE_prev_key0_reg_89_) );
  DFFHQX1 top_core_KE_Nk0_reg_1_ ( .D(top_core_Nk[1]), .CK(n3687), .Q(
        top_core_KE_Nk0_1_) );
  DFFHQX1 top_core_KE_Nk0_reg_2_ ( .D(top_core_Nk[2]), .CK(n3695), .Q(
        top_core_KE_Nk0_2_) );
  DFFRHQX1 top_core_io_k_ready_reg ( .D(top_core_io_inter_ok), .CK(n3795), 
        .RN(n_RSTB), .Q(top_core_k_ready) );
  DFFRHQX1 top_core_EC_c_ready_reg ( .D(n6305), .CK(n3721), .RN(n_RSTB), .Q(
        top_core_c_ready) );
  DFFRHQX1 top_core_io_t_ready_reg ( .D(top_core_io_inter_ok), .CK(n3795), 
        .RN(n_RSTB), .Q(top_core_t_ready) );
  DFFRHQX1 top_core_EC_operation_reg ( .D(top_core_EC_n1295), .CK(n3721), .RN(
        n_RSTB), .Q(top_core_EC_operation) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_57_ ( .D(top_core_KE_n4734), .CK(n3900), .Q(top_core_KE_prev_key0_reg_57_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_47_ ( .D(top_core_KE_n4744), .CK(n3898), .Q(top_core_KE_prev_key0_reg_47_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_55_ ( .D(top_core_KE_n4736), .CK(n3897), .Q(top_core_KE_prev_key0_reg_55_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_46_ ( .D(top_core_KE_n4745), .CK(n3905), .Q(top_core_KE_prev_key0_reg_46_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_54_ ( .D(top_core_KE_n4737), .CK(n3893), .Q(top_core_KE_prev_key0_reg_54_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_62_ ( .D(top_core_KE_n4729), .CK(n3896), .Q(top_core_KE_prev_key0_reg_62_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_53_ ( .D(top_core_KE_n4738), .CK(n3896), .Q(top_core_KE_prev_key0_reg_53_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_61_ ( .D(top_core_KE_n4730), .CK(n3894), .Q(top_core_KE_prev_key0_reg_61_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_52_ ( .D(top_core_KE_n4739), .CK(n3893), .Q(top_core_KE_prev_key0_reg_52_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_60_ ( .D(top_core_KE_n4731), .CK(n3892), .Q(top_core_KE_prev_key0_reg_60_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_51_ ( .D(top_core_KE_n4740), .CK(n3905), .Q(top_core_KE_prev_key0_reg_51_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_59_ ( .D(top_core_KE_n4732), .CK(n3904), .Q(top_core_KE_prev_key0_reg_59_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_50_ ( .D(top_core_KE_n4741), .CK(n3902), .Q(top_core_KE_prev_key0_reg_50_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_58_ ( .D(top_core_KE_n4733), .CK(n3901), .Q(top_core_KE_prev_key0_reg_58_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_49_ ( .D(top_core_KE_n4742), .CK(n3897), .Q(top_core_KE_prev_key0_reg_49_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_48_ ( .D(top_core_KE_n4743), .CK(n3897), .Q(top_core_KE_prev_key0_reg_48_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_56_ ( .D(top_core_KE_n4735), .CK(n3898), .Q(top_core_KE_prev_key0_reg_56_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_45_ ( .D(top_core_KE_n4746), .CK(n3900), .Q(top_core_KE_prev_key0_reg_45_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_44_ ( .D(top_core_KE_n4747), .CK(n3902), .Q(top_core_KE_prev_key0_reg_44_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_43_ ( .D(top_core_KE_n4748), .CK(n3904), .Q(top_core_KE_prev_key0_reg_43_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_34_ ( .D(top_core_KE_n4757), .CK(n3905), .Q(top_core_KE_prev_key0_reg_34_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_42_ ( .D(top_core_KE_n4749), .CK(n3906), .Q(top_core_KE_prev_key0_reg_42_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_33_ ( .D(top_core_KE_n4758), .CK(n3891), .Q(top_core_KE_prev_key0_reg_33_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_32_ ( .D(top_core_KE_n4759), .CK(n3893), .Q(top_core_KE_prev_key0_reg_32_) );
  DFFRHQX1 top_core_io_DOUT_reg_0_ ( .D(top_core_io_N90), .CK(n_CLK), .RN(
        n_RSTB), .Q(n_DOUT[0]) );
  DFFRHQX1 top_core_io_DOUT_reg_1_ ( .D(top_core_io_N91), .CK(n_CLK), .RN(
        n_RSTB), .Q(n_DOUT[1]) );
  DFFRHQX1 top_core_io_DOUT_reg_2_ ( .D(top_core_io_N92), .CK(n_CLK), .RN(
        n_RSTB), .Q(n_DOUT[2]) );
  DFFRHQX1 top_core_io_DOUT_reg_3_ ( .D(top_core_io_N93), .CK(n_CLK), .RN(
        n_RSTB), .Q(n_DOUT[3]) );
  DFFRHQX1 top_core_io_DOUT_reg_4_ ( .D(top_core_io_N94), .CK(n_CLK), .RN(
        n_RSTB), .Q(n_DOUT[4]) );
  DFFRHQX1 top_core_io_DOUT_reg_5_ ( .D(top_core_io_N95), .CK(n_CLK), .RN(
        n_RSTB), .Q(n_DOUT[5]) );
  DFFRHQX1 top_core_io_DOUT_reg_6_ ( .D(top_core_io_N96), .CK(n_CLK), .RN(
        n_RSTB), .Q(n_DOUT[6]) );
  DFFRHQX1 top_core_io_DOUT_reg_7_ ( .D(top_core_io_N97), .CK(n_CLK), .RN(
        n_RSTB), .Q(n_DOUT[7]) );
  DFFHQX1 top_core_KE_CipherKey0_reg_64_ ( .D(top_core_CipherKey[64]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_64_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_65_ ( .D(top_core_CipherKey[65]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_65_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_66_ ( .D(top_core_CipherKey[66]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_66_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_67_ ( .D(top_core_CipherKey[67]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_67_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_68_ ( .D(top_core_CipherKey[68]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_68_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_69_ ( .D(top_core_CipherKey[69]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_69_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_70_ ( .D(top_core_CipherKey[70]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_70_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_71_ ( .D(top_core_CipherKey[71]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_71_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_72_ ( .D(top_core_CipherKey[72]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_72_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_73_ ( .D(top_core_CipherKey[73]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_73_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_74_ ( .D(top_core_CipherKey[74]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_74_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_75_ ( .D(top_core_CipherKey[75]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_75_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_76_ ( .D(top_core_CipherKey[76]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_76_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_77_ ( .D(top_core_CipherKey[77]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_77_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_78_ ( .D(top_core_CipherKey[78]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_78_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_79_ ( .D(top_core_CipherKey[79]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_79_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_80_ ( .D(top_core_CipherKey[80]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_80_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_81_ ( .D(top_core_CipherKey[81]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_81_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_82_ ( .D(top_core_CipherKey[82]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_82_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_83_ ( .D(top_core_CipherKey[83]), .CK(
        n3690), .Q(top_core_KE_CipherKey0_83_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_84_ ( .D(top_core_CipherKey[84]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_84_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_85_ ( .D(top_core_CipherKey[85]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_85_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_86_ ( .D(top_core_CipherKey[86]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_86_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_87_ ( .D(top_core_CipherKey[87]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_87_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_112_ ( .D(top_core_CipherKey[112]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_112_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_113_ ( .D(top_core_CipherKey[113]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_113_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_114_ ( .D(top_core_CipherKey[114]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_114_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_115_ ( .D(top_core_CipherKey[115]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_115_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_116_ ( .D(top_core_CipherKey[116]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_116_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_117_ ( .D(top_core_CipherKey[117]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_117_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_118_ ( .D(top_core_CipherKey[118]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_118_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_119_ ( .D(top_core_CipherKey[119]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_119_) );
  DFFRHQX1 top_core_KE_key_mem_ctrl_reg_reg_1_ ( .D(top_core_KE_n4932), .CK(
        n3848), .RN(n_RSTB), .Q(top_core_KE_key_mem_ctrl_reg_1_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_128_ ( .D(top_core_CipherKey[128]), .CK(
        n3704), .Q(top_core_KE_CipherKey0_128_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_129_ ( .D(top_core_CipherKey[129]), .CK(
        n3704), .Q(top_core_KE_CipherKey0_129_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_130_ ( .D(top_core_CipherKey[130]), .CK(
        n3704), .Q(top_core_KE_CipherKey0_130_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_131_ ( .D(top_core_CipherKey[131]), .CK(
        n3704), .Q(top_core_KE_CipherKey0_131_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_132_ ( .D(top_core_CipherKey[132]), .CK(
        n3704), .Q(top_core_KE_CipherKey0_132_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_133_ ( .D(top_core_CipherKey[133]), .CK(
        n3704), .Q(top_core_KE_CipherKey0_133_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_134_ ( .D(top_core_CipherKey[134]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_134_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_135_ ( .D(top_core_CipherKey[135]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_135_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_136_ ( .D(top_core_CipherKey[136]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_136_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_137_ ( .D(top_core_CipherKey[137]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_137_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_138_ ( .D(top_core_CipherKey[138]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_138_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_139_ ( .D(top_core_CipherKey[139]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_139_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_140_ ( .D(top_core_CipherKey[140]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_140_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_141_ ( .D(top_core_CipherKey[141]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_141_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_142_ ( .D(top_core_CipherKey[142]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_142_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_143_ ( .D(top_core_CipherKey[143]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_143_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_144_ ( .D(top_core_CipherKey[144]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_144_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_145_ ( .D(top_core_CipherKey[145]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_145_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_146_ ( .D(top_core_CipherKey[146]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_146_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_147_ ( .D(top_core_CipherKey[147]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_147_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_148_ ( .D(top_core_CipherKey[148]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_148_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_149_ ( .D(top_core_CipherKey[149]), .CK(
        n3703), .Q(top_core_KE_CipherKey0_149_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_150_ ( .D(top_core_CipherKey[150]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_150_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_151_ ( .D(top_core_CipherKey[151]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_151_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_152_ ( .D(top_core_CipherKey[152]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_152_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_153_ ( .D(top_core_CipherKey[153]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_153_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_154_ ( .D(top_core_CipherKey[154]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_154_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_155_ ( .D(top_core_CipherKey[155]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_155_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_156_ ( .D(top_core_CipherKey[156]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_156_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_157_ ( .D(top_core_CipherKey[157]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_157_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_158_ ( .D(top_core_CipherKey[158]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_158_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_159_ ( .D(top_core_CipherKey[159]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_159_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_160_ ( .D(top_core_CipherKey[160]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_160_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_161_ ( .D(top_core_CipherKey[161]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_161_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_162_ ( .D(top_core_CipherKey[162]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_162_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_163_ ( .D(top_core_CipherKey[163]), .CK(
        n3702), .Q(top_core_KE_CipherKey0_163_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_164_ ( .D(top_core_CipherKey[164]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_164_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_165_ ( .D(top_core_CipherKey[165]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_165_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_166_ ( .D(top_core_CipherKey[166]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_166_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_167_ ( .D(top_core_CipherKey[167]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_167_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_168_ ( .D(top_core_CipherKey[168]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_168_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_169_ ( .D(top_core_CipherKey[169]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_169_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_170_ ( .D(top_core_CipherKey[170]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_170_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_171_ ( .D(top_core_CipherKey[171]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_171_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_172_ ( .D(top_core_CipherKey[172]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_172_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_173_ ( .D(top_core_CipherKey[173]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_173_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_174_ ( .D(top_core_CipherKey[174]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_174_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_175_ ( .D(top_core_CipherKey[175]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_175_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_176_ ( .D(top_core_CipherKey[176]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_176_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_177_ ( .D(top_core_CipherKey[177]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_177_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_178_ ( .D(top_core_CipherKey[178]), .CK(
        n3701), .Q(top_core_KE_CipherKey0_178_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_179_ ( .D(top_core_CipherKey[179]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_179_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_180_ ( .D(top_core_CipherKey[180]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_180_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_181_ ( .D(top_core_CipherKey[181]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_181_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_182_ ( .D(top_core_CipherKey[182]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_182_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_183_ ( .D(top_core_CipherKey[183]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_183_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_184_ ( .D(top_core_CipherKey[184]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_184_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_185_ ( .D(top_core_CipherKey[185]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_185_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_186_ ( .D(top_core_CipherKey[186]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_186_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_187_ ( .D(top_core_CipherKey[187]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_187_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_188_ ( .D(top_core_CipherKey[188]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_188_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_189_ ( .D(top_core_CipherKey[189]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_189_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_190_ ( .D(top_core_CipherKey[190]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_190_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_191_ ( .D(top_core_CipherKey[191]), .CK(
        n3700), .Q(top_core_KE_CipherKey0_191_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_111_ ( .D(top_core_KE_n4808), .CK(
        n3897), .Q(top_core_KE_prev_key1_reg_111_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_103_ ( .D(top_core_KE_n4816), .CK(
        n3903), .Q(top_core_KE_prev_key1_reg_103_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_102_ ( .D(top_core_KE_n4817), .CK(
        n3905), .Q(top_core_KE_prev_key1_reg_102_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_119_ ( .D(top_core_KE_n4800), .CK(
        n3893), .Q(top_core_KE_prev_key1_reg_119_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_118_ ( .D(top_core_KE_n4801), .CK(
        n3896), .Q(top_core_KE_prev_key1_reg_118_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_117_ ( .D(top_core_KE_n4802), .CK(
        n3894), .Q(top_core_KE_prev_key1_reg_117_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_116_ ( .D(top_core_KE_n4803), .CK(
        n3892), .Q(top_core_KE_prev_key1_reg_116_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_115_ ( .D(top_core_KE_n4804), .CK(
        n3904), .Q(top_core_KE_prev_key1_reg_115_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_114_ ( .D(top_core_KE_n4805), .CK(
        n3901), .Q(top_core_KE_prev_key1_reg_114_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_113_ ( .D(top_core_KE_n4806), .CK(
        n3897), .Q(top_core_KE_prev_key1_reg_113_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_112_ ( .D(top_core_KE_n4807), .CK(
        n3898), .Q(top_core_KE_prev_key1_reg_112_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_110_ ( .D(top_core_KE_n4809), .CK(
        n3899), .Q(top_core_KE_prev_key1_reg_110_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_101_ ( .D(top_core_KE_n4818), .CK(
        n3900), .Q(top_core_KE_prev_key1_reg_101_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_109_ ( .D(top_core_KE_n4810), .CK(
        n3901), .Q(top_core_KE_prev_key1_reg_109_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_100_ ( .D(top_core_KE_n4819), .CK(
        n3902), .Q(top_core_KE_prev_key1_reg_100_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_108_ ( .D(top_core_KE_n4811), .CK(
        n3903), .Q(top_core_KE_prev_key1_reg_108_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_99_ ( .D(top_core_KE_n4820), .CK(n3904), .Q(top_core_KE_prev_key1_reg_99_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_107_ ( .D(top_core_KE_n4812), .CK(
        n3905), .Q(top_core_KE_prev_key1_reg_107_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_98_ ( .D(top_core_KE_n4821), .CK(n3906), .Q(top_core_KE_prev_key1_reg_98_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_106_ ( .D(top_core_KE_n4813), .CK(
        n3891), .Q(top_core_KE_prev_key1_reg_106_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_97_ ( .D(top_core_KE_n4822), .CK(n3892), .Q(top_core_KE_prev_key1_reg_97_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_105_ ( .D(top_core_KE_n4814), .CK(
        n3893), .Q(top_core_KE_prev_key1_reg_105_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_96_ ( .D(top_core_KE_n4823), .CK(n3894), .Q(top_core_KE_prev_key1_reg_96_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_104_ ( .D(top_core_KE_n4815), .CK(
        n3895), .Q(top_core_KE_prev_key1_reg_104_) );
  DFFRHQX1 top_core_io_Plain_text_reg_0_ ( .D(top_core_io_N131), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_Plain_text[0]) );
  DFFRHQX1 top_core_io_Plain_text_reg_1_ ( .D(top_core_io_N132), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_Plain_text[1]) );
  DFFRHQX1 top_core_io_Plain_text_reg_2_ ( .D(top_core_io_N133), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_Plain_text[2]) );
  DFFRHQX1 top_core_io_Plain_text_reg_3_ ( .D(top_core_io_N134), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_Plain_text[3]) );
  DFFRHQX1 top_core_io_Plain_text_reg_4_ ( .D(top_core_io_N135), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_Plain_text[4]) );
  DFFRHQX1 top_core_io_Plain_text_reg_5_ ( .D(top_core_io_N136), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[5]) );
  DFFRHQX1 top_core_io_Plain_text_reg_6_ ( .D(top_core_io_N137), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[6]) );
  DFFRHQX1 top_core_io_Plain_text_reg_7_ ( .D(top_core_io_N138), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[7]) );
  DFFRHQX1 top_core_io_Plain_text_reg_8_ ( .D(top_core_io_N139), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[8]) );
  DFFRHQX1 top_core_io_Plain_text_reg_9_ ( .D(top_core_io_N140), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[9]) );
  DFFRHQX1 top_core_io_Plain_text_reg_10_ ( .D(top_core_io_N141), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[10]) );
  DFFRHQX1 top_core_io_Plain_text_reg_11_ ( .D(top_core_io_N142), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[11]) );
  DFFRHQX1 top_core_io_Plain_text_reg_12_ ( .D(top_core_io_N143), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[12]) );
  DFFRHQX1 top_core_io_Plain_text_reg_13_ ( .D(top_core_io_N144), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[13]) );
  DFFRHQX1 top_core_io_Plain_text_reg_14_ ( .D(top_core_io_N145), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[14]) );
  DFFRHQX1 top_core_io_Plain_text_reg_15_ ( .D(top_core_io_N146), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[15]) );
  DFFRHQX1 top_core_io_Plain_text_reg_16_ ( .D(top_core_io_N147), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[16]) );
  DFFRHQX1 top_core_io_Plain_text_reg_17_ ( .D(top_core_io_N148), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[17]) );
  DFFRHQX1 top_core_io_Plain_text_reg_18_ ( .D(top_core_io_N149), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[18]) );
  DFFRHQX1 top_core_io_Plain_text_reg_19_ ( .D(top_core_io_N150), .CK(n3770), 
        .RN(n_RSTB), .Q(top_core_Plain_text[19]) );
  DFFRHQX1 top_core_io_Plain_text_reg_20_ ( .D(top_core_io_N151), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[20]) );
  DFFRHQX1 top_core_io_Plain_text_reg_21_ ( .D(top_core_io_N152), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[21]) );
  DFFRHQX1 top_core_io_Plain_text_reg_22_ ( .D(top_core_io_N153), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[22]) );
  DFFRHQX1 top_core_io_Plain_text_reg_23_ ( .D(top_core_io_N154), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[23]) );
  DFFRHQX1 top_core_io_Plain_text_reg_24_ ( .D(top_core_io_N155), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[24]) );
  DFFRHQX1 top_core_io_Plain_text_reg_25_ ( .D(top_core_io_N156), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[25]) );
  DFFRHQX1 top_core_io_Plain_text_reg_26_ ( .D(top_core_io_N157), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[26]) );
  DFFRHQX1 top_core_io_Plain_text_reg_27_ ( .D(top_core_io_N158), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[27]) );
  DFFRHQX1 top_core_io_Plain_text_reg_28_ ( .D(top_core_io_N159), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[28]) );
  DFFRHQX1 top_core_io_Plain_text_reg_29_ ( .D(top_core_io_N160), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[29]) );
  DFFRHQX1 top_core_io_Plain_text_reg_30_ ( .D(top_core_io_N161), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[30]) );
  DFFRHQX1 top_core_io_Plain_text_reg_31_ ( .D(top_core_io_N162), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[31]) );
  DFFRHQX1 top_core_io_Plain_text_reg_32_ ( .D(top_core_io_N163), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[32]) );
  DFFRHQX1 top_core_io_Plain_text_reg_33_ ( .D(top_core_io_N164), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[33]) );
  DFFRHQX1 top_core_io_Plain_text_reg_34_ ( .D(top_core_io_N165), .CK(n3771), 
        .RN(n_RSTB), .Q(top_core_Plain_text[34]) );
  DFFRHQX1 top_core_io_Plain_text_reg_35_ ( .D(top_core_io_N166), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[35]) );
  DFFRHQX1 top_core_io_Plain_text_reg_36_ ( .D(top_core_io_N167), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[36]) );
  DFFRHQX1 top_core_io_Plain_text_reg_37_ ( .D(top_core_io_N168), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[37]) );
  DFFRHQX1 top_core_io_Plain_text_reg_38_ ( .D(top_core_io_N169), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[38]) );
  DFFRHQX1 top_core_io_Plain_text_reg_39_ ( .D(top_core_io_N170), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[39]) );
  DFFRHQX1 top_core_io_Plain_text_reg_40_ ( .D(top_core_io_N171), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[40]) );
  DFFRHQX1 top_core_io_Plain_text_reg_41_ ( .D(top_core_io_N172), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[41]) );
  DFFRHQX1 top_core_io_Plain_text_reg_42_ ( .D(top_core_io_N173), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[42]) );
  DFFRHQX1 top_core_io_Plain_text_reg_43_ ( .D(top_core_io_N174), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[43]) );
  DFFRHQX1 top_core_io_Plain_text_reg_44_ ( .D(top_core_io_N175), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[44]) );
  DFFRHQX1 top_core_io_Plain_text_reg_45_ ( .D(top_core_io_N176), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[45]) );
  DFFRHQX1 top_core_io_Plain_text_reg_46_ ( .D(top_core_io_N177), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[46]) );
  DFFRHQX1 top_core_io_Plain_text_reg_47_ ( .D(top_core_io_N178), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[47]) );
  DFFRHQX1 top_core_io_Plain_text_reg_48_ ( .D(top_core_io_N179), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[48]) );
  DFFRHQX1 top_core_io_Plain_text_reg_49_ ( .D(top_core_io_N180), .CK(n3772), 
        .RN(n_RSTB), .Q(top_core_Plain_text[49]) );
  DFFRHQX1 top_core_io_Plain_text_reg_50_ ( .D(top_core_io_N181), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[50]) );
  DFFRHQX1 top_core_io_Plain_text_reg_51_ ( .D(top_core_io_N182), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[51]) );
  DFFRHQX1 top_core_io_Plain_text_reg_52_ ( .D(top_core_io_N183), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[52]) );
  DFFRHQX1 top_core_io_Plain_text_reg_53_ ( .D(top_core_io_N184), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[53]) );
  DFFRHQX1 top_core_io_Plain_text_reg_54_ ( .D(top_core_io_N185), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[54]) );
  DFFRHQX1 top_core_io_Plain_text_reg_55_ ( .D(top_core_io_N186), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[55]) );
  DFFRHQX1 top_core_io_Plain_text_reg_56_ ( .D(top_core_io_N187), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[56]) );
  DFFRHQX1 top_core_io_Plain_text_reg_57_ ( .D(top_core_io_N188), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[57]) );
  DFFRHQX1 top_core_io_Plain_text_reg_58_ ( .D(top_core_io_N189), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[58]) );
  DFFRHQX1 top_core_io_Plain_text_reg_59_ ( .D(top_core_io_N190), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[59]) );
  DFFRHQX1 top_core_io_Plain_text_reg_60_ ( .D(top_core_io_N191), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[60]) );
  DFFRHQX1 top_core_io_Plain_text_reg_61_ ( .D(top_core_io_N192), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[61]) );
  DFFRHQX1 top_core_io_Plain_text_reg_62_ ( .D(top_core_io_N193), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[62]) );
  DFFRHQX1 top_core_io_Plain_text_reg_63_ ( .D(top_core_io_N194), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[63]) );
  DFFRHQX1 top_core_io_Plain_text_reg_66_ ( .D(top_core_io_N197), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[66]) );
  DFFRHQX1 top_core_io_Plain_text_reg_67_ ( .D(top_core_io_N198), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[67]) );
  DFFRHQX1 top_core_io_Plain_text_reg_68_ ( .D(top_core_io_N199), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[68]) );
  DFFRHQX1 top_core_io_Plain_text_reg_69_ ( .D(top_core_io_N200), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[69]) );
  DFFRHQX1 top_core_io_Plain_text_reg_70_ ( .D(top_core_io_N201), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[70]) );
  DFFRHQX1 top_core_io_Plain_text_reg_71_ ( .D(top_core_io_N202), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[71]) );
  DFFRHQX1 top_core_KE_rcon_reg_reg_6_ ( .D(top_core_KE_n4921), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_rcon_reg_6_) );
  DFFRHQX1 top_core_KE_rcon_reg_reg_5_ ( .D(top_core_KE_n4922), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_rcon_reg_5_) );
  DFFRHQX1 top_core_KE_rcon_reg_reg_4_ ( .D(top_core_KE_n4923), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_rcon_reg_4_) );
  DFFRHQX1 top_core_KE_rcon_reg_reg_1_ ( .D(top_core_KE_n4926), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_rcon_reg_1_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_127_ ( .D(top_core_CipherKey[127]), .CK(
        n3704), .Q(top_core_KE_CipherKey0_127_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_127_ ( .D(top_core_EC_n1163), .CK(
        n3787), .RN(n_RSTB), .Q(top_core_EC_round_result_r_127_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_126_ ( .D(top_core_EC_n1164), .CK(
        n3787), .RN(n_RSTB), .Q(top_core_EC_round_result_r_126_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_125_ ( .D(top_core_EC_n1165), .CK(
        n3787), .RN(n_RSTB), .Q(top_core_EC_round_result_r_125_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_124_ ( .D(top_core_EC_n1166), .CK(
        n3787), .RN(n_RSTB), .Q(top_core_EC_round_result_r_124_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_123_ ( .D(top_core_EC_n1167), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_123_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_122_ ( .D(top_core_EC_n1168), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_122_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_121_ ( .D(top_core_EC_n1169), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_121_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_120_ ( .D(top_core_EC_n1170), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_120_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_119_ ( .D(top_core_EC_n1171), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_119_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_118_ ( .D(top_core_EC_n1172), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_118_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_117_ ( .D(top_core_EC_n1173), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_117_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_116_ ( .D(top_core_EC_n1174), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_116_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_115_ ( .D(top_core_EC_n1175), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_115_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_114_ ( .D(top_core_EC_n1176), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_114_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_113_ ( .D(top_core_EC_n1177), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_113_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_112_ ( .D(top_core_EC_n1178), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_112_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_111_ ( .D(top_core_EC_n1179), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_111_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_110_ ( .D(top_core_EC_n1180), .CK(
        n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_r_110_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_109_ ( .D(top_core_EC_n1181), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_109_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_108_ ( .D(top_core_EC_n1182), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_108_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_107_ ( .D(top_core_EC_n1183), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_107_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_106_ ( .D(top_core_EC_n1184), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_106_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_105_ ( .D(top_core_EC_n1185), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_105_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_104_ ( .D(top_core_EC_n1186), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_104_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_103_ ( .D(top_core_EC_n1187), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_103_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_102_ ( .D(top_core_EC_n1188), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_102_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_101_ ( .D(top_core_EC_n1189), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_101_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_100_ ( .D(top_core_EC_n1190), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_100_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_99_ ( .D(top_core_EC_n1191), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_99_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_98_ ( .D(top_core_EC_n1192), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_98_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_97_ ( .D(top_core_EC_n1193), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_97_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_96_ ( .D(top_core_EC_n1194), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_96_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_95_ ( .D(top_core_EC_n1195), .CK(
        n3789), .RN(n_RSTB), .Q(top_core_EC_round_result_r_95_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_94_ ( .D(top_core_EC_n1196), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_94_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_93_ ( .D(top_core_EC_n1197), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_93_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_92_ ( .D(top_core_EC_n1198), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_92_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_91_ ( .D(top_core_EC_n1199), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_91_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_90_ ( .D(top_core_EC_n1200), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_90_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_89_ ( .D(top_core_EC_n1201), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_89_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_88_ ( .D(top_core_EC_n1202), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_88_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_87_ ( .D(top_core_EC_n1203), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_87_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_86_ ( .D(top_core_EC_n1204), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_86_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_85_ ( .D(top_core_EC_n1205), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_85_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_84_ ( .D(top_core_EC_n1206), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_84_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_83_ ( .D(top_core_EC_n1207), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_83_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_82_ ( .D(top_core_EC_n1208), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_82_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_81_ ( .D(top_core_EC_n1209), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_81_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_80_ ( .D(top_core_EC_n1210), .CK(
        n3790), .RN(n_RSTB), .Q(top_core_EC_round_result_r_80_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_79_ ( .D(top_core_EC_n1211), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_79_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_78_ ( .D(top_core_EC_n1212), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_78_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_77_ ( .D(top_core_EC_n1213), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_77_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_76_ ( .D(top_core_EC_n1214), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_76_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_75_ ( .D(top_core_EC_n1215), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_75_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_74_ ( .D(top_core_EC_n1216), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_74_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_73_ ( .D(top_core_EC_n1217), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_73_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_72_ ( .D(top_core_EC_n1218), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_72_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_71_ ( .D(top_core_EC_n1219), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_71_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_70_ ( .D(top_core_EC_n1220), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_70_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_69_ ( .D(top_core_EC_n1221), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_69_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_68_ ( .D(top_core_EC_n1222), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_68_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_67_ ( .D(top_core_EC_n1223), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_67_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_66_ ( .D(top_core_EC_n1224), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_66_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_65_ ( .D(top_core_EC_n1225), .CK(
        n3791), .RN(n_RSTB), .Q(top_core_EC_round_result_r_65_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_64_ ( .D(top_core_EC_n1226), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_64_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_63_ ( .D(top_core_EC_n1227), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_63_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_62_ ( .D(top_core_EC_n1228), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_62_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_61_ ( .D(top_core_EC_n1229), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_61_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_60_ ( .D(top_core_EC_n1230), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_60_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_59_ ( .D(top_core_EC_n1231), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_59_) );
  DFFRHQX1 top_core_EC_round_result_r_reg_58_ ( .D(top_core_EC_n1232), .CK(
        n3792), .RN(n_RSTB), .Q(top_core_EC_round_result_r_58_) );
  DFFRHQX1 top_core_io_Plain_text_reg_64_ ( .D(top_core_io_N195), .CK(n3773), 
        .RN(n_RSTB), .Q(top_core_Plain_text[64]) );
  DFFRHQX1 top_core_io_Plain_text_reg_65_ ( .D(top_core_io_N196), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[65]) );
  DFFRHQX1 top_core_io_Plain_text_reg_72_ ( .D(top_core_io_N203), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[72]) );
  DFFRHQX1 top_core_io_Plain_text_reg_73_ ( .D(top_core_io_N204), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[73]) );
  DFFRHQX1 top_core_io_Plain_text_reg_74_ ( .D(top_core_io_N205), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[74]) );
  DFFRHQX1 top_core_io_Plain_text_reg_75_ ( .D(top_core_io_N206), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[75]) );
  DFFRHQX1 top_core_io_Plain_text_reg_76_ ( .D(top_core_io_N207), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[76]) );
  DFFRHQX1 top_core_io_Plain_text_reg_77_ ( .D(top_core_io_N208), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[77]) );
  DFFRHQX1 top_core_io_Plain_text_reg_78_ ( .D(top_core_io_N209), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[78]) );
  DFFRHQX1 top_core_io_Plain_text_reg_79_ ( .D(top_core_io_N210), .CK(n3774), 
        .RN(n_RSTB), .Q(top_core_Plain_text[79]) );
  DFFRHQX1 top_core_io_Plain_text_reg_80_ ( .D(top_core_io_N211), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[80]) );
  DFFRHQX1 top_core_io_Plain_text_reg_81_ ( .D(top_core_io_N212), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[81]) );
  DFFRHQX1 top_core_io_Plain_text_reg_82_ ( .D(top_core_io_N213), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[82]) );
  DFFRHQX1 top_core_io_Plain_text_reg_83_ ( .D(top_core_io_N214), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[83]) );
  DFFRHQX1 top_core_io_Plain_text_reg_84_ ( .D(top_core_io_N215), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[84]) );
  DFFRHQX1 top_core_io_Plain_text_reg_85_ ( .D(top_core_io_N216), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[85]) );
  DFFRHQX1 top_core_io_Plain_text_reg_86_ ( .D(top_core_io_N217), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[86]) );
  DFFRHQX1 top_core_io_Plain_text_reg_87_ ( .D(top_core_io_N218), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[87]) );
  DFFRHQX1 top_core_io_Plain_text_reg_88_ ( .D(top_core_io_N219), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[88]) );
  DFFRHQX1 top_core_io_Plain_text_reg_89_ ( .D(top_core_io_N220), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[89]) );
  DFFRHQX1 top_core_io_Plain_text_reg_90_ ( .D(top_core_io_N221), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[90]) );
  DFFRHQX1 top_core_io_Plain_text_reg_91_ ( .D(top_core_io_N222), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[91]) );
  DFFRHQX1 top_core_io_Plain_text_reg_92_ ( .D(top_core_io_N223), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[92]) );
  DFFRHQX1 top_core_io_Plain_text_reg_93_ ( .D(top_core_io_N224), .CK(n3775), 
        .RN(n_RSTB), .Q(top_core_Plain_text[93]) );
  DFFRHQX1 top_core_io_Plain_text_reg_94_ ( .D(top_core_io_N225), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[94]) );
  DFFRHQX1 top_core_io_Plain_text_reg_95_ ( .D(top_core_io_N226), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[95]) );
  DFFRHQX1 top_core_io_Plain_text_reg_96_ ( .D(top_core_io_N227), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[96]) );
  DFFRHQX1 top_core_io_Plain_text_reg_97_ ( .D(top_core_io_N228), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[97]) );
  DFFRHQX1 top_core_io_Plain_text_reg_98_ ( .D(top_core_io_N229), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[98]) );
  DFFRHQX1 top_core_io_Plain_text_reg_99_ ( .D(top_core_io_N230), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[99]) );
  DFFRHQX1 top_core_io_Plain_text_reg_100_ ( .D(top_core_io_N231), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[100]) );
  DFFRHQX1 top_core_io_Plain_text_reg_101_ ( .D(top_core_io_N232), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[101]) );
  DFFRHQX1 top_core_io_Plain_text_reg_102_ ( .D(top_core_io_N233), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[102]) );
  DFFRHQX1 top_core_io_Plain_text_reg_103_ ( .D(top_core_io_N234), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[103]) );
  DFFRHQX1 top_core_io_Plain_text_reg_104_ ( .D(top_core_io_N235), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[104]) );
  DFFRHQX1 top_core_io_Plain_text_reg_105_ ( .D(top_core_io_N236), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[105]) );
  DFFRHQX1 top_core_io_Plain_text_reg_106_ ( .D(top_core_io_N237), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[106]) );
  DFFRHQX1 top_core_io_Plain_text_reg_107_ ( .D(top_core_io_N238), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[107]) );
  DFFRHQX1 top_core_io_Plain_text_reg_108_ ( .D(top_core_io_N239), .CK(n3776), 
        .RN(n_RSTB), .Q(top_core_Plain_text[108]) );
  DFFRHQX1 top_core_io_Plain_text_reg_109_ ( .D(top_core_io_N240), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[109]) );
  DFFRHQX1 top_core_io_Plain_text_reg_110_ ( .D(top_core_io_N241), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[110]) );
  DFFRHQX1 top_core_io_Plain_text_reg_111_ ( .D(top_core_io_N242), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[111]) );
  DFFRHQX1 top_core_io_Plain_text_reg_112_ ( .D(top_core_io_N243), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[112]) );
  DFFRHQX1 top_core_io_Plain_text_reg_113_ ( .D(top_core_io_N244), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[113]) );
  DFFRHQX1 top_core_io_Plain_text_reg_114_ ( .D(top_core_io_N245), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[114]) );
  DFFRHQX1 top_core_io_Plain_text_reg_115_ ( .D(top_core_io_N246), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[115]) );
  DFFRHQX1 top_core_io_Plain_text_reg_116_ ( .D(top_core_io_N247), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[116]) );
  DFFRHQX1 top_core_io_Plain_text_reg_117_ ( .D(top_core_io_N248), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[117]) );
  DFFRHQX1 top_core_io_Plain_text_reg_118_ ( .D(top_core_io_N249), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[118]) );
  DFFRHQX1 top_core_io_Plain_text_reg_119_ ( .D(top_core_io_N250), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[119]) );
  DFFRHQX1 top_core_io_Plain_text_reg_120_ ( .D(top_core_io_N251), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[120]) );
  DFFRHQX1 top_core_io_Plain_text_reg_121_ ( .D(top_core_io_N252), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[121]) );
  DFFRHQX1 top_core_io_Plain_text_reg_122_ ( .D(top_core_io_N253), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[122]) );
  DFFRHQX1 top_core_io_Plain_text_reg_123_ ( .D(top_core_io_N254), .CK(n3777), 
        .RN(n_RSTB), .Q(top_core_Plain_text[123]) );
  DFFRHQX1 top_core_io_Plain_text_reg_124_ ( .D(top_core_io_N255), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_Plain_text[124]) );
  DFFRHQX1 top_core_io_Plain_text_reg_125_ ( .D(top_core_io_N256), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_Plain_text[125]) );
  DFFRHQX1 top_core_io_Plain_text_reg_126_ ( .D(top_core_io_N257), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_Plain_text[126]) );
  DFFRHQX1 top_core_io_Plain_text_reg_127_ ( .D(top_core_io_N258), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_Plain_text[127]) );
  DFFHQX1 top_core_KE_CipherKey0_reg_88_ ( .D(top_core_CipherKey[88]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_88_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_89_ ( .D(top_core_CipherKey[89]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_89_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_90_ ( .D(top_core_CipherKey[90]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_90_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_91_ ( .D(top_core_CipherKey[91]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_91_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_92_ ( .D(top_core_CipherKey[92]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_92_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_93_ ( .D(top_core_CipherKey[93]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_93_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_94_ ( .D(top_core_CipherKey[94]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_94_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_95_ ( .D(top_core_CipherKey[95]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_95_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_96_ ( .D(top_core_CipherKey[96]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_96_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_97_ ( .D(top_core_CipherKey[97]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_97_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_98_ ( .D(top_core_CipherKey[98]), .CK(
        n3689), .Q(top_core_KE_CipherKey0_98_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_99_ ( .D(top_core_CipherKey[99]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_99_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_100_ ( .D(top_core_CipherKey[100]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_100_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_101_ ( .D(top_core_CipherKey[101]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_101_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_102_ ( .D(top_core_CipherKey[102]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_102_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_103_ ( .D(top_core_CipherKey[103]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_103_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_104_ ( .D(top_core_CipherKey[104]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_104_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_105_ ( .D(top_core_CipherKey[105]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_105_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_106_ ( .D(top_core_CipherKey[106]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_106_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_107_ ( .D(top_core_CipherKey[107]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_107_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_108_ ( .D(top_core_CipherKey[108]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_108_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_109_ ( .D(top_core_CipherKey[109]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_109_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_110_ ( .D(top_core_CipherKey[110]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_110_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_111_ ( .D(top_core_CipherKey[111]), .CK(
        n3688), .Q(top_core_KE_CipherKey0_111_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_120_ ( .D(top_core_CipherKey[120]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_120_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_121_ ( .D(top_core_CipherKey[121]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_121_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_122_ ( .D(top_core_CipherKey[122]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_122_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_123_ ( .D(top_core_CipherKey[123]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_123_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_124_ ( .D(top_core_CipherKey[124]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_124_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_125_ ( .D(top_core_CipherKey[125]), .CK(
        n3687), .Q(top_core_KE_CipherKey0_125_) );
  DFFHQX1 top_core_KE_CipherKey0_reg_126_ ( .D(top_core_CipherKey[126]), .CK(
        n3691), .Q(top_core_KE_CipherKey0_126_) );
  DFFRHQX1 top_core_EC_round_result_reg_127_ ( .D(top_core_EC_n1035), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_127_) );
  DFFRHQX1 top_core_EC_round_result_reg_126_ ( .D(top_core_EC_n1036), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_126_) );
  DFFRHQX1 top_core_EC_round_result_reg_125_ ( .D(top_core_EC_n1037), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_125_) );
  DFFRHQX1 top_core_EC_round_result_reg_124_ ( .D(top_core_EC_n1038), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_124_) );
  DFFRHQX1 top_core_EC_round_result_reg_123_ ( .D(top_core_EC_n1039), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_123_) );
  DFFRHQX1 top_core_EC_round_result_reg_122_ ( .D(top_core_EC_n1040), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_122_) );
  DFFRHQX1 top_core_EC_round_result_reg_121_ ( .D(top_core_EC_n1041), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_121_) );
  DFFRHQX1 top_core_EC_round_result_reg_120_ ( .D(top_core_EC_n1042), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_120_) );
  DFFRHQX1 top_core_EC_round_result_reg_119_ ( .D(top_core_EC_n1043), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_119_) );
  DFFRHQX1 top_core_EC_round_result_reg_118_ ( .D(top_core_EC_n1044), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_118_) );
  DFFRHQX1 top_core_EC_round_result_reg_117_ ( .D(top_core_EC_n1045), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_117_) );
  DFFRHQX1 top_core_EC_round_result_reg_116_ ( .D(top_core_EC_n1046), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_116_) );
  DFFRHQX1 top_core_EC_round_result_reg_115_ ( .D(top_core_EC_n1047), .CK(
        n3804), .RN(n_RSTB), .Q(top_core_EC_round_result_115_) );
  DFFRHQX1 top_core_EC_round_result_reg_114_ ( .D(top_core_EC_n1048), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_114_) );
  DFFRHQX1 top_core_EC_round_result_reg_113_ ( .D(top_core_EC_n1049), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_113_) );
  DFFRHQX1 top_core_EC_round_result_reg_112_ ( .D(top_core_EC_n1050), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_112_) );
  DFFRHQX1 top_core_EC_round_result_reg_111_ ( .D(top_core_EC_n1051), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_111_) );
  DFFRHQX1 top_core_EC_round_result_reg_110_ ( .D(top_core_EC_n1052), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_110_) );
  DFFRHQX1 top_core_EC_round_result_reg_109_ ( .D(top_core_EC_n1053), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_109_) );
  DFFRHQX1 top_core_EC_round_result_reg_108_ ( .D(top_core_EC_n1054), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_108_) );
  DFFRHQX1 top_core_EC_round_result_reg_107_ ( .D(top_core_EC_n1055), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_107_) );
  DFFRHQX1 top_core_EC_round_result_reg_106_ ( .D(top_core_EC_n1056), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_106_) );
  DFFRHQX1 top_core_EC_round_result_reg_105_ ( .D(top_core_EC_n1057), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_105_) );
  DFFRHQX1 top_core_EC_round_result_reg_104_ ( .D(top_core_EC_n1058), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_104_) );
  DFFRHQX1 top_core_EC_round_result_reg_103_ ( .D(top_core_EC_n1059), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_103_) );
  DFFRHQX1 top_core_EC_round_result_reg_102_ ( .D(top_core_EC_n1060), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_102_) );
  DFFRHQX1 top_core_EC_round_result_reg_101_ ( .D(top_core_EC_n1061), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_101_) );
  DFFRHQX1 top_core_EC_round_result_reg_100_ ( .D(top_core_EC_n1062), .CK(
        n3805), .RN(n_RSTB), .Q(top_core_EC_round_result_100_) );
  DFFRHQX1 top_core_EC_round_result_reg_99_ ( .D(top_core_EC_n1063), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_99_) );
  DFFRHQX1 top_core_EC_round_result_reg_98_ ( .D(top_core_EC_n1064), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_98_) );
  DFFRHQX1 top_core_EC_round_result_reg_97_ ( .D(top_core_EC_n1065), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_97_) );
  DFFRHQX1 top_core_EC_round_result_reg_96_ ( .D(top_core_EC_n1066), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_96_) );
  DFFRHQX1 top_core_EC_round_result_reg_95_ ( .D(top_core_EC_n1067), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_95_) );
  DFFRHQX1 top_core_EC_round_result_reg_94_ ( .D(top_core_EC_n1068), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_94_) );
  DFFRHQX1 top_core_EC_round_result_reg_93_ ( .D(top_core_EC_n1069), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_93_) );
  DFFRHQX1 top_core_EC_round_result_reg_92_ ( .D(top_core_EC_n1070), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_92_) );
  DFFRHQX1 top_core_EC_round_result_reg_91_ ( .D(top_core_EC_n1071), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_91_) );
  DFFRHQX1 top_core_EC_round_result_reg_90_ ( .D(top_core_EC_n1072), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_90_) );
  DFFRHQX1 top_core_EC_round_result_reg_89_ ( .D(top_core_EC_n1073), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_89_) );
  DFFRHQX1 top_core_EC_round_result_reg_88_ ( .D(top_core_EC_n1074), .CK(n3806), .RN(n_RSTB), .Q(top_core_EC_round_result_88_) );
  DFFRHQX1 top_core_EC_round_result_reg_87_ ( .D(top_core_EC_n1075), .CK(n3788), .RN(n_RSTB), .Q(top_core_EC_round_result_87_) );
  DFFRHQX1 top_core_EC_round_result_reg_86_ ( .D(top_core_EC_n1076), .CK(n3781), .RN(n_RSTB), .Q(top_core_EC_round_result_86_) );
  DFFRHQX1 top_core_EC_round_result_reg_85_ ( .D(top_core_EC_n1077), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_85_) );
  DFFRHQX1 top_core_EC_round_result_reg_84_ ( .D(top_core_EC_n1078), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_84_) );
  DFFRHQX1 top_core_EC_round_result_reg_83_ ( .D(top_core_EC_n1079), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_83_) );
  DFFRHQX1 top_core_EC_round_result_reg_82_ ( .D(top_core_EC_n1080), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_82_) );
  DFFRHQX1 top_core_EC_round_result_reg_81_ ( .D(top_core_EC_n1081), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_81_) );
  DFFRHQX1 top_core_EC_round_result_reg_80_ ( .D(top_core_EC_n1082), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_80_) );
  DFFRHQX1 top_core_EC_round_result_reg_79_ ( .D(top_core_EC_n1083), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_79_) );
  DFFRHQX1 top_core_EC_round_result_reg_78_ ( .D(top_core_EC_n1084), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_78_) );
  DFFRHQX1 top_core_EC_round_result_reg_77_ ( .D(top_core_EC_n1085), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_77_) );
  DFFRHQX1 top_core_EC_round_result_reg_76_ ( .D(top_core_EC_n1086), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_76_) );
  DFFRHQX1 top_core_EC_round_result_reg_75_ ( .D(top_core_EC_n1087), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_75_) );
  DFFRHQX1 top_core_EC_round_result_reg_74_ ( .D(top_core_EC_n1088), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_74_) );
  DFFRHQX1 top_core_EC_round_result_reg_73_ ( .D(top_core_EC_n1089), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_73_) );
  DFFRHQX1 top_core_EC_round_result_reg_72_ ( .D(top_core_EC_n1090), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_72_) );
  DFFRHQX1 top_core_EC_round_result_reg_71_ ( .D(top_core_EC_n1091), .CK(n3782), .RN(n_RSTB), .Q(top_core_EC_round_result_71_) );
  DFFRHQX1 top_core_EC_round_result_reg_70_ ( .D(top_core_EC_n1092), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_70_) );
  DFFRHQX1 top_core_EC_round_result_reg_69_ ( .D(top_core_EC_n1093), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_69_) );
  DFFRHQX1 top_core_EC_round_result_reg_68_ ( .D(top_core_EC_n1094), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_68_) );
  DFFRHQX1 top_core_EC_round_result_reg_67_ ( .D(top_core_EC_n1095), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_67_) );
  DFFRHQX1 top_core_EC_round_result_reg_66_ ( .D(top_core_EC_n1096), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_66_) );
  DFFRHQX1 top_core_EC_round_result_reg_65_ ( .D(top_core_EC_n1097), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_65_) );
  DFFRHQX1 top_core_EC_round_result_reg_64_ ( .D(top_core_EC_n1098), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_64_) );
  DFFRHQX1 top_core_EC_round_result_reg_63_ ( .D(top_core_EC_n1099), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_63_) );
  DFFRHQX1 top_core_EC_round_result_reg_62_ ( .D(top_core_EC_n1100), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_62_) );
  DFFRHQX1 top_core_EC_round_result_reg_61_ ( .D(top_core_EC_n1101), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_61_) );
  DFFRHQX1 top_core_EC_round_result_reg_60_ ( .D(top_core_EC_n1102), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_60_) );
  DFFRHQX1 top_core_EC_round_result_reg_59_ ( .D(top_core_EC_n1103), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_59_) );
  DFFRHQX1 top_core_EC_round_result_reg_58_ ( .D(top_core_EC_n1104), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_58_) );
  DFFRHQX1 top_core_EC_round_result_reg_57_ ( .D(top_core_EC_n1105), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_57_) );
  DFFRHQX1 top_core_EC_round_result_reg_56_ ( .D(top_core_EC_n1106), .CK(n3783), .RN(n_RSTB), .Q(top_core_EC_round_result_56_) );
  DFFRHQX1 top_core_EC_round_result_reg_55_ ( .D(top_core_EC_n1107), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_55_) );
  DFFRHQX1 top_core_EC_round_result_reg_54_ ( .D(top_core_EC_n1108), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_54_) );
  DFFRHQX1 top_core_EC_round_result_reg_53_ ( .D(top_core_EC_n1109), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_53_) );
  DFFRHQX1 top_core_EC_round_result_reg_52_ ( .D(top_core_EC_n1110), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_52_) );
  DFFRHQX1 top_core_EC_round_result_reg_51_ ( .D(top_core_EC_n1111), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_51_) );
  DFFRHQX1 top_core_EC_round_result_reg_50_ ( .D(top_core_EC_n1112), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_50_) );
  DFFRHQX1 top_core_EC_round_result_reg_49_ ( .D(top_core_EC_n1113), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_49_) );
  DFFRHQX1 top_core_EC_round_result_reg_48_ ( .D(top_core_EC_n1114), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_48_) );
  DFFRHQX1 top_core_EC_round_result_reg_47_ ( .D(top_core_EC_n1115), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_47_) );
  DFFRHQX1 top_core_EC_round_result_reg_46_ ( .D(top_core_EC_n1116), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_46_) );
  DFFRHQX1 top_core_EC_round_result_reg_45_ ( .D(top_core_EC_n1117), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_45_) );
  DFFRHQX1 top_core_EC_round_result_reg_44_ ( .D(top_core_EC_n1118), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_44_) );
  DFFRHQX1 top_core_EC_round_result_reg_43_ ( .D(top_core_EC_n1119), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_43_) );
  DFFRHQX1 top_core_EC_round_result_reg_42_ ( .D(top_core_EC_n1120), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_42_) );
  DFFRHQX1 top_core_EC_round_result_reg_41_ ( .D(top_core_EC_n1121), .CK(n3784), .RN(n_RSTB), .Q(top_core_EC_round_result_41_) );
  DFFRHQX1 top_core_EC_round_result_reg_40_ ( .D(top_core_EC_n1122), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_40_) );
  DFFRHQX1 top_core_EC_round_result_reg_39_ ( .D(top_core_EC_n1123), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_39_) );
  DFFRHQX1 top_core_EC_round_result_reg_38_ ( .D(top_core_EC_n1124), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_38_) );
  DFFRHQX1 top_core_EC_round_result_reg_37_ ( .D(top_core_EC_n1125), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_37_) );
  DFFRHQX1 top_core_EC_round_result_reg_36_ ( .D(top_core_EC_n1126), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_36_) );
  DFFRHQX1 top_core_EC_round_result_reg_35_ ( .D(top_core_EC_n1127), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_35_) );
  DFFRHQX1 top_core_EC_round_result_reg_34_ ( .D(top_core_EC_n1128), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_34_) );
  DFFRHQX1 top_core_EC_round_result_reg_33_ ( .D(top_core_EC_n1129), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_33_) );
  DFFRHQX1 top_core_EC_round_result_reg_32_ ( .D(top_core_EC_n1130), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_32_) );
  DFFRHQX1 top_core_EC_round_result_reg_31_ ( .D(top_core_EC_n1131), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_31_) );
  DFFRHQX1 top_core_EC_round_result_reg_30_ ( .D(top_core_EC_n1132), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_30_) );
  DFFRHQX1 top_core_EC_round_result_reg_29_ ( .D(top_core_EC_n1133), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_29_) );
  DFFRHQX1 top_core_EC_round_result_reg_28_ ( .D(top_core_EC_n1134), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_28_) );
  DFFRHQX1 top_core_EC_round_result_reg_27_ ( .D(top_core_EC_n1135), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_27_) );
  DFFRHQX1 top_core_EC_round_result_reg_26_ ( .D(top_core_EC_n1136), .CK(n3785), .RN(n_RSTB), .Q(top_core_EC_round_result_26_) );
  DFFRHQX1 top_core_EC_round_result_reg_25_ ( .D(top_core_EC_n1137), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_25_) );
  DFFRHQX1 top_core_EC_round_result_reg_24_ ( .D(top_core_EC_n1138), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_24_) );
  DFFRHQX1 top_core_EC_round_result_reg_23_ ( .D(top_core_EC_n1139), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_23_) );
  DFFRHQX1 top_core_EC_round_result_reg_22_ ( .D(top_core_EC_n1140), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_22_) );
  DFFRHQX1 top_core_EC_round_result_reg_21_ ( .D(top_core_EC_n1141), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_21_) );
  DFFRHQX1 top_core_EC_round_result_reg_20_ ( .D(top_core_EC_n1142), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_20_) );
  DFFRHQX1 top_core_EC_round_result_reg_19_ ( .D(top_core_EC_n1143), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_19_) );
  DFFRHQX1 top_core_EC_round_result_reg_18_ ( .D(top_core_EC_n1144), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_18_) );
  DFFRHQX1 top_core_EC_round_result_reg_17_ ( .D(top_core_EC_n1145), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_17_) );
  DFFRHQX1 top_core_EC_round_result_reg_16_ ( .D(top_core_EC_n1146), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_16_) );
  DFFRHQX1 top_core_EC_round_result_reg_15_ ( .D(top_core_EC_n1147), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_15_) );
  DFFRHQX1 top_core_EC_round_result_reg_14_ ( .D(top_core_EC_n1148), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_14_) );
  DFFRHQX1 top_core_EC_round_result_reg_13_ ( .D(top_core_EC_n1149), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_13_) );
  DFFRHQX1 top_core_EC_round_result_reg_12_ ( .D(top_core_EC_n1150), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_12_) );
  DFFRHQX1 top_core_EC_round_result_reg_11_ ( .D(top_core_EC_n1151), .CK(n3786), .RN(n_RSTB), .Q(top_core_EC_round_result_11_) );
  DFFRHQX1 top_core_EC_round_result_reg_10_ ( .D(top_core_EC_n1152), .CK(n3787), .RN(n_RSTB), .Q(top_core_EC_round_result_10_) );
  DFFRHQX1 top_core_EC_round_result_reg_9_ ( .D(top_core_EC_n1153), .CK(n3787), 
        .RN(n_RSTB), .Q(top_core_EC_round_result_9_) );
  DFFRHQX1 top_core_EC_round_result_reg_8_ ( .D(top_core_EC_n1154), .CK(n3787), 
        .RN(n_RSTB), .Q(top_core_EC_round_result_8_) );
  DFFRHQX1 top_core_EC_round_result_reg_7_ ( .D(top_core_EC_n1155), .CK(n3787), 
        .RN(n_RSTB), .Q(top_core_EC_round_result_7_) );
  DFFRHQX1 top_core_EC_round_result_reg_6_ ( .D(top_core_EC_n1156), .CK(n3787), 
        .RN(n_RSTB), .Q(top_core_EC_round_result_6_) );
  DFFRHQX1 top_core_EC_round_result_reg_5_ ( .D(top_core_EC_n1157), .CK(n3787), 
        .RN(n_RSTB), .Q(top_core_EC_round_result_5_) );
  DFFRHQX1 top_core_EC_round_result_reg_4_ ( .D(top_core_EC_n1158), .CK(n3787), 
        .RN(n_RSTB), .Q(top_core_EC_round_result_4_) );
  DFFRHQX1 top_core_EC_round_result_reg_3_ ( .D(top_core_EC_n1159), .CK(n3787), 
        .RN(n_RSTB), .Q(top_core_EC_round_result_3_) );
  DFFRHQX1 top_core_EC_round_result_reg_2_ ( .D(top_core_EC_n1160), .CK(n3787), 
        .RN(n_RSTB), .Q(top_core_EC_round_result_2_) );
  DFFRHQX1 top_core_EC_round_result_reg_1_ ( .D(top_core_EC_n1161), .CK(n3787), 
        .RN(n_RSTB), .Q(top_core_EC_round_result_1_) );
  DFFRHQX1 top_core_EC_round_result_reg_0_ ( .D(top_core_EC_n1162), .CK(n3787), 
        .RN(n_RSTB), .Q(top_core_EC_round_result_0_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_57_ ( .D(top_core_KE_n4862), .CK(n3900), .Q(top_core_KE_prev_key1_reg_57_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_62_ ( .D(top_core_KE_n4857), .CK(n3896), .Q(top_core_KE_prev_key1_reg_62_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_61_ ( .D(top_core_KE_n4858), .CK(n3894), .Q(top_core_KE_prev_key1_reg_61_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_60_ ( .D(top_core_KE_n4859), .CK(n3891), .Q(top_core_KE_prev_key1_reg_60_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_59_ ( .D(top_core_KE_n4860), .CK(n3904), .Q(top_core_KE_prev_key1_reg_59_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_58_ ( .D(top_core_KE_n4861), .CK(n3900), .Q(top_core_KE_prev_key1_reg_58_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_56_ ( .D(top_core_KE_n4863), .CK(n3898), .Q(top_core_KE_prev_key1_reg_56_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_121_ ( .D(top_core_KE_n4671), .CK(
        n3899), .Q(top_core_KE_prev_key0_reg_121_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_25_ ( .D(top_core_KE_n4766), .CK(n3899), .Q(top_core_KE_prev_key0_reg_25_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_15_ ( .D(top_core_KE_n4776), .CK(n3897), .Q(top_core_KE_prev_key0_reg_15_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_31_ ( .D(top_core_KE_n4760), .CK(n3902), .Q(top_core_KE_prev_key0_reg_31_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_22_ ( .D(top_core_KE_n4769), .CK(n3896), .Q(top_core_KE_prev_key0_reg_22_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_126_ ( .D(top_core_KE_n4666), .CK(
        n3896), .Q(top_core_KE_prev_key0_reg_126_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_30_ ( .D(top_core_KE_n4761), .CK(n3897), .Q(top_core_KE_prev_key0_reg_30_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_21_ ( .D(top_core_KE_n4770), .CK(n3894), .Q(top_core_KE_prev_key0_reg_21_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_125_ ( .D(top_core_KE_n4667), .CK(
        n3894), .Q(top_core_KE_prev_key0_reg_125_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_29_ ( .D(top_core_KE_n4762), .CK(n3893), .Q(top_core_KE_prev_key0_reg_29_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_20_ ( .D(top_core_KE_n4771), .CK(n3891), .Q(top_core_KE_prev_key0_reg_20_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_124_ ( .D(top_core_KE_n4668), .CK(
        n3892), .Q(top_core_KE_prev_key0_reg_124_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_28_ ( .D(top_core_KE_n4763), .CK(n3892), .Q(top_core_KE_prev_key0_reg_28_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_19_ ( .D(top_core_KE_n4772), .CK(n3904), .Q(top_core_KE_prev_key0_reg_19_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_123_ ( .D(top_core_KE_n4669), .CK(
        n3903), .Q(top_core_KE_prev_key0_reg_123_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_27_ ( .D(top_core_KE_n4764), .CK(n3903), .Q(top_core_KE_prev_key0_reg_27_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_18_ ( .D(top_core_KE_n4773), .CK(n3901), .Q(top_core_KE_prev_key0_reg_18_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_122_ ( .D(top_core_KE_n4670), .CK(
        n3900), .Q(top_core_KE_prev_key0_reg_122_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_26_ ( .D(top_core_KE_n4765), .CK(n3900), .Q(top_core_KE_prev_key0_reg_26_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_17_ ( .D(top_core_KE_n4774), .CK(n3897), .Q(top_core_KE_prev_key0_reg_17_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_16_ ( .D(top_core_KE_n4775), .CK(n3898), .Q(top_core_KE_prev_key0_reg_16_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_120_ ( .D(top_core_KE_n4672), .CK(
        n3898), .Q(top_core_KE_prev_key0_reg_120_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_24_ ( .D(top_core_KE_n4767), .CK(n3898), .Q(top_core_KE_prev_key0_reg_24_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_14_ ( .D(top_core_KE_n4777), .CK(n3899), .Q(top_core_KE_prev_key0_reg_14_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_13_ ( .D(top_core_KE_n4778), .CK(n3901), .Q(top_core_KE_prev_key0_reg_13_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_12_ ( .D(top_core_KE_n4779), .CK(n3903), .Q(top_core_KE_prev_key0_reg_12_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_11_ ( .D(top_core_KE_n4780), .CK(n3905), .Q(top_core_KE_prev_key0_reg_11_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_2_ ( .D(top_core_KE_n4789), .CK(n3906), 
        .Q(top_core_KE_prev_key0_reg_2_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_10_ ( .D(top_core_KE_n4781), .CK(n3891), .Q(top_core_KE_prev_key0_reg_10_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_1_ ( .D(top_core_KE_n4790), .CK(n3892), 
        .Q(top_core_KE_prev_key0_reg_1_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_0_ ( .D(top_core_KE_n4791), .CK(n3894), 
        .Q(top_core_KE_prev_key0_reg_0_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_23_ ( .D(top_core_KE_n4768), .CK(n3895), .Q(top_core_KE_prev_key0_reg_23_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_111_ ( .D(top_core_KE_n4681), .CK(
        n3897), .Q(top_core_KE_prev_key0_reg_111_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_103_ ( .D(top_core_KE_n4689), .CK(
        n3903), .Q(top_core_KE_prev_key0_reg_103_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_102_ ( .D(top_core_KE_n4690), .CK(
        n3905), .Q(top_core_KE_prev_key0_reg_102_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_6_ ( .D(top_core_KE_n4785), .CK(n3905), 
        .Q(top_core_KE_prev_key0_reg_6_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_110_ ( .D(top_core_KE_n4682), .CK(
        n3899), .Q(top_core_KE_prev_key0_reg_110_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_101_ ( .D(top_core_KE_n4691), .CK(
        n3900), .Q(top_core_KE_prev_key0_reg_101_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_5_ ( .D(top_core_KE_n4786), .CK(n3900), 
        .Q(top_core_KE_prev_key0_reg_5_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_109_ ( .D(top_core_KE_n4683), .CK(
        n3901), .Q(top_core_KE_prev_key0_reg_109_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_100_ ( .D(top_core_KE_n4692), .CK(
        n3902), .Q(top_core_KE_prev_key0_reg_100_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_4_ ( .D(top_core_KE_n4787), .CK(n3902), 
        .Q(top_core_KE_prev_key0_reg_4_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_108_ ( .D(top_core_KE_n4684), .CK(
        n3903), .Q(top_core_KE_prev_key0_reg_108_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_99_ ( .D(top_core_KE_n4693), .CK(n3904), .Q(top_core_KE_prev_key0_reg_99_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_3_ ( .D(top_core_KE_n4788), .CK(n3904), 
        .Q(top_core_KE_prev_key0_reg_3_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_107_ ( .D(top_core_KE_n4685), .CK(
        n3905), .Q(top_core_KE_prev_key0_reg_107_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_98_ ( .D(top_core_KE_n4920), .CK(n3906), .Q(top_core_KE_prev_key0_reg_98_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_106_ ( .D(top_core_KE_n4686), .CK(
        n3891), .Q(top_core_KE_prev_key0_reg_106_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_97_ ( .D(top_core_KE_n4694), .CK(n3892), .Q(top_core_KE_prev_key0_reg_97_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_105_ ( .D(top_core_KE_n4687), .CK(
        n3893), .Q(top_core_KE_prev_key0_reg_105_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_9_ ( .D(top_core_KE_n4782), .CK(n3893), 
        .Q(top_core_KE_prev_key0_reg_9_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_96_ ( .D(top_core_KE_n4695), .CK(n3893), .Q(top_core_KE_prev_key0_reg_96_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_104_ ( .D(top_core_KE_n4688), .CK(
        n3895), .Q(top_core_KE_prev_key0_reg_104_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_8_ ( .D(top_core_KE_n4783), .CK(n3895), 
        .Q(top_core_KE_prev_key0_reg_8_) );
  DFFHQX1 top_core_KE_prev_key0_reg_reg_7_ ( .D(top_core_KE_n4784), .CK(n3892), 
        .Q(top_core_KE_prev_key0_reg_7_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_121_ ( .D(top_core_KE_n4798), .CK(
        n3899), .Q(top_core_KE_prev_key1_reg_121_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_126_ ( .D(top_core_KE_n4793), .CK(
        n3896), .Q(top_core_KE_prev_key1_reg_126_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_125_ ( .D(top_core_KE_n4794), .CK(
        n3894), .Q(top_core_KE_prev_key1_reg_125_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_124_ ( .D(top_core_KE_n4795), .CK(
        n3892), .Q(top_core_KE_prev_key1_reg_124_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_123_ ( .D(top_core_KE_n4796), .CK(
        n3903), .Q(top_core_KE_prev_key1_reg_123_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_122_ ( .D(top_core_KE_n4797), .CK(
        n3900), .Q(top_core_KE_prev_key1_reg_122_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_120_ ( .D(top_core_KE_n4799), .CK(
        n3898), .Q(top_core_KE_prev_key1_reg_120_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_127_ ( .D(top_core_KE_n4792), .CK(
        n3902), .Q(top_core_KE_prev_key1_reg_127_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_21_ ( .D(top_core_KE_n4898), .CK(n3894), .Q(top_core_KE_prev_key1_reg_21_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_93_ ( .D(top_core_KE_n4826), .CK(n3894), .Q(top_core_KE_prev_key1_reg_93_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_29_ ( .D(top_core_KE_n4890), .CK(n3893), .Q(top_core_KE_prev_key1_reg_29_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_90_ ( .D(top_core_KE_n4829), .CK(n3900), .Q(top_core_KE_prev_key1_reg_90_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_5_ ( .D(top_core_KE_n4914), .CK(n3900), 
        .Q(top_core_KE_prev_key1_reg_5_) );
  DFFHQX1 top_core_KE_prev_key1_reg_reg_13_ ( .D(top_core_KE_n4906), .CK(n3901), .Q(top_core_KE_prev_key1_reg_13_) );
  DFFRHQX1 top_core_KE_rcon_reg_reg_3_ ( .D(top_core_KE_n4924), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_rcon_reg_3_) );
  DFFRHQX1 top_core_KE_rcon_reg_reg_2_ ( .D(top_core_KE_n4925), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_rcon_reg_2_) );
  DFFRHQX1 top_core_KE_rcon_reg_reg_0_ ( .D(top_core_KE_n4927), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_rcon_reg_0_) );
  DFFRHQX1 top_core_EC_rounds_reg_2_ ( .D(top_core_EC_n1297), .CK(n3721), .RN(
        n_RSTB), .Q(top_core_EC_rounds_2_) );
  DFFRHQX1 top_core_EC_rounds_reg_1_ ( .D(top_core_EC_n1296), .CK(n3721), .RN(
        n_RSTB), .Q(n7246) );
  DFFRHQX1 top_core_EC_rounds_reg_3_ ( .D(top_core_EC_n1298), .CK(n3721), .RN(
        n_RSTB), .Q(top_core_EC_rounds_3_) );
  DFFRHQX2 top_core_KE_rcon_reg_reg_7_ ( .D(top_core_KE_n4928), .CK(n3836), 
        .RN(n_RSTB), .Q(top_core_KE_rcon_reg_7_) );
  DFFRHQX2 top_core_EC_Core_Full_reg ( .D(top_core_EC_n1299), .CK(n3721), .RN(
        n_RSTB), .Q(top_core_Core_Full) );
  DFFHQX1 top_core_io_div_16_c_reg_2_ ( .D(top_core_io_div_16_N8), .CK(n_CLK), 
        .Q(top_core_io_div_16_c_2_) );
  JKFFX1 top_core_io_div_16_c_reg_0_ ( .J(1'b1), .K(1'b1), .CK(n_CLK), .QN(
        top_core_io_div_16_n5) );
  DFFHQX1 top_core_io_div_16_c_reg_1_ ( .D(top_core_io_div_16_N7), .CK(n_CLK), 
        .Q(top_core_io_div_16_c_1_) );
  DFFRHQX1 top_core_io_NK_reg_1_ ( .D(top_core_io_n665), .CK(n_CLK), .RN(
        n_RSTB), .Q(top_core_io_NK_1_) );
  DFFRHQX1 top_core_io_NK_reg_2_ ( .D(top_core_io_n666), .CK(n_CLK), .RN(
        n_RSTB), .Q(top_core_io_NK_2_) );
  DFFRHQX1 top_core_io_CORE_FULL_reg ( .D(top_core_Core_Full), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CORE_FULL) );
  DFFRHQX1 top_core_io_operation_reg ( .D(top_core_io_n663), .CK(n_CLK), .RN(
        n_RSTB), .Q(top_core_io_operation) );
  DFFRHQX1 top_core_io_OK_reg ( .D(top_core_io_n1182), .CK(n_CLK), .RN(n_RSTB), 
        .Q(n_OK) );
  DFFRHQX1 top_core_io_Data_reg_reg_29__0_ ( .D(n4535), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_29__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_29__1_ ( .D(n4536), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_29__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_29__2_ ( .D(n4537), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_29__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_29__3_ ( .D(n4538), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_29__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_29__4_ ( .D(n4539), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_29__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_29__5_ ( .D(n4540), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_29__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_29__6_ ( .D(n4541), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_29__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_29__7_ ( .D(n4542), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_29__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_25__0_ ( .D(n4567), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_25__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_25__1_ ( .D(n4568), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_25__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_25__2_ ( .D(n4569), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_25__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_25__3_ ( .D(n4570), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_25__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_25__4_ ( .D(n4571), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_25__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_25__5_ ( .D(n4572), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_25__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_25__6_ ( .D(n4573), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_25__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_25__7_ ( .D(n4574), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_25__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_21__0_ ( .D(n4599), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_21__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_21__1_ ( .D(n4600), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_21__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_21__2_ ( .D(n4601), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_21__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_21__3_ ( .D(n4602), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_21__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_21__4_ ( .D(n4603), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_21__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_21__5_ ( .D(n4604), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_21__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_21__6_ ( .D(n4605), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_21__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_21__7_ ( .D(n4606), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_21__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_17__0_ ( .D(n4631), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_17__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_17__1_ ( .D(n4632), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_17__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_17__2_ ( .D(n4633), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_17__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_17__3_ ( .D(n4634), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_17__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_17__4_ ( .D(n4635), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_17__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_17__5_ ( .D(n4636), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_17__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_17__6_ ( .D(n4637), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_17__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_17__7_ ( .D(n4638), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_17__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_31__0_ ( .D(n4519), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_31__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_31__1_ ( .D(n4520), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_31__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_31__2_ ( .D(n4521), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_31__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_31__3_ ( .D(n4522), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_31__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_31__4_ ( .D(n4523), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_31__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_31__5_ ( .D(n4524), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_31__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_31__6_ ( .D(n4525), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_31__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_31__7_ ( .D(n4526), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_31__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_27__0_ ( .D(n4551), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_27__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_27__1_ ( .D(n4552), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_27__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_27__2_ ( .D(n4553), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_27__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_27__3_ ( .D(n4554), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_27__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_27__4_ ( .D(n4555), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_27__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_27__5_ ( .D(n4556), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_27__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_27__6_ ( .D(n4557), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_27__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_27__7_ ( .D(n4558), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_27__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_23__0_ ( .D(n4583), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_23__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_23__1_ ( .D(n4584), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_23__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_23__2_ ( .D(n4585), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_23__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_23__3_ ( .D(n4586), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_23__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_23__4_ ( .D(n4587), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_23__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_23__5_ ( .D(n4588), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_23__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_23__6_ ( .D(n4589), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_23__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_23__7_ ( .D(n4590), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_23__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_19__0_ ( .D(n4615), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_19__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_19__1_ ( .D(n4616), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_19__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_19__2_ ( .D(n4617), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_19__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_19__3_ ( .D(n4618), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_19__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_19__4_ ( .D(n4619), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_19__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_19__5_ ( .D(n4620), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_19__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_19__6_ ( .D(n4621), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_19__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_19__7_ ( .D(n4622), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_19__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_28__0_ ( .D(n4543), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_28__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_28__1_ ( .D(n4544), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_28__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_28__2_ ( .D(n4545), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_28__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_28__3_ ( .D(n4546), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_28__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_28__4_ ( .D(n4547), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_28__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_28__5_ ( .D(n4548), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_28__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_28__6_ ( .D(n4549), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_28__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_28__7_ ( .D(n4550), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_28__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_24__0_ ( .D(n4575), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_24__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_24__1_ ( .D(n4576), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_24__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_24__2_ ( .D(n4577), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_24__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_24__3_ ( .D(n4578), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_24__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_24__4_ ( .D(n4579), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_24__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_24__5_ ( .D(n4580), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_24__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_24__6_ ( .D(n4581), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_24__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_24__7_ ( .D(n4582), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_24__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_20__0_ ( .D(n4607), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_20__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_20__1_ ( .D(n4608), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_20__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_20__2_ ( .D(n4609), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_20__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_20__3_ ( .D(n4610), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_20__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_20__4_ ( .D(n4611), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_20__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_20__5_ ( .D(n4612), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_20__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_20__6_ ( .D(n4613), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_20__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_20__7_ ( .D(n4614), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_20__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_16__0_ ( .D(n4639), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_16__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_16__1_ ( .D(n4640), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_16__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_16__2_ ( .D(n4641), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_16__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_16__3_ ( .D(n4642), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_16__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_16__4_ ( .D(n4643), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_16__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_16__5_ ( .D(n4644), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_16__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_16__6_ ( .D(n4645), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_16__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_16__7_ ( .D(n4646), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_16__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_30__0_ ( .D(n4527), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_30__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_30__1_ ( .D(n4528), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_30__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_30__2_ ( .D(n4529), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_30__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_30__3_ ( .D(n4530), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_30__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_30__4_ ( .D(n4531), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_30__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_30__5_ ( .D(n4532), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_30__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_30__6_ ( .D(n4533), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_30__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_30__7_ ( .D(n4534), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_30__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_26__0_ ( .D(n4559), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_26__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_26__1_ ( .D(n4560), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_26__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_26__2_ ( .D(n4561), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_26__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_26__3_ ( .D(n4562), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_26__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_26__4_ ( .D(n4563), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_26__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_26__5_ ( .D(n4564), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_26__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_26__6_ ( .D(n4565), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_26__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_26__7_ ( .D(n4566), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_26__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_22__0_ ( .D(n4591), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_22__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_22__1_ ( .D(n4592), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_22__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_22__2_ ( .D(n4593), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_22__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_22__3_ ( .D(n4594), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_22__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_22__4_ ( .D(n4595), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_22__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_22__5_ ( .D(n4596), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_22__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_22__6_ ( .D(n4597), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_22__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_22__7_ ( .D(n4598), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_22__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_18__0_ ( .D(n4623), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_18__0_) );
  DFFRHQX1 top_core_io_Data_reg_reg_18__1_ ( .D(n4624), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_18__1_) );
  DFFRHQX1 top_core_io_Data_reg_reg_18__2_ ( .D(n4625), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_18__2_) );
  DFFRHQX1 top_core_io_Data_reg_reg_18__3_ ( .D(n4626), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_18__3_) );
  DFFRHQX1 top_core_io_Data_reg_reg_18__4_ ( .D(n4627), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_18__4_) );
  DFFRHQX1 top_core_io_Data_reg_reg_18__5_ ( .D(n4628), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_18__5_) );
  DFFRHQX1 top_core_io_Data_reg_reg_18__6_ ( .D(n4629), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_18__6_) );
  DFFRHQX1 top_core_io_Data_reg_reg_18__7_ ( .D(n4630), .CK(n_CLK), .RN(n_RSTB), .Q(top_core_io_Data_reg_18__7_) );
  DFFRHQX1 top_core_io_Data_reg_reg_61__0_ ( .D(top_core_io_n683), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_232_) );
  DFFRHQX1 top_core_io_Data_reg_reg_61__1_ ( .D(top_core_io_n684), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_233_) );
  DFFRHQX1 top_core_io_Data_reg_reg_61__2_ ( .D(top_core_io_n685), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_234_) );
  DFFRHQX1 top_core_io_Data_reg_reg_61__3_ ( .D(top_core_io_n686), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_235_) );
  DFFRHQX1 top_core_io_Data_reg_reg_61__4_ ( .D(top_core_io_n687), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_236_) );
  DFFRHQX1 top_core_io_Data_reg_reg_61__5_ ( .D(top_core_io_n688), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_237_) );
  DFFRHQX1 top_core_io_Data_reg_reg_61__6_ ( .D(top_core_io_n689), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_238_) );
  DFFRHQX1 top_core_io_Data_reg_reg_61__7_ ( .D(top_core_io_n690), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_239_) );
  DFFRHQX1 top_core_io_Data_reg_reg_57__0_ ( .D(top_core_io_n715), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_200_) );
  DFFRHQX1 top_core_io_Data_reg_reg_57__1_ ( .D(top_core_io_n716), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_201_) );
  DFFRHQX1 top_core_io_Data_reg_reg_57__2_ ( .D(top_core_io_n717), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_202_) );
  DFFRHQX1 top_core_io_Data_reg_reg_57__3_ ( .D(top_core_io_n718), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_203_) );
  DFFRHQX1 top_core_io_Data_reg_reg_57__4_ ( .D(top_core_io_n719), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_204_) );
  DFFRHQX1 top_core_io_Data_reg_reg_57__5_ ( .D(top_core_io_n720), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_205_) );
  DFFRHQX1 top_core_io_Data_reg_reg_57__6_ ( .D(top_core_io_n721), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_206_) );
  DFFRHQX1 top_core_io_Data_reg_reg_57__7_ ( .D(top_core_io_n722), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_207_) );
  DFFRHQX1 top_core_io_Data_reg_reg_45__0_ ( .D(top_core_io_n811), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_104_) );
  DFFRHQX1 top_core_io_Data_reg_reg_45__1_ ( .D(top_core_io_n812), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_105_) );
  DFFRHQX1 top_core_io_Data_reg_reg_45__2_ ( .D(top_core_io_n813), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_106_) );
  DFFRHQX1 top_core_io_Data_reg_reg_45__3_ ( .D(top_core_io_n814), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_107_) );
  DFFRHQX1 top_core_io_Data_reg_reg_45__4_ ( .D(top_core_io_n815), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_108_) );
  DFFRHQX1 top_core_io_Data_reg_reg_45__5_ ( .D(top_core_io_n816), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_109_) );
  DFFRHQX1 top_core_io_Data_reg_reg_45__6_ ( .D(top_core_io_n817), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_110_) );
  DFFRHQX1 top_core_io_Data_reg_reg_45__7_ ( .D(top_core_io_n818), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_111_) );
  DFFRHQX1 top_core_io_Data_reg_reg_41__0_ ( .D(top_core_io_n843), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_72_) );
  DFFRHQX1 top_core_io_Data_reg_reg_41__1_ ( .D(top_core_io_n844), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_73_) );
  DFFRHQX1 top_core_io_Data_reg_reg_41__2_ ( .D(top_core_io_n845), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_74_) );
  DFFRHQX1 top_core_io_Data_reg_reg_41__3_ ( .D(top_core_io_n846), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_75_) );
  DFFRHQX1 top_core_io_Data_reg_reg_41__4_ ( .D(top_core_io_n847), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_76_) );
  DFFRHQX1 top_core_io_Data_reg_reg_41__5_ ( .D(top_core_io_n848), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_77_) );
  DFFRHQX1 top_core_io_Data_reg_reg_41__6_ ( .D(top_core_io_n849), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_78_) );
  DFFRHQX1 top_core_io_Data_reg_reg_41__7_ ( .D(top_core_io_n850), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_79_) );
  DFFRHQX1 top_core_io_Data_reg_reg_13__0_ ( .D(top_core_io_n1067), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_104_) );
  DFFRHQX1 top_core_io_Data_reg_reg_13__1_ ( .D(top_core_io_n1068), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_105_) );
  DFFRHQX1 top_core_io_Data_reg_reg_13__2_ ( .D(top_core_io_n1069), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_106_) );
  DFFRHQX1 top_core_io_Data_reg_reg_13__3_ ( .D(top_core_io_n1070), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_107_) );
  DFFRHQX1 top_core_io_Data_reg_reg_13__4_ ( .D(top_core_io_n1071), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_108_) );
  DFFRHQX1 top_core_io_Data_reg_reg_13__5_ ( .D(top_core_io_n1072), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_109_) );
  DFFRHQX1 top_core_io_Data_reg_reg_13__6_ ( .D(top_core_io_n1073), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_110_) );
  DFFRHQX1 top_core_io_Data_reg_reg_13__7_ ( .D(top_core_io_n1074), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_111_) );
  DFFRHQX1 top_core_io_Data_reg_reg_9__0_ ( .D(top_core_io_n1099), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_72_) );
  DFFRHQX1 top_core_io_Data_reg_reg_9__1_ ( .D(top_core_io_n1100), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_73_) );
  DFFRHQX1 top_core_io_Data_reg_reg_9__2_ ( .D(top_core_io_n1101), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_74_) );
  DFFRHQX1 top_core_io_Data_reg_reg_9__3_ ( .D(top_core_io_n1102), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_75_) );
  DFFRHQX1 top_core_io_Data_reg_reg_9__4_ ( .D(top_core_io_n1103), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_76_) );
  DFFRHQX1 top_core_io_Data_reg_reg_9__5_ ( .D(top_core_io_n1104), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_77_) );
  DFFRHQX1 top_core_io_Data_reg_reg_9__6_ ( .D(top_core_io_n1105), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_78_) );
  DFFRHQX1 top_core_io_Data_reg_reg_9__7_ ( .D(top_core_io_n1106), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_79_) );
  DFFRHQX1 top_core_io_Data_reg_reg_63__0_ ( .D(top_core_io_n667), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_248_) );
  DFFRHQX1 top_core_io_Data_reg_reg_63__1_ ( .D(top_core_io_n668), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_249_) );
  DFFRHQX1 top_core_io_Data_reg_reg_63__2_ ( .D(top_core_io_n669), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_250_) );
  DFFRHQX1 top_core_io_Data_reg_reg_63__3_ ( .D(top_core_io_n670), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_251_) );
  DFFRHQX1 top_core_io_Data_reg_reg_63__4_ ( .D(top_core_io_n671), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_252_) );
  DFFRHQX1 top_core_io_Data_reg_reg_63__5_ ( .D(top_core_io_n672), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_253_) );
  DFFRHQX1 top_core_io_Data_reg_reg_63__6_ ( .D(top_core_io_n673), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_254_) );
  DFFRHQX1 top_core_io_Data_reg_reg_63__7_ ( .D(top_core_io_n674), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_255_) );
  DFFRHQX1 top_core_io_Data_reg_reg_59__0_ ( .D(top_core_io_n699), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_216_) );
  DFFRHQX1 top_core_io_Data_reg_reg_59__1_ ( .D(top_core_io_n700), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_217_) );
  DFFRHQX1 top_core_io_Data_reg_reg_59__2_ ( .D(top_core_io_n701), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_218_) );
  DFFRHQX1 top_core_io_Data_reg_reg_59__3_ ( .D(top_core_io_n702), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_219_) );
  DFFRHQX1 top_core_io_Data_reg_reg_59__4_ ( .D(top_core_io_n703), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_220_) );
  DFFRHQX1 top_core_io_Data_reg_reg_59__5_ ( .D(top_core_io_n704), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_221_) );
  DFFRHQX1 top_core_io_Data_reg_reg_59__6_ ( .D(top_core_io_n705), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_222_) );
  DFFRHQX1 top_core_io_Data_reg_reg_59__7_ ( .D(top_core_io_n706), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_223_) );
  DFFRHQX1 top_core_io_Data_reg_reg_47__0_ ( .D(top_core_io_n795), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_120_) );
  DFFRHQX1 top_core_io_Data_reg_reg_47__1_ ( .D(top_core_io_n796), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_121_) );
  DFFRHQX1 top_core_io_Data_reg_reg_47__2_ ( .D(top_core_io_n797), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_122_) );
  DFFRHQX1 top_core_io_Data_reg_reg_47__3_ ( .D(top_core_io_n798), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_123_) );
  DFFRHQX1 top_core_io_Data_reg_reg_47__4_ ( .D(top_core_io_n799), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_124_) );
  DFFRHQX1 top_core_io_Data_reg_reg_47__5_ ( .D(top_core_io_n800), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_125_) );
  DFFRHQX1 top_core_io_Data_reg_reg_47__6_ ( .D(top_core_io_n801), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_126_) );
  DFFRHQX1 top_core_io_Data_reg_reg_47__7_ ( .D(top_core_io_n802), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_127_) );
  DFFRHQX1 top_core_io_Data_reg_reg_43__0_ ( .D(top_core_io_n827), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_88_) );
  DFFRHQX1 top_core_io_Data_reg_reg_43__1_ ( .D(top_core_io_n828), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_89_) );
  DFFRHQX1 top_core_io_Data_reg_reg_43__2_ ( .D(top_core_io_n829), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_90_) );
  DFFRHQX1 top_core_io_Data_reg_reg_43__3_ ( .D(top_core_io_n830), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_91_) );
  DFFRHQX1 top_core_io_Data_reg_reg_43__4_ ( .D(top_core_io_n831), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_92_) );
  DFFRHQX1 top_core_io_Data_reg_reg_43__5_ ( .D(top_core_io_n832), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_93_) );
  DFFRHQX1 top_core_io_Data_reg_reg_43__6_ ( .D(top_core_io_n833), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_94_) );
  DFFRHQX1 top_core_io_Data_reg_reg_43__7_ ( .D(top_core_io_n834), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_95_) );
  DFFRHQX1 top_core_io_Data_reg_reg_15__0_ ( .D(top_core_io_n1051), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_120_) );
  DFFRHQX1 top_core_io_Data_reg_reg_15__1_ ( .D(top_core_io_n1052), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_121_) );
  DFFRHQX1 top_core_io_Data_reg_reg_15__2_ ( .D(top_core_io_n1053), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_122_) );
  DFFRHQX1 top_core_io_Data_reg_reg_15__3_ ( .D(top_core_io_n1054), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_123_) );
  DFFRHQX1 top_core_io_Data_reg_reg_15__4_ ( .D(top_core_io_n1055), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_124_) );
  DFFRHQX1 top_core_io_Data_reg_reg_15__5_ ( .D(top_core_io_n1056), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_125_) );
  DFFRHQX1 top_core_io_Data_reg_reg_15__6_ ( .D(top_core_io_n1057), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_126_) );
  DFFRHQX1 top_core_io_Data_reg_reg_15__7_ ( .D(top_core_io_n1058), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_127_) );
  DFFRHQX1 top_core_io_Data_reg_reg_11__0_ ( .D(top_core_io_n1083), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_88_) );
  DFFRHQX1 top_core_io_Data_reg_reg_11__1_ ( .D(top_core_io_n1084), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_89_) );
  DFFRHQX1 top_core_io_Data_reg_reg_11__2_ ( .D(top_core_io_n1085), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_90_) );
  DFFRHQX1 top_core_io_Data_reg_reg_11__3_ ( .D(top_core_io_n1086), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_91_) );
  DFFRHQX1 top_core_io_Data_reg_reg_11__4_ ( .D(top_core_io_n1087), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_92_) );
  DFFRHQX1 top_core_io_Data_reg_reg_11__5_ ( .D(top_core_io_n1088), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_93_) );
  DFFRHQX1 top_core_io_Data_reg_reg_11__6_ ( .D(top_core_io_n1089), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_94_) );
  DFFRHQX1 top_core_io_Data_reg_reg_11__7_ ( .D(top_core_io_n1090), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_95_) );
  DFFRHQX1 top_core_io_Data_reg_reg_60__0_ ( .D(top_core_io_n691), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_224_) );
  DFFRHQX1 top_core_io_Data_reg_reg_60__1_ ( .D(top_core_io_n692), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_225_) );
  DFFRHQX1 top_core_io_Data_reg_reg_60__2_ ( .D(top_core_io_n693), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_226_) );
  DFFRHQX1 top_core_io_Data_reg_reg_60__3_ ( .D(top_core_io_n694), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_227_) );
  DFFRHQX1 top_core_io_Data_reg_reg_60__4_ ( .D(top_core_io_n695), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_228_) );
  DFFRHQX1 top_core_io_Data_reg_reg_60__5_ ( .D(top_core_io_n696), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_229_) );
  DFFRHQX1 top_core_io_Data_reg_reg_60__6_ ( .D(top_core_io_n697), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_230_) );
  DFFRHQX1 top_core_io_Data_reg_reg_60__7_ ( .D(top_core_io_n698), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_231_) );
  DFFRHQX1 top_core_io_Data_reg_reg_44__0_ ( .D(top_core_io_n819), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_96_) );
  DFFRHQX1 top_core_io_Data_reg_reg_44__1_ ( .D(top_core_io_n820), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_97_) );
  DFFRHQX1 top_core_io_Data_reg_reg_44__2_ ( .D(top_core_io_n821), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_98_) );
  DFFRHQX1 top_core_io_Data_reg_reg_44__3_ ( .D(top_core_io_n822), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_99_) );
  DFFRHQX1 top_core_io_Data_reg_reg_44__4_ ( .D(top_core_io_n823), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_100_) );
  DFFRHQX1 top_core_io_Data_reg_reg_44__5_ ( .D(top_core_io_n824), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_101_) );
  DFFRHQX1 top_core_io_Data_reg_reg_44__6_ ( .D(top_core_io_n825), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_102_) );
  DFFRHQX1 top_core_io_Data_reg_reg_44__7_ ( .D(top_core_io_n826), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_103_) );
  DFFRHQX1 top_core_io_Data_reg_reg_12__0_ ( .D(top_core_io_n1075), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_96_) );
  DFFRHQX1 top_core_io_Data_reg_reg_12__1_ ( .D(top_core_io_n1076), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_97_) );
  DFFRHQX1 top_core_io_Data_reg_reg_12__2_ ( .D(top_core_io_n1077), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_98_) );
  DFFRHQX1 top_core_io_Data_reg_reg_12__3_ ( .D(top_core_io_n1078), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_99_) );
  DFFRHQX1 top_core_io_Data_reg_reg_12__4_ ( .D(top_core_io_n1079), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_100_) );
  DFFRHQX1 top_core_io_Data_reg_reg_12__5_ ( .D(top_core_io_n1080), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_101_) );
  DFFRHQX1 top_core_io_Data_reg_reg_12__6_ ( .D(top_core_io_n1081), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_102_) );
  DFFRHQX1 top_core_io_Data_reg_reg_12__7_ ( .D(top_core_io_n1082), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_103_) );
  DFFRHQX1 top_core_io_Data_reg_reg_62__0_ ( .D(top_core_io_n675), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_240_) );
  DFFRHQX1 top_core_io_Data_reg_reg_62__1_ ( .D(top_core_io_n676), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_241_) );
  DFFRHQX1 top_core_io_Data_reg_reg_62__2_ ( .D(top_core_io_n677), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_242_) );
  DFFRHQX1 top_core_io_Data_reg_reg_62__3_ ( .D(top_core_io_n678), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_243_) );
  DFFRHQX1 top_core_io_Data_reg_reg_62__4_ ( .D(top_core_io_n679), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_244_) );
  DFFRHQX1 top_core_io_Data_reg_reg_62__5_ ( .D(top_core_io_n680), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_245_) );
  DFFRHQX1 top_core_io_Data_reg_reg_62__6_ ( .D(top_core_io_n681), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_246_) );
  DFFRHQX1 top_core_io_Data_reg_reg_62__7_ ( .D(top_core_io_n682), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_247_) );
  DFFRHQX1 top_core_io_Data_reg_reg_58__0_ ( .D(top_core_io_n707), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_208_) );
  DFFRHQX1 top_core_io_Data_reg_reg_58__1_ ( .D(top_core_io_n708), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_209_) );
  DFFRHQX1 top_core_io_Data_reg_reg_58__2_ ( .D(top_core_io_n709), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_210_) );
  DFFRHQX1 top_core_io_Data_reg_reg_58__3_ ( .D(top_core_io_n710), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_211_) );
  DFFRHQX1 top_core_io_Data_reg_reg_58__4_ ( .D(top_core_io_n711), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_212_) );
  DFFRHQX1 top_core_io_Data_reg_reg_58__5_ ( .D(top_core_io_n712), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_213_) );
  DFFRHQX1 top_core_io_Data_reg_reg_58__6_ ( .D(top_core_io_n713), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_214_) );
  DFFRHQX1 top_core_io_Data_reg_reg_58__7_ ( .D(top_core_io_n714), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_215_) );
  DFFRHQX1 top_core_io_Data_reg_reg_46__0_ ( .D(top_core_io_n803), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_112_) );
  DFFRHQX1 top_core_io_Data_reg_reg_46__1_ ( .D(top_core_io_n804), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_113_) );
  DFFRHQX1 top_core_io_Data_reg_reg_46__2_ ( .D(top_core_io_n805), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_114_) );
  DFFRHQX1 top_core_io_Data_reg_reg_46__3_ ( .D(top_core_io_n806), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_115_) );
  DFFRHQX1 top_core_io_Data_reg_reg_46__4_ ( .D(top_core_io_n807), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_116_) );
  DFFRHQX1 top_core_io_Data_reg_reg_46__5_ ( .D(top_core_io_n808), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_117_) );
  DFFRHQX1 top_core_io_Data_reg_reg_46__6_ ( .D(top_core_io_n809), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_118_) );
  DFFRHQX1 top_core_io_Data_reg_reg_46__7_ ( .D(top_core_io_n810), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_119_) );
  DFFRHQX1 top_core_io_Data_reg_reg_42__0_ ( .D(top_core_io_n835), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_80_) );
  DFFRHQX1 top_core_io_Data_reg_reg_42__1_ ( .D(top_core_io_n836), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_81_) );
  DFFRHQX1 top_core_io_Data_reg_reg_42__2_ ( .D(top_core_io_n837), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_82_) );
  DFFRHQX1 top_core_io_Data_reg_reg_42__3_ ( .D(top_core_io_n838), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_83_) );
  DFFRHQX1 top_core_io_Data_reg_reg_42__4_ ( .D(top_core_io_n839), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_84_) );
  DFFRHQX1 top_core_io_Data_reg_reg_42__5_ ( .D(top_core_io_n840), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_85_) );
  DFFRHQX1 top_core_io_Data_reg_reg_42__6_ ( .D(top_core_io_n841), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_86_) );
  DFFRHQX1 top_core_io_Data_reg_reg_42__7_ ( .D(top_core_io_n842), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_87_) );
  DFFRHQX1 top_core_io_Data_reg_reg_14__0_ ( .D(top_core_io_n1059), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_112_) );
  DFFRHQX1 top_core_io_Data_reg_reg_14__1_ ( .D(top_core_io_n1060), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_113_) );
  DFFRHQX1 top_core_io_Data_reg_reg_14__2_ ( .D(top_core_io_n1061), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_114_) );
  DFFRHQX1 top_core_io_Data_reg_reg_14__3_ ( .D(top_core_io_n1062), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_115_) );
  DFFRHQX1 top_core_io_Data_reg_reg_14__4_ ( .D(top_core_io_n1063), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_116_) );
  DFFRHQX1 top_core_io_Data_reg_reg_14__5_ ( .D(top_core_io_n1064), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_117_) );
  DFFRHQX1 top_core_io_Data_reg_reg_14__6_ ( .D(top_core_io_n1065), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_118_) );
  DFFRHQX1 top_core_io_Data_reg_reg_14__7_ ( .D(top_core_io_n1066), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_119_) );
  DFFRHQX1 top_core_io_Data_reg_reg_10__0_ ( .D(top_core_io_n1091), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_80_) );
  DFFRHQX1 top_core_io_Data_reg_reg_10__1_ ( .D(top_core_io_n1092), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_81_) );
  DFFRHQX1 top_core_io_Data_reg_reg_10__2_ ( .D(top_core_io_n1093), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_82_) );
  DFFRHQX1 top_core_io_Data_reg_reg_10__3_ ( .D(top_core_io_n1094), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_83_) );
  DFFRHQX1 top_core_io_Data_reg_reg_10__4_ ( .D(top_core_io_n1095), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_84_) );
  DFFRHQX1 top_core_io_Data_reg_reg_10__5_ ( .D(top_core_io_n1096), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_85_) );
  DFFRHQX1 top_core_io_Data_reg_reg_10__6_ ( .D(top_core_io_n1097), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_86_) );
  DFFRHQX1 top_core_io_Data_reg_reg_10__7_ ( .D(top_core_io_n1098), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_87_) );
  DFFHQX1 top_core_io_div_16_clk_slow_reg ( .D(top_core_io_div_16_n3), .CK(
        n_CLK), .Q(top_core_clk_slow) );
  AND2X2 top_core_KE_U5608 ( .A(top_core_KE_key_mem_14__103_), .B(n4078), .Y(
        top_core_KE_n5553) );
  AND2X2 top_core_KE_U5160 ( .A(top_core_KE_key_mem_14__39_), .B(n4080), .Y(
        top_core_KE_n5169) );
  AND2X2 top_core_KE_U5440 ( .A(top_core_KE_key_mem_14__79_), .B(n4073), .Y(
        top_core_KE_n5409) );
  AND2X2 top_core_KE_U5272 ( .A(top_core_KE_key_mem_14__55_), .B(n4067), .Y(
        top_core_KE_n5265) );
  AND2X2 top_core_KE_U5720 ( .A(top_core_KE_key_mem_14__119_), .B(n4114), .Y(
        top_core_KE_n5649) );
  AND2X2 top_core_KE_U5104 ( .A(top_core_KE_key_mem_14__31_), .B(n4095), .Y(
        top_core_KE_n5121) );
  AND2X2 top_core_KE_U4936 ( .A(top_core_KE_key_mem_14__7_), .B(n4092), .Y(
        top_core_KE_n4977) );
  AND2X2 top_core_KE_U5384 ( .A(top_core_KE_key_mem_14__71_), .B(n4076), .Y(
        top_core_KE_n5361) );
  AND2X2 top_core_KE_U5664 ( .A(top_core_KE_key_mem_14__111_), .B(n4092), .Y(
        top_core_KE_n5601) );
  AND2X2 top_core_KE_U5496 ( .A(top_core_KE_key_mem_14__87_), .B(n4074), .Y(
        top_core_KE_n5457) );
  AND2X2 top_core_KE_U5048 ( .A(top_core_KE_key_mem_14__23_), .B(n4084), .Y(
        top_core_KE_n5073) );
  AND2X2 top_core_KE_U5328 ( .A(top_core_KE_key_mem_14__63_), .B(n4080), .Y(
        top_core_KE_n5313) );
  AND2X2 top_core_KE_U5552 ( .A(top_core_KE_key_mem_14__95_), .B(n4070), .Y(
        top_core_KE_n5505) );
  AND2X2 top_core_KE_U4992 ( .A(top_core_KE_key_mem_14__15_), .B(n4088), .Y(
        top_core_KE_n5025) );
  AND2X2 top_core_KE_U5216 ( .A(top_core_KE_key_mem_14__47_), .B(n4083), .Y(
        top_core_KE_n5217) );
  AND2X2 top_core_KE_U5776 ( .A(top_core_KE_key_mem_14__127_), .B(n4079), .Y(
        top_core_KE_n5697) );
  AND2X2 top_core_KE_U5783 ( .A(top_core_KE_key_mem_14__128_), .B(n4093), .Y(
        top_core_KE_n5703) );
  AND2X2 top_core_KE_U5132 ( .A(top_core_KE_key_mem_14__35_), .B(n4034), .Y(
        top_core_KE_n5145) );
  AND2X2 top_core_KE_U5412 ( .A(top_core_KE_key_mem_14__75_), .B(n4088), .Y(
        top_core_KE_n5385) );
  AND2X2 top_core_KE_U5692 ( .A(top_core_KE_key_mem_14__115_), .B(n4067), .Y(
        top_core_KE_n5625) );
  AND2X2 top_core_KE_U5076 ( .A(top_core_KE_key_mem_14__27_), .B(n4083), .Y(
        top_core_KE_n5097) );
  AND2X2 top_core_KE_U5356 ( .A(top_core_KE_key_mem_14__67_), .B(n4078), .Y(
        top_core_KE_n5337) );
  AND2X2 top_core_KE_U5636 ( .A(top_core_KE_key_mem_14__107_), .B(n4091), .Y(
        top_core_KE_n5577) );
  AND2X2 top_core_KE_U5020 ( .A(top_core_KE_key_mem_14__19_), .B(n4086), .Y(
        top_core_KE_n5049) );
  AND2X2 top_core_KE_U5300 ( .A(top_core_KE_key_mem_14__59_), .B(n4115), .Y(
        top_core_KE_n5289) );
  AND2X2 top_core_KE_U5580 ( .A(top_core_KE_key_mem_14__99_), .B(n4081), .Y(
        top_core_KE_n5529) );
  AND2X2 top_core_KE_U4908 ( .A(top_core_KE_key_mem_14__3_), .B(n4094), .Y(
        top_core_KE_n4953) );
  AND2X2 top_core_KE_U5244 ( .A(top_core_KE_key_mem_14__51_), .B(n4082), .Y(
        top_core_KE_n5241) );
  AND2X2 top_core_KE_U5468 ( .A(top_core_KE_key_mem_14__83_), .B(n4087), .Y(
        top_core_KE_n5433) );
  AND2X2 top_core_KE_U5601 ( .A(top_core_KE_key_mem_14__102_), .B(n4069), .Y(
        top_core_KE_n5547) );
  AND2X2 top_core_KE_U5153 ( .A(top_core_KE_key_mem_14__38_), .B(n4081), .Y(
        top_core_KE_n5163) );
  AND2X2 top_core_KE_U5433 ( .A(top_core_KE_key_mem_14__78_), .B(n4113), .Y(
        top_core_KE_n5403) );
  AND2X2 top_core_KE_U5097 ( .A(top_core_KE_key_mem_14__30_), .B(n4111), .Y(
        top_core_KE_n5115) );
  AND2X2 top_core_KE_U5657 ( .A(top_core_KE_key_mem_14__110_), .B(n4075), .Y(
        top_core_KE_n5595) );
  AND2X2 top_core_KE_U5321 ( .A(top_core_KE_key_mem_14__62_), .B(n4080), .Y(
        top_core_KE_n5307) );
  AND2X2 top_core_KE_U5524 ( .A(top_core_KE_key_mem_14__91_), .B(n4072), .Y(
        top_core_KE_n5481) );
  AND2X2 top_core_KE_U4964 ( .A(top_core_KE_key_mem_14__11_), .B(n4090), .Y(
        top_core_KE_n5001) );
  AND2X2 top_core_KE_U5713 ( .A(top_core_KE_key_mem_14__118_), .B(n4068), .Y(
        top_core_KE_n5643) );
  AND2X2 top_core_KE_U4929 ( .A(top_core_KE_key_mem_14__6_), .B(n4092), .Y(
        top_core_KE_n4971) );
  AND2X2 top_core_KE_U5377 ( .A(top_core_KE_key_mem_14__70_), .B(n4076), .Y(
        top_core_KE_n5355) );
  AND2X2 top_core_KE_U5748 ( .A(top_core_KE_key_mem_14__123_), .B(n4070), .Y(
        top_core_KE_n5673) );
  AND2X2 top_core_KE_U5188 ( .A(top_core_KE_key_mem_14__43_), .B(n4070), .Y(
        top_core_KE_n5193) );
  AND2X2 top_core_KE_U5041 ( .A(top_core_KE_key_mem_14__22_), .B(n4084), .Y(
        top_core_KE_n5067) );
  AND2X2 top_core_KE_U5265 ( .A(top_core_KE_key_mem_14__54_), .B(n4068), .Y(
        top_core_KE_n5259) );
  AND2X2 top_core_KE_U5699 ( .A(top_core_KE_key_mem_14__116_), .B(n4066), .Y(
        top_core_KE_n5631) );
  AND2X2 top_core_KE_U5146 ( .A(top_core_KE_key_mem_14__37_), .B(n4076), .Y(
        top_core_KE_n5157) );
  AND2X2 top_core_KE_U5587 ( .A(top_core_KE_key_mem_14__100_), .B(n4086), .Y(
        top_core_KE_n5535) );
  AND2X2 top_core_KE_U5594 ( .A(top_core_KE_key_mem_14__101_), .B(n4088), .Y(
        top_core_KE_n5541) );
  AND2X2 top_core_KE_U5363 ( .A(top_core_KE_key_mem_14__68_), .B(n4077), .Y(
        top_core_KE_n5343) );
  AND2X2 top_core_KE_U5489 ( .A(top_core_KE_key_mem_14__86_), .B(n4074), .Y(
        top_core_KE_n5451) );
  AND2X2 top_core_KE_U5139 ( .A(top_core_KE_key_mem_14__36_), .B(n4077), .Y(
        top_core_KE_n5151) );
  AND2X2 top_core_KE_U5426 ( .A(top_core_KE_key_mem_14__77_), .B(n4070), .Y(
        top_core_KE_n5397) );
  AND2X2 top_core_KE_U5419 ( .A(top_core_KE_key_mem_14__76_), .B(n4071), .Y(
        top_core_KE_n5391) );
  AND2X2 top_core_KE_U5090 ( .A(top_core_KE_key_mem_14__29_), .B(n4087), .Y(
        top_core_KE_n5109) );
  AND2X2 top_core_KE_U5083 ( .A(top_core_KE_key_mem_14__28_), .B(n4090), .Y(
        top_core_KE_n5103) );
  AND2X2 top_core_KE_U5650 ( .A(top_core_KE_key_mem_14__109_), .B(n4069), .Y(
        top_core_KE_n5589) );
  AND2X2 top_core_KE_U5643 ( .A(top_core_KE_key_mem_14__108_), .B(n4069), .Y(
        top_core_KE_n5583) );
  AND2X2 top_core_KE_U5314 ( .A(top_core_KE_key_mem_14__61_), .B(n4081), .Y(
        top_core_KE_n5301) );
  AND2X2 top_core_KE_U5307 ( .A(top_core_KE_key_mem_14__60_), .B(n4081), .Y(
        top_core_KE_n5295) );
  AND2X2 top_core_KE_U5545 ( .A(top_core_KE_key_mem_14__94_), .B(n4070), .Y(
        top_core_KE_n5499) );
  AND2X2 top_core_KE_U4985 ( .A(top_core_KE_key_mem_14__14_), .B(n4088), .Y(
        top_core_KE_n5019) );
  AND2X2 top_core_KE_U5706 ( .A(top_core_KE_key_mem_14__117_), .B(n4066), .Y(
        top_core_KE_n5637) );
  AND2X2 top_core_KE_U5370 ( .A(top_core_KE_key_mem_14__69_), .B(n4077), .Y(
        top_core_KE_n5349) );
  AND2X2 top_core_KE_U5209 ( .A(top_core_KE_key_mem_14__46_), .B(n4113), .Y(
        top_core_KE_n5211) );
  AND2X2 top_core_KE_U5027 ( .A(top_core_KE_key_mem_14__20_), .B(n4085), .Y(
        top_core_KE_n5055) );
  AND2X2 top_core_KE_U5034 ( .A(top_core_KE_key_mem_14__21_), .B(n4085), .Y(
        top_core_KE_n5061) );
  AND2X2 top_core_KE_U4922 ( .A(top_core_KE_key_mem_14__5_), .B(n4093), .Y(
        top_core_KE_n4965) );
  AND2X2 top_core_KE_U5251 ( .A(top_core_KE_key_mem_14__52_), .B(n4078), .Y(
        top_core_KE_n5247) );
  AND2X2 top_core_KE_U5258 ( .A(top_core_KE_key_mem_14__53_), .B(n4067), .Y(
        top_core_KE_n5253) );
  AND2X2 top_core_KE_U4915 ( .A(top_core_KE_key_mem_14__4_), .B(n4093), .Y(
        top_core_KE_n4959) );
  AND2X2 top_core_KE_U5769 ( .A(top_core_KE_key_mem_14__126_), .B(n4111), .Y(
        top_core_KE_n5691) );
  AND2X2 top_core_KE_U5685 ( .A(top_core_KE_key_mem_14__114_), .B(n4067), .Y(
        top_core_KE_n5619) );
  AND2X2 top_core_KE_U5349 ( .A(top_core_KE_key_mem_14__66_), .B(n4078), .Y(
        top_core_KE_n5331) );
  AND2X2 top_core_KE_U5475 ( .A(top_core_KE_key_mem_14__84_), .B(n4075), .Y(
        top_core_KE_n5439) );
  AND2X2 top_core_KE_U5482 ( .A(top_core_KE_key_mem_14__85_), .B(n4075), .Y(
        top_core_KE_n5445) );
  AND2X2 top_core_KE_U5013 ( .A(top_core_KE_key_mem_14__18_), .B(n4086), .Y(
        top_core_KE_n5043) );
  AND2X2 top_core_KE_U5111 ( .A(top_core_KE_key_mem_14__32_), .B(n4082), .Y(
        top_core_KE_n5127) );
  AND2X2 top_core_KE_U5391 ( .A(top_core_KE_key_mem_14__72_), .B(n4069), .Y(
        top_core_KE_n5367) );
  AND2X2 top_core_KE_U5055 ( .A(top_core_KE_key_mem_14__24_), .B(n4077), .Y(
        top_core_KE_n5079) );
  AND2X2 top_core_KE_U5615 ( .A(top_core_KE_key_mem_14__104_), .B(n4085), .Y(
        top_core_KE_n5559) );
  AND2X2 top_core_KE_U5279 ( .A(top_core_KE_key_mem_14__56_), .B(n4082), .Y(
        top_core_KE_n5271) );
  AND2X2 top_core_KE_U5559 ( .A(top_core_KE_key_mem_14__96_), .B(n4111), .Y(
        top_core_KE_n5511) );
  AND2X2 top_core_KE_U5531 ( .A(top_core_KE_key_mem_14__92_), .B(n4071), .Y(
        top_core_KE_n5487) );
  AND2X2 top_core_KE_U5538 ( .A(top_core_KE_key_mem_14__93_), .B(n4071), .Y(
        top_core_KE_n5493) );
  AND2X2 top_core_KE_U4971 ( .A(top_core_KE_key_mem_14__12_), .B(n4089), .Y(
        top_core_KE_n5007) );
  AND2X2 top_core_KE_U4978 ( .A(top_core_KE_key_mem_14__13_), .B(n4089), .Y(
        top_core_KE_n5013) );
  AND2X2 top_core_KE_U5230 ( .A(top_core_KE_key_mem_14__49_), .B(n4084), .Y(
        top_core_KE_n5229) );
  AND2X2 top_core_KE_U5223 ( .A(top_core_KE_key_mem_14__48_), .B(n4083), .Y(
        top_core_KE_n5223) );
  AND2X2 top_core_KE_U5671 ( .A(top_core_KE_key_mem_14__112_), .B(n4068), .Y(
        top_core_KE_n5607) );
  AND2X2 top_core_KE_U4887 ( .A(top_core_KE_key_mem_14__0_), .B(n4095), .Y(
        top_core_KE_n4935) );
  AND2X2 top_core_KE_U5755 ( .A(top_core_KE_key_mem_14__124_), .B(n4112), .Y(
        top_core_KE_n5679) );
  AND2X2 top_core_KE_U5762 ( .A(top_core_KE_key_mem_14__125_), .B(n4069), .Y(
        top_core_KE_n5685) );
  AND2X2 top_core_KE_U5454 ( .A(top_core_KE_key_mem_14__81_), .B(n4090), .Y(
        top_core_KE_n5421) );
  AND2X2 top_core_KE_U5335 ( .A(top_core_KE_key_mem_14__64_), .B(n4079), .Y(
        top_core_KE_n5319) );
  AND2X2 top_core_KE_U5195 ( .A(top_core_KE_key_mem_14__44_), .B(n4115), .Y(
        top_core_KE_n5199) );
  AND2X2 top_core_KE_U5202 ( .A(top_core_KE_key_mem_14__45_), .B(n4113), .Y(
        top_core_KE_n5205) );
  AND2X2 top_core_KE_U5006 ( .A(top_core_KE_key_mem_14__17_), .B(n4087), .Y(
        top_core_KE_n5037) );
  AND2X2 top_core_KE_U5447 ( .A(top_core_KE_key_mem_14__80_), .B(n4072), .Y(
        top_core_KE_n5415) );
  AND2X2 top_core_KE_U4999 ( .A(top_core_KE_key_mem_14__16_), .B(n4087), .Y(
        top_core_KE_n5031) );
  AND2X2 top_core_KE_U5566 ( .A(top_core_KE_key_mem_14__97_), .B(n4084), .Y(
        top_core_KE_n5517) );
  AND2X2 top_core_KE_U5125 ( .A(top_core_KE_key_mem_14__34_), .B(n4094), .Y(
        top_core_KE_n5139) );
  AND2X2 top_core_KE_U5398 ( .A(top_core_KE_key_mem_14__73_), .B(n4068), .Y(
        top_core_KE_n5373) );
  AND2X2 top_core_KE_U5405 ( .A(top_core_KE_key_mem_14__74_), .B(n4093), .Y(
        top_core_KE_n5379) );
  AND2X2 top_core_KE_U5062 ( .A(top_core_KE_key_mem_14__25_), .B(n4080), .Y(
        top_core_KE_n5085) );
  AND2X2 top_core_KE_U5069 ( .A(top_core_KE_key_mem_14__26_), .B(n4083), .Y(
        top_core_KE_n5091) );
  AND2X2 top_core_KE_U4894 ( .A(top_core_KE_key_mem_14__1_), .B(n4095), .Y(
        top_core_KE_n4941) );
  AND2X2 top_core_KE_U5622 ( .A(top_core_KE_key_mem_14__105_), .B(n4034), .Y(
        top_core_KE_n5565) );
  AND2X2 top_core_KE_U5629 ( .A(top_core_KE_key_mem_14__106_), .B(n4079), .Y(
        top_core_KE_n5571) );
  AND2X2 top_core_KE_U5286 ( .A(top_core_KE_key_mem_14__57_), .B(n4089), .Y(
        top_core_KE_n5277) );
  AND2X2 top_core_KE_U5293 ( .A(top_core_KE_key_mem_14__58_), .B(n4074), .Y(
        top_core_KE_n5283) );
  AND2X2 top_core_KE_U5118 ( .A(top_core_KE_key_mem_14__33_), .B(n4082), .Y(
        top_core_KE_n5133) );
  AND2X2 top_core_KE_U5573 ( .A(top_core_KE_key_mem_14__98_), .B(n4112), .Y(
        top_core_KE_n5523) );
  AND2X2 top_core_KE_U5517 ( .A(top_core_KE_key_mem_14__90_), .B(n4072), .Y(
        top_core_KE_n5475) );
  AND2X2 top_core_KE_U4957 ( .A(top_core_KE_key_mem_14__10_), .B(n4090), .Y(
        top_core_KE_n4995) );
  AND2X2 top_core_KE_U5678 ( .A(top_core_KE_key_mem_14__113_), .B(n4068), .Y(
        top_core_KE_n5613) );
  AND2X2 top_core_KE_U5181 ( .A(top_core_KE_key_mem_14__42_), .B(n4071), .Y(
        top_core_KE_n5187) );
  AND2X2 top_core_KE_U5342 ( .A(top_core_KE_key_mem_14__65_), .B(n4079), .Y(
        top_core_KE_n5325) );
  AND2X2 top_core_KE_U5741 ( .A(top_core_KE_key_mem_14__122_), .B(n4071), .Y(
        top_core_KE_n5667) );
  AND2X2 top_core_KE_U4901 ( .A(top_core_KE_key_mem_14__2_), .B(n4094), .Y(
        top_core_KE_n4947) );
  AND2X2 top_core_KE_U5503 ( .A(top_core_KE_key_mem_14__88_), .B(n4073), .Y(
        top_core_KE_n5463) );
  AND2X2 top_core_KE_U4943 ( .A(top_core_KE_key_mem_14__8_), .B(n4091), .Y(
        top_core_KE_n4983) );
  AND2X2 top_core_KE_U5237 ( .A(top_core_KE_key_mem_14__50_), .B(n4091), .Y(
        top_core_KE_n5235) );
  AND2X2 top_core_KE_U5167 ( .A(top_core_KE_key_mem_14__40_), .B(n4067), .Y(
        top_core_KE_n5175) );
  AND2X2 top_core_KE_U5510 ( .A(top_core_KE_key_mem_14__89_), .B(n4073), .Y(
        top_core_KE_n5469) );
  AND2X2 top_core_KE_U4950 ( .A(top_core_KE_key_mem_14__9_), .B(n4091), .Y(
        top_core_KE_n4989) );
  AND2X2 top_core_KE_U5174 ( .A(top_core_KE_key_mem_14__41_), .B(n4114), .Y(
        top_core_KE_n5181) );
  AND2X2 top_core_KE_U5734 ( .A(top_core_KE_key_mem_14__121_), .B(n4079), .Y(
        top_core_KE_n5661) );
  AND2X2 top_core_KE_U5461 ( .A(top_core_KE_key_mem_14__82_), .B(n4093), .Y(
        top_core_KE_n5427) );
  AND2X2 top_core_KE_U5727 ( .A(top_core_KE_key_mem_14__120_), .B(n4078), .Y(
        top_core_KE_n5655) );
  MX2X1 top_core_KE_U5131 ( .A(top_core_KE_key_mem_12__35_), .B(
        top_core_KE_key_mem_13__35_), .S0(n4046), .Y(top_core_KE_n5144) );
  MX2X1 top_core_KE_U5257 ( .A(top_core_KE_key_mem_12__53_), .B(
        top_core_KE_key_mem_13__53_), .S0(n4047), .Y(top_core_KE_n5252) );
  MX2X1 top_core_KE_U5502 ( .A(top_core_KE_key_mem_12__88_), .B(
        top_core_KE_key_mem_13__88_), .S0(n4101), .Y(top_core_KE_n5462) );
  MX2X1 top_core_KE_U5607 ( .A(top_core_KE_key_mem_12__103_), .B(
        top_core_KE_key_mem_13__103_), .S0(n4065), .Y(top_core_KE_n5552) );
  MX2X1 top_core_KE_U5159 ( .A(top_core_KE_key_mem_12__39_), .B(
        top_core_KE_key_mem_13__39_), .S0(n4063), .Y(top_core_KE_n5168) );
  MX2X1 top_core_KE_U5439 ( .A(top_core_KE_key_mem_12__79_), .B(
        top_core_KE_key_mem_13__79_), .S0(n4061), .Y(top_core_KE_n5408) );
  MX2X1 top_core_KE_U5271 ( .A(top_core_KE_key_mem_12__55_), .B(
        top_core_KE_key_mem_13__55_), .S0(n4065), .Y(top_core_KE_n5264) );
  MX2X1 top_core_KE_U5719 ( .A(top_core_KE_key_mem_12__119_), .B(
        top_core_KE_key_mem_13__119_), .S0(n4061), .Y(top_core_KE_n5648) );
  MX2X1 top_core_KE_U5103 ( .A(top_core_KE_key_mem_12__31_), .B(
        top_core_KE_key_mem_13__31_), .S0(n4065), .Y(top_core_KE_n5120) );
  MX2X1 top_core_KE_U4935 ( .A(top_core_KE_key_mem_12__7_), .B(
        top_core_KE_key_mem_13__7_), .S0(n4059), .Y(top_core_KE_n4976) );
  MX2X1 top_core_KE_U5663 ( .A(top_core_KE_key_mem_12__111_), .B(
        top_core_KE_key_mem_13__111_), .S0(n4063), .Y(top_core_KE_n5600) );
  MX2X1 top_core_KE_U5495 ( .A(top_core_KE_key_mem_12__87_), .B(
        top_core_KE_key_mem_13__87_), .S0(n4065), .Y(top_core_KE_n5456) );
  MX2X1 top_core_KE_U5047 ( .A(top_core_KE_key_mem_12__23_), .B(
        top_core_KE_key_mem_13__23_), .S0(n4063), .Y(top_core_KE_n5072) );
  MX2X1 top_core_KE_U5327 ( .A(top_core_KE_key_mem_12__63_), .B(
        top_core_KE_key_mem_13__63_), .S0(n4062), .Y(top_core_KE_n5312) );
  MX2X1 top_core_KE_U5551 ( .A(top_core_KE_key_mem_12__95_), .B(
        top_core_KE_key_mem_13__95_), .S0(n4059), .Y(top_core_KE_n5504) );
  MX2X1 top_core_KE_U4991 ( .A(top_core_KE_key_mem_12__15_), .B(
        top_core_KE_key_mem_13__15_), .S0(n4061), .Y(top_core_KE_n5024) );
  MX2X1 top_core_KE_U5691 ( .A(top_core_KE_key_mem_12__115_), .B(
        top_core_KE_key_mem_13__115_), .S0(n4062), .Y(top_core_KE_n5624) );
  MX2X1 top_core_KE_U5075 ( .A(top_core_KE_key_mem_12__27_), .B(
        top_core_KE_key_mem_13__27_), .S0(n4064), .Y(top_core_KE_n5096) );
  MX2X1 top_core_KE_U5355 ( .A(top_core_KE_key_mem_12__67_), .B(
        top_core_KE_key_mem_13__67_), .S0(n4060), .Y(top_core_KE_n5336) );
  MX2X1 top_core_KE_U5635 ( .A(top_core_KE_key_mem_12__107_), .B(
        top_core_KE_key_mem_13__107_), .S0(n4064), .Y(top_core_KE_n5576) );
  MX2X1 top_core_KE_U5019 ( .A(top_core_KE_key_mem_12__19_), .B(
        top_core_KE_key_mem_13__19_), .S0(n4062), .Y(top_core_KE_n5048) );
  MX2X1 top_core_KE_U5299 ( .A(top_core_KE_key_mem_12__59_), .B(
        top_core_KE_key_mem_13__59_), .S0(n4063), .Y(top_core_KE_n5288) );
  MX2X1 top_core_KE_U5579 ( .A(top_core_KE_key_mem_12__99_), .B(
        top_core_KE_key_mem_13__99_), .S0(n4063), .Y(top_core_KE_n5528) );
  MX2X1 top_core_KE_U5243 ( .A(top_core_KE_key_mem_12__51_), .B(
        top_core_KE_key_mem_13__51_), .S0(n4063), .Y(top_core_KE_n5240) );
  MX2X1 top_core_KE_U5467 ( .A(top_core_KE_key_mem_12__83_), .B(
        top_core_KE_key_mem_13__83_), .S0(n4063), .Y(top_core_KE_n5432) );
  MX2X1 top_core_KE_U5152 ( .A(top_core_KE_key_mem_12__38_), .B(
        top_core_KE_key_mem_13__38_), .S0(n4064), .Y(top_core_KE_n5162) );
  MX2X1 top_core_KE_U5432 ( .A(top_core_KE_key_mem_12__78_), .B(
        top_core_KE_key_mem_13__78_), .S0(n4060), .Y(top_core_KE_n5402) );
  MX2X1 top_core_KE_U5096 ( .A(top_core_KE_key_mem_12__30_), .B(
        top_core_KE_key_mem_13__30_), .S0(n4065), .Y(top_core_KE_n5114) );
  MX2X1 top_core_KE_U5656 ( .A(top_core_KE_key_mem_12__110_), .B(
        top_core_KE_key_mem_13__110_), .S0(n4063), .Y(top_core_KE_n5594) );
  MX2X1 top_core_KE_U5320 ( .A(top_core_KE_key_mem_12__62_), .B(
        top_core_KE_key_mem_13__62_), .S0(n4062), .Y(top_core_KE_n5306) );
  MX2X1 top_core_KE_U5523 ( .A(top_core_KE_key_mem_12__91_), .B(
        top_core_KE_key_mem_13__91_), .S0(n4062), .Y(top_core_KE_n5480) );
  MX2X1 top_core_KE_U4963 ( .A(top_core_KE_key_mem_12__11_), .B(
        top_core_KE_key_mem_13__11_), .S0(n4060), .Y(top_core_KE_n5000) );
  MX2X1 top_core_KE_U5712 ( .A(top_core_KE_key_mem_12__118_), .B(
        top_core_KE_key_mem_13__118_), .S0(n4061), .Y(top_core_KE_n5642) );
  MX2X1 top_core_KE_U4928 ( .A(top_core_KE_key_mem_12__6_), .B(
        top_core_KE_key_mem_13__6_), .S0(n4059), .Y(top_core_KE_n4970) );
  MX2X1 top_core_KE_U5376 ( .A(top_core_KE_key_mem_12__70_), .B(
        top_core_KE_key_mem_13__70_), .S0(n4059), .Y(top_core_KE_n5354) );
  MX2X1 top_core_KE_U5747 ( .A(top_core_KE_key_mem_12__123_), .B(
        top_core_KE_key_mem_13__123_), .S0(n4060), .Y(top_core_KE_n5672) );
  MX2X1 top_core_KE_U5187 ( .A(top_core_KE_key_mem_12__43_), .B(
        top_core_KE_key_mem_13__43_), .S0(n4060), .Y(top_core_KE_n5192) );
  MX2X1 top_core_KE_U5040 ( .A(top_core_KE_key_mem_12__22_), .B(
        top_core_KE_key_mem_13__22_), .S0(n4063), .Y(top_core_KE_n5066) );
  MX2X1 top_core_KE_U5264 ( .A(top_core_KE_key_mem_12__54_), .B(
        top_core_KE_key_mem_13__54_), .S0(n4065), .Y(top_core_KE_n5258) );
  MX2X1 top_core_KE_U5698 ( .A(top_core_KE_key_mem_12__116_), .B(
        top_core_KE_key_mem_13__116_), .S0(n4061), .Y(top_core_KE_n5630) );
  MX2X1 top_core_KE_U5145 ( .A(top_core_KE_key_mem_12__37_), .B(
        top_core_KE_key_mem_13__37_), .S0(n4065), .Y(top_core_KE_n5156) );
  MX2X1 top_core_KE_U5586 ( .A(top_core_KE_key_mem_12__100_), .B(
        top_core_KE_key_mem_13__100_), .S0(n4064), .Y(top_core_KE_n5534) );
  MX2X1 top_core_KE_U5593 ( .A(top_core_KE_key_mem_12__101_), .B(
        top_core_KE_key_mem_13__101_), .S0(n4065), .Y(top_core_KE_n5540) );
  MX2X1 top_core_KE_U5362 ( .A(top_core_KE_key_mem_12__68_), .B(
        top_core_KE_key_mem_13__68_), .S0(n4060), .Y(top_core_KE_n5342) );
  MX2X1 top_core_KE_U5488 ( .A(top_core_KE_key_mem_12__86_), .B(
        top_core_KE_key_mem_13__86_), .S0(n4064), .Y(top_core_KE_n5450) );
  MX2X1 top_core_KE_U5138 ( .A(top_core_KE_key_mem_12__36_), .B(
        top_core_KE_key_mem_13__36_), .S0(n4065), .Y(top_core_KE_n5150) );
  MX2X1 top_core_KE_U5425 ( .A(top_core_KE_key_mem_12__77_), .B(
        top_core_KE_key_mem_13__77_), .S0(n4061), .Y(top_core_KE_n5396) );
  MX2X1 top_core_KE_U5418 ( .A(top_core_KE_key_mem_12__76_), .B(
        top_core_KE_key_mem_13__76_), .S0(n4059), .Y(top_core_KE_n5390) );
  MX2X1 top_core_KE_U5089 ( .A(top_core_KE_key_mem_12__29_), .B(
        top_core_KE_key_mem_13__29_), .S0(n4064), .Y(top_core_KE_n5108) );
  MX2X1 top_core_KE_U5082 ( .A(top_core_KE_key_mem_12__28_), .B(
        top_core_KE_key_mem_13__28_), .S0(n4064), .Y(top_core_KE_n5102) );
  MX2X1 top_core_KE_U5649 ( .A(top_core_KE_key_mem_12__109_), .B(
        top_core_KE_key_mem_13__109_), .S0(n4064), .Y(top_core_KE_n5588) );
  MX2X1 top_core_KE_U5642 ( .A(top_core_KE_key_mem_12__108_), .B(
        top_core_KE_key_mem_13__108_), .S0(n4064), .Y(top_core_KE_n5582) );
  MX2X1 top_core_KE_U5313 ( .A(top_core_KE_key_mem_12__61_), .B(
        top_core_KE_key_mem_13__61_), .S0(n4063), .Y(top_core_KE_n5300) );
  MX2X1 top_core_KE_U5306 ( .A(top_core_KE_key_mem_12__60_), .B(
        top_core_KE_key_mem_13__60_), .S0(n4063), .Y(top_core_KE_n5294) );
  MX2X1 top_core_KE_U4984 ( .A(top_core_KE_key_mem_12__14_), .B(
        top_core_KE_key_mem_13__14_), .S0(n4061), .Y(top_core_KE_n5018) );
  MX2X1 top_core_KE_U5705 ( .A(top_core_KE_key_mem_12__117_), .B(
        top_core_KE_key_mem_13__117_), .S0(n4061), .Y(top_core_KE_n5636) );
  MX2X1 top_core_KE_U5369 ( .A(top_core_KE_key_mem_12__69_), .B(
        top_core_KE_key_mem_13__69_), .S0(n4059), .Y(top_core_KE_n5348) );
  MX2X1 top_core_KE_U5026 ( .A(top_core_KE_key_mem_12__20_), .B(
        top_core_KE_key_mem_13__20_), .S0(n4062), .Y(top_core_KE_n5054) );
  MX2X1 top_core_KE_U5033 ( .A(top_core_KE_key_mem_12__21_), .B(
        top_core_KE_key_mem_13__21_), .S0(n4063), .Y(top_core_KE_n5060) );
  MX2X1 top_core_KE_U4921 ( .A(top_core_KE_key_mem_12__5_), .B(
        top_core_KE_key_mem_13__5_), .S0(n4059), .Y(top_core_KE_n4964) );
  MX2X1 top_core_KE_U5250 ( .A(top_core_KE_key_mem_12__52_), .B(
        top_core_KE_key_mem_13__52_), .S0(n4064), .Y(top_core_KE_n5246) );
  MX2X1 top_core_KE_U5768 ( .A(top_core_KE_key_mem_12__126_), .B(
        top_core_KE_key_mem_13__126_), .S0(n4059), .Y(top_core_KE_n5690) );
  MX2X1 top_core_KE_U5684 ( .A(top_core_KE_key_mem_12__114_), .B(
        top_core_KE_key_mem_13__114_), .S0(n4062), .Y(top_core_KE_n5618) );
  MX2X1 top_core_KE_U5348 ( .A(top_core_KE_key_mem_12__66_), .B(
        top_core_KE_key_mem_13__66_), .S0(n4060), .Y(top_core_KE_n5330) );
  MX2X1 top_core_KE_U5474 ( .A(top_core_KE_key_mem_12__84_), .B(
        top_core_KE_key_mem_13__84_), .S0(n4063), .Y(top_core_KE_n5438) );
  MX2X1 top_core_KE_U5481 ( .A(top_core_KE_key_mem_12__85_), .B(
        top_core_KE_key_mem_13__85_), .S0(n4064), .Y(top_core_KE_n5444) );
  MX2X1 top_core_KE_U5012 ( .A(top_core_KE_key_mem_12__18_), .B(
        top_core_KE_key_mem_13__18_), .S0(n4062), .Y(top_core_KE_n5042) );
  MX2X1 top_core_KE_U5110 ( .A(top_core_KE_key_mem_12__32_), .B(
        top_core_KE_key_mem_13__32_), .S0(n4065), .Y(top_core_KE_n5126) );
  MX2X1 top_core_KE_U5054 ( .A(top_core_KE_key_mem_12__24_), .B(
        top_core_KE_key_mem_13__24_), .S0(n4063), .Y(top_core_KE_n5078) );
  MX2X1 top_core_KE_U5614 ( .A(top_core_KE_key_mem_12__104_), .B(
        top_core_KE_key_mem_13__104_), .S0(n4065), .Y(top_core_KE_n5558) );
  MX2X1 top_core_KE_U5278 ( .A(top_core_KE_key_mem_12__56_), .B(
        top_core_KE_key_mem_13__56_), .S0(n4065), .Y(top_core_KE_n5270) );
  MX2X1 top_core_KE_U5558 ( .A(top_core_KE_key_mem_12__96_), .B(
        top_core_KE_key_mem_13__96_), .S0(n4060), .Y(top_core_KE_n5510) );
  MX2X1 top_core_KE_U5530 ( .A(top_core_KE_key_mem_12__92_), .B(
        top_core_KE_key_mem_13__92_), .S0(n4060), .Y(top_core_KE_n5486) );
  MX2X1 top_core_KE_U5537 ( .A(top_core_KE_key_mem_12__93_), .B(
        top_core_KE_key_mem_13__93_), .S0(n4059), .Y(top_core_KE_n5492) );
  MX2X1 top_core_KE_U4970 ( .A(top_core_KE_key_mem_12__12_), .B(
        top_core_KE_key_mem_13__12_), .S0(n4060), .Y(top_core_KE_n5006) );
  MX2X1 top_core_KE_U4977 ( .A(top_core_KE_key_mem_12__13_), .B(
        top_core_KE_key_mem_13__13_), .S0(n4061), .Y(top_core_KE_n5012) );
  MX2X1 top_core_KE_U5229 ( .A(top_core_KE_key_mem_12__49_), .B(
        top_core_KE_key_mem_13__49_), .S0(n4060), .Y(top_core_KE_n5228) );
  MX2X1 top_core_KE_U5222 ( .A(top_core_KE_key_mem_12__48_), .B(
        top_core_KE_key_mem_13__48_), .S0(n4060), .Y(top_core_KE_n5222) );
  MX2X1 top_core_KE_U5670 ( .A(top_core_KE_key_mem_12__112_), .B(
        top_core_KE_key_mem_13__112_), .S0(n4063), .Y(top_core_KE_n5606) );
  MX2X1 top_core_KE_U4886 ( .A(top_core_KE_key_mem_12__0_), .B(
        top_core_KE_key_mem_13__0_), .S0(n4059), .Y(top_core_KE_n4934) );
  MX2X1 top_core_KE_U5754 ( .A(top_core_KE_key_mem_12__124_), .B(
        top_core_KE_key_mem_13__124_), .S0(n4059), .Y(top_core_KE_n5678) );
  MX2X1 top_core_KE_U5453 ( .A(top_core_KE_key_mem_12__81_), .B(
        top_core_KE_key_mem_13__81_), .S0(n4062), .Y(top_core_KE_n5420) );
  MX2X1 top_core_KE_U5334 ( .A(top_core_KE_key_mem_12__64_), .B(
        top_core_KE_key_mem_13__64_), .S0(n4061), .Y(top_core_KE_n5318) );
  MX2X1 top_core_KE_U5194 ( .A(top_core_KE_key_mem_12__44_), .B(
        top_core_KE_key_mem_13__44_), .S0(n4059), .Y(top_core_KE_n5198) );
  MX2X1 top_core_KE_U5201 ( .A(top_core_KE_key_mem_12__45_), .B(
        top_core_KE_key_mem_13__45_), .S0(n4059), .Y(top_core_KE_n5204) );
  MX2X1 top_core_KE_U5005 ( .A(top_core_KE_key_mem_12__17_), .B(
        top_core_KE_key_mem_13__17_), .S0(n4062), .Y(top_core_KE_n5036) );
  MX2X1 top_core_KE_U5446 ( .A(top_core_KE_key_mem_12__80_), .B(
        top_core_KE_key_mem_13__80_), .S0(n4061), .Y(top_core_KE_n5414) );
  MX2X1 top_core_KE_U4998 ( .A(top_core_KE_key_mem_12__16_), .B(
        top_core_KE_key_mem_13__16_), .S0(n4061), .Y(top_core_KE_n5030) );
  MX2X1 top_core_KE_U5565 ( .A(top_core_KE_key_mem_12__97_), .B(
        top_core_KE_key_mem_13__97_), .S0(n4061), .Y(top_core_KE_n5516) );
  MX2X1 top_core_KE_U5124 ( .A(top_core_KE_key_mem_12__34_), .B(
        top_core_KE_key_mem_13__34_), .S0(n4065), .Y(top_core_KE_n5138) );
  MX2X1 top_core_KE_U5061 ( .A(top_core_KE_key_mem_12__25_), .B(
        top_core_KE_key_mem_13__25_), .S0(n4063), .Y(top_core_KE_n5084) );
  MX2X1 top_core_KE_U5068 ( .A(top_core_KE_key_mem_12__26_), .B(
        top_core_KE_key_mem_13__26_), .S0(n4064), .Y(top_core_KE_n5090) );
  MX2X1 top_core_KE_U4893 ( .A(top_core_KE_key_mem_12__1_), .B(
        top_core_KE_key_mem_13__1_), .S0(n4059), .Y(top_core_KE_n4940) );
  MX2X1 top_core_KE_U5621 ( .A(top_core_KE_key_mem_12__105_), .B(
        top_core_KE_key_mem_13__105_), .S0(n4065), .Y(top_core_KE_n5564) );
  MX2X1 top_core_KE_U5628 ( .A(top_core_KE_key_mem_12__106_), .B(
        top_core_KE_key_mem_13__106_), .S0(n4064), .Y(top_core_KE_n5570) );
  MX2X1 top_core_KE_U5285 ( .A(top_core_KE_key_mem_12__57_), .B(
        top_core_KE_key_mem_13__57_), .S0(n4064), .Y(top_core_KE_n5276) );
  MX2X1 top_core_KE_U5292 ( .A(top_core_KE_key_mem_12__58_), .B(
        top_core_KE_key_mem_13__58_), .S0(n4064), .Y(top_core_KE_n5282) );
  MX2X1 top_core_KE_U5117 ( .A(top_core_KE_key_mem_12__33_), .B(
        top_core_KE_key_mem_13__33_), .S0(n4065), .Y(top_core_KE_n5132) );
  MX2X1 top_core_KE_U5572 ( .A(top_core_KE_key_mem_12__98_), .B(
        top_core_KE_key_mem_13__98_), .S0(n4062), .Y(top_core_KE_n5522) );
  MX2X1 top_core_KE_U5516 ( .A(top_core_KE_key_mem_12__90_), .B(
        top_core_KE_key_mem_13__90_), .S0(n4064), .Y(top_core_KE_n5474) );
  MX2X1 top_core_KE_U4956 ( .A(top_core_KE_key_mem_12__10_), .B(
        top_core_KE_key_mem_13__10_), .S0(n4060), .Y(top_core_KE_n4994) );
  MX2X1 top_core_KE_U5677 ( .A(top_core_KE_key_mem_12__113_), .B(
        top_core_KE_key_mem_13__113_), .S0(n4062), .Y(top_core_KE_n5612) );
  MX2X1 top_core_KE_U5180 ( .A(top_core_KE_key_mem_12__42_), .B(
        top_core_KE_key_mem_13__42_), .S0(n4061), .Y(top_core_KE_n5186) );
  MX2X1 top_core_KE_U5341 ( .A(top_core_KE_key_mem_12__65_), .B(
        top_core_KE_key_mem_13__65_), .S0(n4061), .Y(top_core_KE_n5324) );
  MX2X1 top_core_KE_U5740 ( .A(top_core_KE_key_mem_12__122_), .B(
        top_core_KE_key_mem_13__122_), .S0(n4059), .Y(top_core_KE_n5666) );
  MX2X1 top_core_KE_U4900 ( .A(top_core_KE_key_mem_12__2_), .B(
        top_core_KE_key_mem_13__2_), .S0(n4059), .Y(top_core_KE_n4946) );
  MX2X1 top_core_KE_U4942 ( .A(top_core_KE_key_mem_12__8_), .B(
        top_core_KE_key_mem_13__8_), .S0(n4061), .Y(top_core_KE_n4982) );
  MX2X1 top_core_KE_U5236 ( .A(top_core_KE_key_mem_12__50_), .B(
        top_core_KE_key_mem_13__50_), .S0(n4062), .Y(top_core_KE_n5234) );
  MX2X1 top_core_KE_U5166 ( .A(top_core_KE_key_mem_12__40_), .B(
        top_core_KE_key_mem_13__40_), .S0(n4062), .Y(top_core_KE_n5174) );
  MX2X1 top_core_KE_U5509 ( .A(top_core_KE_key_mem_12__89_), .B(
        top_core_KE_key_mem_13__89_), .S0(n4065), .Y(top_core_KE_n5468) );
  MX2X1 top_core_KE_U4949 ( .A(top_core_KE_key_mem_12__9_), .B(
        top_core_KE_key_mem_13__9_), .S0(n4060), .Y(top_core_KE_n4988) );
  MX2X1 top_core_KE_U5173 ( .A(top_core_KE_key_mem_12__41_), .B(
        top_core_KE_key_mem_13__41_), .S0(n4062), .Y(top_core_KE_n5180) );
  MX2X1 top_core_KE_U5733 ( .A(top_core_KE_key_mem_12__121_), .B(
        top_core_KE_key_mem_13__121_), .S0(n4060), .Y(top_core_KE_n5660) );
  MX2X1 top_core_KE_U5460 ( .A(top_core_KE_key_mem_12__82_), .B(
        top_core_KE_key_mem_13__82_), .S0(n4062), .Y(top_core_KE_n5426) );
  MX2X1 top_core_KE_U5726 ( .A(top_core_KE_key_mem_12__120_), .B(
        top_core_KE_key_mem_13__120_), .S0(n4060), .Y(top_core_KE_n5654) );
  MX2X1 top_core_KE_U5383 ( .A(top_core_KE_key_mem_12__71_), .B(
        top_core_KE_key_mem_13__71_), .S0(n4058), .Y(top_core_KE_n5360) );
  MX2X1 top_core_KE_U5215 ( .A(top_core_KE_key_mem_12__47_), .B(
        top_core_KE_key_mem_13__47_), .S0(n4058), .Y(top_core_KE_n5216) );
  MX2X1 top_core_KE_U5775 ( .A(top_core_KE_key_mem_12__127_), .B(
        top_core_KE_key_mem_13__127_), .S0(n4058), .Y(top_core_KE_n5696) );
  MX2X1 top_core_KE_U5782 ( .A(top_core_KE_key_mem_12__128_), .B(
        top_core_KE_key_mem_13__128_), .S0(n4058), .Y(top_core_KE_n5702) );
  MX2X1 top_core_KE_U5411 ( .A(top_core_KE_key_mem_12__75_), .B(
        top_core_KE_key_mem_13__75_), .S0(n4058), .Y(top_core_KE_n5384) );
  MX2X1 top_core_KE_U4907 ( .A(top_core_KE_key_mem_12__3_), .B(
        top_core_KE_key_mem_13__3_), .S0(n4058), .Y(top_core_KE_n4952) );
  MX2X1 top_core_KE_U5600 ( .A(top_core_KE_key_mem_12__102_), .B(
        top_core_KE_key_mem_13__102_), .S0(n4058), .Y(top_core_KE_n5546) );
  MX2X1 top_core_KE_U5544 ( .A(top_core_KE_key_mem_12__94_), .B(
        top_core_KE_key_mem_13__94_), .S0(n4058), .Y(top_core_KE_n5498) );
  MX2X1 top_core_KE_U5208 ( .A(top_core_KE_key_mem_12__46_), .B(
        top_core_KE_key_mem_13__46_), .S0(n4058), .Y(top_core_KE_n5210) );
  MX2X1 top_core_KE_U4914 ( .A(top_core_KE_key_mem_12__4_), .B(
        top_core_KE_key_mem_13__4_), .S0(n4058), .Y(top_core_KE_n4958) );
  MX2X1 top_core_KE_U5390 ( .A(top_core_KE_key_mem_12__72_), .B(
        top_core_KE_key_mem_13__72_), .S0(n4058), .Y(top_core_KE_n5366) );
  MX2X1 top_core_KE_U5761 ( .A(top_core_KE_key_mem_12__125_), .B(
        top_core_KE_key_mem_13__125_), .S0(n4058), .Y(top_core_KE_n5684) );
  MX2X1 top_core_KE_U5397 ( .A(top_core_KE_key_mem_12__73_), .B(
        top_core_KE_key_mem_13__73_), .S0(n4058), .Y(top_core_KE_n5372) );
  MX2X1 top_core_KE_U5404 ( .A(top_core_KE_key_mem_12__74_), .B(
        top_core_KE_key_mem_13__74_), .S0(n4058), .Y(top_core_KE_n5378) );
  MX4X1 top_core_KE_U5787 ( .A(top_core_KE_key_mem_0__128_), .B(
        top_core_KE_key_mem_1__128_), .C(top_core_KE_key_mem_2__128_), .D(
        top_core_KE_key_mem_3__128_), .S0(n4033), .S1(n3989), .Y(
        top_core_KE_n5707) );
  MX4X1 top_core_KE_U5611 ( .A(top_core_KE_key_mem_4__103_), .B(
        top_core_KE_key_mem_5__103_), .C(top_core_KE_key_mem_6__103_), .D(
        top_core_KE_key_mem_7__103_), .S0(n4104), .S1(n4005), .Y(
        top_core_KE_n5556) );
  MX4X1 top_core_KE_U5163 ( .A(top_core_KE_key_mem_4__39_), .B(
        top_core_KE_key_mem_5__39_), .C(top_core_KE_key_mem_6__39_), .D(
        top_core_KE_key_mem_7__39_), .S0(n4035), .S1(n3989), .Y(
        top_core_KE_n5172) );
  MX4X1 top_core_KE_U5443 ( .A(top_core_KE_key_mem_4__79_), .B(
        top_core_KE_key_mem_5__79_), .C(top_core_KE_key_mem_6__79_), .D(
        top_core_KE_key_mem_7__79_), .S0(n4053), .S1(n4010), .Y(
        top_core_KE_n5412) );
  MX4X1 top_core_KE_U5275 ( .A(top_core_KE_key_mem_4__55_), .B(
        top_core_KE_key_mem_5__55_), .C(top_core_KE_key_mem_6__55_), .D(
        top_core_KE_key_mem_7__55_), .S0(n4039), .S1(n3992), .Y(
        top_core_KE_n5268) );
  MX4X1 top_core_KE_U5723 ( .A(top_core_KE_key_mem_4__119_), .B(
        top_core_KE_key_mem_5__119_), .C(top_core_KE_key_mem_6__119_), .D(
        top_core_KE_key_mem_7__119_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5652) );
  MX4X1 top_core_KE_U5107 ( .A(top_core_KE_key_mem_4__31_), .B(
        top_core_KE_key_mem_5__31_), .C(top_core_KE_key_mem_6__31_), .D(
        top_core_KE_key_mem_7__31_), .S0(n4050), .S1(n4002), .Y(
        top_core_KE_n5124) );
  MX4X1 top_core_KE_U4939 ( .A(top_core_KE_key_mem_4__7_), .B(
        top_core_KE_key_mem_5__7_), .C(top_core_KE_key_mem_6__7_), .D(
        top_core_KE_key_mem_7__7_), .S0(n4045), .S1(n3997), .Y(
        top_core_KE_n4980) );
  MX4X1 top_core_KE_U5387 ( .A(top_core_KE_key_mem_4__71_), .B(
        top_core_KE_key_mem_5__71_), .C(top_core_KE_key_mem_6__71_), .D(
        top_core_KE_key_mem_7__71_), .S0(n4043), .S1(n3995), .Y(
        top_core_KE_n5364) );
  MX4X1 top_core_KE_U5667 ( .A(top_core_KE_key_mem_4__111_), .B(
        top_core_KE_key_mem_5__111_), .C(top_core_KE_key_mem_6__111_), .D(
        top_core_KE_key_mem_7__111_), .S0(n4052), .S1(n4006), .Y(
        top_core_KE_n5604) );
  MX4X1 top_core_KE_U5499 ( .A(top_core_KE_key_mem_4__87_), .B(
        top_core_KE_key_mem_5__87_), .C(top_core_KE_key_mem_6__87_), .D(
        top_core_KE_key_mem_7__87_), .S0(n4057), .S1(n4011), .Y(
        top_core_KE_n5460) );
  MX4X1 top_core_KE_U5051 ( .A(top_core_KE_key_mem_4__23_), .B(
        top_core_KE_key_mem_5__23_), .C(top_core_KE_key_mem_6__23_), .D(
        top_core_KE_key_mem_7__23_), .S0(n4048), .S1(n4000), .Y(
        top_core_KE_n5076) );
  MX4X1 top_core_KE_U5331 ( .A(top_core_KE_key_mem_4__63_), .B(
        top_core_KE_key_mem_5__63_), .C(top_core_KE_key_mem_6__63_), .D(
        top_core_KE_key_mem_7__63_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5316) );
  MX4X1 top_core_KE_U5555 ( .A(top_core_KE_key_mem_4__95_), .B(
        top_core_KE_key_mem_5__95_), .C(top_core_KE_key_mem_6__95_), .D(
        top_core_KE_key_mem_7__95_), .S0(n4096), .S1(n4003), .Y(
        top_core_KE_n5508) );
  MX4X1 top_core_KE_U4995 ( .A(top_core_KE_key_mem_4__15_), .B(
        top_core_KE_key_mem_5__15_), .C(top_core_KE_key_mem_6__15_), .D(
        top_core_KE_key_mem_7__15_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5028) );
  MX4X1 top_core_KE_U5219 ( .A(top_core_KE_key_mem_4__47_), .B(
        top_core_KE_key_mem_5__47_), .C(top_core_KE_key_mem_6__47_), .D(
        top_core_KE_key_mem_7__47_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5220) );
  MX4X1 top_core_KE_U5779 ( .A(top_core_KE_key_mem_4__127_), .B(
        top_core_KE_key_mem_5__127_), .C(top_core_KE_key_mem_6__127_), .D(
        top_core_KE_key_mem_7__127_), .S0(n4055), .S1(n4008), .Y(
        top_core_KE_n5700) );
  MX4X1 top_core_KE_U5786 ( .A(top_core_KE_key_mem_4__128_), .B(
        top_core_KE_key_mem_5__128_), .C(top_core_KE_key_mem_6__128_), .D(
        top_core_KE_key_mem_7__128_), .S0(n4042), .S1(n4007), .Y(
        top_core_KE_n5706) );
  MX4X1 top_core_KE_U5135 ( .A(top_core_KE_key_mem_4__35_), .B(
        top_core_KE_key_mem_5__35_), .C(top_core_KE_key_mem_6__35_), .D(
        top_core_KE_key_mem_7__35_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5148) );
  MX4X1 top_core_KE_U5415 ( .A(top_core_KE_key_mem_4__75_), .B(
        top_core_KE_key_mem_5__75_), .C(top_core_KE_key_mem_6__75_), .D(
        top_core_KE_key_mem_7__75_), .S0(n4041), .S1(n4010), .Y(
        top_core_KE_n5388) );
  MX4X1 top_core_KE_U5695 ( .A(top_core_KE_key_mem_4__115_), .B(
        top_core_KE_key_mem_5__115_), .C(top_core_KE_key_mem_6__115_), .D(
        top_core_KE_key_mem_7__115_), .S0(n4053), .S1(n3989), .Y(
        top_core_KE_n5628) );
  MX4X1 top_core_KE_U5079 ( .A(top_core_KE_key_mem_4__27_), .B(
        top_core_KE_key_mem_5__27_), .C(top_core_KE_key_mem_6__27_), .D(
        top_core_KE_key_mem_7__27_), .S0(n4049), .S1(n4001), .Y(
        top_core_KE_n5100) );
  MX4X1 top_core_KE_U5359 ( .A(top_core_KE_key_mem_4__67_), .B(
        top_core_KE_key_mem_5__67_), .C(top_core_KE_key_mem_6__67_), .D(
        top_core_KE_key_mem_7__67_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5340) );
  MX4X1 top_core_KE_U5639 ( .A(top_core_KE_key_mem_4__107_), .B(
        top_core_KE_key_mem_5__107_), .C(top_core_KE_key_mem_6__107_), .D(
        top_core_KE_key_mem_7__107_), .S0(n4107), .S1(n4005), .Y(
        top_core_KE_n5580) );
  MX4X1 top_core_KE_U5023 ( .A(top_core_KE_key_mem_4__19_), .B(
        top_core_KE_key_mem_5__19_), .C(top_core_KE_key_mem_6__19_), .D(
        top_core_KE_key_mem_7__19_), .S0(n4048), .S1(n3999), .Y(
        top_core_KE_n5052) );
  MX4X1 top_core_KE_U5303 ( .A(top_core_KE_key_mem_4__59_), .B(
        top_core_KE_key_mem_5__59_), .C(top_core_KE_key_mem_6__59_), .D(
        top_core_KE_key_mem_7__59_), .S0(n4040), .S1(n3993), .Y(
        top_core_KE_n5292) );
  MX4X1 top_core_KE_U5583 ( .A(top_core_KE_key_mem_4__99_), .B(
        top_core_KE_key_mem_5__99_), .C(top_core_KE_key_mem_6__99_), .D(
        top_core_KE_key_mem_7__99_), .S0(n4104), .S1(n4004), .Y(
        top_core_KE_n5532) );
  MX4X1 top_core_KE_U4911 ( .A(top_core_KE_key_mem_4__3_), .B(
        top_core_KE_key_mem_5__3_), .C(top_core_KE_key_mem_6__3_), .D(
        top_core_KE_key_mem_7__3_), .S0(n4044), .S1(n3996), .Y(
        top_core_KE_n4956) );
  MX4X1 top_core_KE_U5247 ( .A(top_core_KE_key_mem_4__51_), .B(
        top_core_KE_key_mem_5__51_), .C(top_core_KE_key_mem_6__51_), .D(
        top_core_KE_key_mem_7__51_), .S0(n4038), .S1(n3992), .Y(
        top_core_KE_n5244) );
  MX4X1 top_core_KE_U5471 ( .A(top_core_KE_key_mem_4__83_), .B(
        top_core_KE_key_mem_5__83_), .C(top_core_KE_key_mem_6__83_), .D(
        top_core_KE_key_mem_7__83_), .S0(n4056), .S1(n4011), .Y(
        top_core_KE_n5436) );
  MX4X1 top_core_KE_U5604 ( .A(top_core_KE_key_mem_4__102_), .B(
        top_core_KE_key_mem_5__102_), .C(top_core_KE_key_mem_6__102_), .D(
        top_core_KE_key_mem_7__102_), .S0(n4031), .S1(n4004), .Y(
        top_core_KE_n5550) );
  MX4X1 top_core_KE_U5156 ( .A(top_core_KE_key_mem_4__38_), .B(
        top_core_KE_key_mem_5__38_), .C(top_core_KE_key_mem_6__38_), .D(
        top_core_KE_key_mem_7__38_), .S0(n4035), .S1(n3989), .Y(
        top_core_KE_n5166) );
  MX4X1 top_core_KE_U5436 ( .A(top_core_KE_key_mem_4__78_), .B(
        top_core_KE_key_mem_5__78_), .C(top_core_KE_key_mem_6__78_), .D(
        top_core_KE_key_mem_7__78_), .S0(n4050), .S1(n4010), .Y(
        top_core_KE_n5406) );
  MX4X1 top_core_KE_U5100 ( .A(top_core_KE_key_mem_4__30_), .B(
        top_core_KE_key_mem_5__30_), .C(top_core_KE_key_mem_6__30_), .D(
        top_core_KE_key_mem_7__30_), .S0(n4050), .S1(n4001), .Y(
        top_core_KE_n5118) );
  MX4X1 top_core_KE_U5660 ( .A(top_core_KE_key_mem_4__110_), .B(
        top_core_KE_key_mem_5__110_), .C(top_core_KE_key_mem_6__110_), .D(
        top_core_KE_key_mem_7__110_), .S0(n4096), .S1(n4006), .Y(
        top_core_KE_n5598) );
  MX4X1 top_core_KE_U5324 ( .A(top_core_KE_key_mem_4__62_), .B(
        top_core_KE_key_mem_5__62_), .C(top_core_KE_key_mem_6__62_), .D(
        top_core_KE_key_mem_7__62_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5310) );
  MX4X1 top_core_KE_U5527 ( .A(top_core_KE_key_mem_4__91_), .B(
        top_core_KE_key_mem_5__91_), .C(top_core_KE_key_mem_6__91_), .D(
        top_core_KE_key_mem_7__91_), .S0(top_core_EC_n864), .S1(n4009), .Y(
        top_core_KE_n5484) );
  MX4X1 top_core_KE_U4967 ( .A(top_core_KE_key_mem_4__11_), .B(
        top_core_KE_key_mem_5__11_), .C(top_core_KE_key_mem_6__11_), .D(
        top_core_KE_key_mem_7__11_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5004) );
  MX4X1 top_core_KE_U5716 ( .A(top_core_KE_key_mem_4__118_), .B(
        top_core_KE_key_mem_5__118_), .C(top_core_KE_key_mem_6__118_), .D(
        top_core_KE_key_mem_7__118_), .S0(n4053), .S1(n4020), .Y(
        top_core_KE_n5646) );
  MX4X1 top_core_KE_U4932 ( .A(top_core_KE_key_mem_4__6_), .B(
        top_core_KE_key_mem_5__6_), .C(top_core_KE_key_mem_6__6_), .D(
        top_core_KE_key_mem_7__6_), .S0(n4044), .S1(n3997), .Y(
        top_core_KE_n4974) );
  MX4X1 top_core_KE_U5380 ( .A(top_core_KE_key_mem_4__70_), .B(
        top_core_KE_key_mem_5__70_), .C(top_core_KE_key_mem_6__70_), .D(
        top_core_KE_key_mem_7__70_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5358) );
  MX4X1 top_core_KE_U5751 ( .A(top_core_KE_key_mem_4__123_), .B(
        top_core_KE_key_mem_5__123_), .C(top_core_KE_key_mem_6__123_), .D(
        top_core_KE_key_mem_7__123_), .S0(n4055), .S1(n4007), .Y(
        top_core_KE_n5676) );
  MX4X1 top_core_KE_U5191 ( .A(top_core_KE_key_mem_4__43_), .B(
        top_core_KE_key_mem_5__43_), .C(top_core_KE_key_mem_6__43_), .D(
        top_core_KE_key_mem_7__43_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5196) );
  MX4X1 top_core_KE_U5044 ( .A(top_core_KE_key_mem_4__22_), .B(
        top_core_KE_key_mem_5__22_), .C(top_core_KE_key_mem_6__22_), .D(
        top_core_KE_key_mem_7__22_), .S0(n4048), .S1(n4000), .Y(
        top_core_KE_n5070) );
  MX4X1 top_core_KE_U5268 ( .A(top_core_KE_key_mem_4__54_), .B(
        top_core_KE_key_mem_5__54_), .C(top_core_KE_key_mem_6__54_), .D(
        top_core_KE_key_mem_7__54_), .S0(n4039), .S1(n3992), .Y(
        top_core_KE_n5262) );
  MX4X1 top_core_KE_U5702 ( .A(top_core_KE_key_mem_4__116_), .B(
        top_core_KE_key_mem_5__116_), .C(top_core_KE_key_mem_6__116_), .D(
        top_core_KE_key_mem_7__116_), .S0(n4053), .S1(n4020), .Y(
        top_core_KE_n5634) );
  MX4X1 top_core_KE_U5149 ( .A(top_core_KE_key_mem_4__37_), .B(
        top_core_KE_key_mem_5__37_), .C(top_core_KE_key_mem_6__37_), .D(
        top_core_KE_key_mem_7__37_), .S0(n4035), .S1(n3989), .Y(
        top_core_KE_n5160) );
  MX4X1 top_core_KE_U5590 ( .A(top_core_KE_key_mem_4__100_), .B(
        top_core_KE_key_mem_5__100_), .C(top_core_KE_key_mem_6__100_), .D(
        top_core_KE_key_mem_7__100_), .S0(n4109), .S1(n4004), .Y(
        top_core_KE_n5538) );
  MX4X1 top_core_KE_U5597 ( .A(top_core_KE_key_mem_4__101_), .B(
        top_core_KE_key_mem_5__101_), .C(top_core_KE_key_mem_6__101_), .D(
        top_core_KE_key_mem_7__101_), .S0(n4109), .S1(n4004), .Y(
        top_core_KE_n5544) );
  MX4X1 top_core_KE_U5366 ( .A(top_core_KE_key_mem_4__68_), .B(
        top_core_KE_key_mem_5__68_), .C(top_core_KE_key_mem_6__68_), .D(
        top_core_KE_key_mem_7__68_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5346) );
  MX4X1 top_core_KE_U5492 ( .A(top_core_KE_key_mem_4__86_), .B(
        top_core_KE_key_mem_5__86_), .C(top_core_KE_key_mem_6__86_), .D(
        top_core_KE_key_mem_7__86_), .S0(n4057), .S1(n4011), .Y(
        top_core_KE_n5454) );
  MX4X1 top_core_KE_U5142 ( .A(top_core_KE_key_mem_4__36_), .B(
        top_core_KE_key_mem_5__36_), .C(top_core_KE_key_mem_6__36_), .D(
        top_core_KE_key_mem_7__36_), .S0(n4051), .S1(n4003), .Y(
        top_core_KE_n5154) );
  MX4X1 top_core_KE_U5429 ( .A(top_core_KE_key_mem_4__77_), .B(
        top_core_KE_key_mem_5__77_), .C(top_core_KE_key_mem_6__77_), .D(
        top_core_KE_key_mem_7__77_), .S0(n4051), .S1(n4011), .Y(
        top_core_KE_n5400) );
  MX4X1 top_core_KE_U5422 ( .A(top_core_KE_key_mem_4__76_), .B(
        top_core_KE_key_mem_5__76_), .C(top_core_KE_key_mem_6__76_), .D(
        top_core_KE_key_mem_7__76_), .S0(n4040), .S1(n4011), .Y(
        top_core_KE_n5394) );
  MX4X1 top_core_KE_U5093 ( .A(top_core_KE_key_mem_4__29_), .B(
        top_core_KE_key_mem_5__29_), .C(top_core_KE_key_mem_6__29_), .D(
        top_core_KE_key_mem_7__29_), .S0(n4050), .S1(n4001), .Y(
        top_core_KE_n5112) );
  MX4X1 top_core_KE_U5086 ( .A(top_core_KE_key_mem_4__28_), .B(
        top_core_KE_key_mem_5__28_), .C(top_core_KE_key_mem_6__28_), .D(
        top_core_KE_key_mem_7__28_), .S0(n4050), .S1(n4001), .Y(
        top_core_KE_n5106) );
  MX4X1 top_core_KE_U5653 ( .A(top_core_KE_key_mem_4__109_), .B(
        top_core_KE_key_mem_5__109_), .C(top_core_KE_key_mem_6__109_), .D(
        top_core_KE_key_mem_7__109_), .S0(n4097), .S1(n4006), .Y(
        top_core_KE_n5592) );
  MX4X1 top_core_KE_U5646 ( .A(top_core_KE_key_mem_4__108_), .B(
        top_core_KE_key_mem_5__108_), .C(top_core_KE_key_mem_6__108_), .D(
        top_core_KE_key_mem_7__108_), .S0(n4107), .S1(n4005), .Y(
        top_core_KE_n5586) );
  MX4X1 top_core_KE_U5317 ( .A(top_core_KE_key_mem_4__61_), .B(
        top_core_KE_key_mem_5__61_), .C(top_core_KE_key_mem_6__61_), .D(
        top_core_KE_key_mem_7__61_), .S0(n4040), .S1(n3994), .Y(
        top_core_KE_n5304) );
  MX4X1 top_core_KE_U5310 ( .A(top_core_KE_key_mem_4__60_), .B(
        top_core_KE_key_mem_5__60_), .C(top_core_KE_key_mem_6__60_), .D(
        top_core_KE_key_mem_7__60_), .S0(n4040), .S1(n3993), .Y(
        top_core_KE_n5298) );
  MX4X1 top_core_KE_U5548 ( .A(top_core_KE_key_mem_4__94_), .B(
        top_core_KE_key_mem_5__94_), .C(top_core_KE_key_mem_6__94_), .D(
        top_core_KE_key_mem_7__94_), .S0(top_core_Addr[0]), .S1(n4003), .Y(
        top_core_KE_n5502) );
  MX4X1 top_core_KE_U4988 ( .A(top_core_KE_key_mem_4__14_), .B(
        top_core_KE_key_mem_5__14_), .C(top_core_KE_key_mem_6__14_), .D(
        top_core_KE_key_mem_7__14_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5022) );
  MX4X1 top_core_KE_U5709 ( .A(top_core_KE_key_mem_4__117_), .B(
        top_core_KE_key_mem_5__117_), .C(top_core_KE_key_mem_6__117_), .D(
        top_core_KE_key_mem_7__117_), .S0(n4053), .S1(n4020), .Y(
        top_core_KE_n5640) );
  MX4X1 top_core_KE_U5373 ( .A(top_core_KE_key_mem_4__69_), .B(
        top_core_KE_key_mem_5__69_), .C(top_core_KE_key_mem_6__69_), .D(
        top_core_KE_key_mem_7__69_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5352) );
  MX4X1 top_core_KE_U5212 ( .A(top_core_KE_key_mem_4__46_), .B(
        top_core_KE_key_mem_5__46_), .C(top_core_KE_key_mem_6__46_), .D(
        top_core_KE_key_mem_7__46_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5214) );
  MX4X1 top_core_KE_U5030 ( .A(top_core_KE_key_mem_4__20_), .B(
        top_core_KE_key_mem_5__20_), .C(top_core_KE_key_mem_6__20_), .D(
        top_core_KE_key_mem_7__20_), .S0(n4048), .S1(n4000), .Y(
        top_core_KE_n5058) );
  MX4X1 top_core_KE_U5037 ( .A(top_core_KE_key_mem_4__21_), .B(
        top_core_KE_key_mem_5__21_), .C(top_core_KE_key_mem_6__21_), .D(
        top_core_KE_key_mem_7__21_), .S0(n4048), .S1(n4000), .Y(
        top_core_KE_n5064) );
  MX4X1 top_core_KE_U4925 ( .A(top_core_KE_key_mem_4__5_), .B(
        top_core_KE_key_mem_5__5_), .C(top_core_KE_key_mem_6__5_), .D(
        top_core_KE_key_mem_7__5_), .S0(n4044), .S1(n3997), .Y(
        top_core_KE_n4968) );
  MX4X1 top_core_KE_U5254 ( .A(top_core_KE_key_mem_4__52_), .B(
        top_core_KE_key_mem_5__52_), .C(top_core_KE_key_mem_6__52_), .D(
        top_core_KE_key_mem_7__52_), .S0(n4038), .S1(n3992), .Y(
        top_core_KE_n5250) );
  MX4X1 top_core_KE_U5261 ( .A(top_core_KE_key_mem_4__53_), .B(
        top_core_KE_key_mem_5__53_), .C(top_core_KE_key_mem_6__53_), .D(
        top_core_KE_key_mem_7__53_), .S0(n4038), .S1(n3992), .Y(
        top_core_KE_n5256) );
  MX4X1 top_core_KE_U4918 ( .A(top_core_KE_key_mem_4__4_), .B(
        top_core_KE_key_mem_5__4_), .C(top_core_KE_key_mem_6__4_), .D(
        top_core_KE_key_mem_7__4_), .S0(n4044), .S1(n3997), .Y(
        top_core_KE_n4962) );
  MX4X1 top_core_KE_U5772 ( .A(top_core_KE_key_mem_4__126_), .B(
        top_core_KE_key_mem_5__126_), .C(top_core_KE_key_mem_6__126_), .D(
        top_core_KE_key_mem_7__126_), .S0(n4055), .S1(n4008), .Y(
        top_core_KE_n5694) );
  MX4X1 top_core_KE_U5688 ( .A(top_core_KE_key_mem_4__114_), .B(
        top_core_KE_key_mem_5__114_), .C(top_core_KE_key_mem_6__114_), .D(
        top_core_KE_key_mem_7__114_), .S0(n4052), .S1(n4020), .Y(
        top_core_KE_n5622) );
  MX4X1 top_core_KE_U5352 ( .A(top_core_KE_key_mem_4__66_), .B(
        top_core_KE_key_mem_5__66_), .C(top_core_KE_key_mem_6__66_), .D(
        top_core_KE_key_mem_7__66_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5334) );
  MX4X1 top_core_KE_U5478 ( .A(top_core_KE_key_mem_4__84_), .B(
        top_core_KE_key_mem_5__84_), .C(top_core_KE_key_mem_6__84_), .D(
        top_core_KE_key_mem_7__84_), .S0(n4056), .S1(n4012), .Y(
        top_core_KE_n5442) );
  MX4X1 top_core_KE_U5485 ( .A(top_core_KE_key_mem_4__85_), .B(
        top_core_KE_key_mem_5__85_), .C(top_core_KE_key_mem_6__85_), .D(
        top_core_KE_key_mem_7__85_), .S0(n4056), .S1(n4012), .Y(
        top_core_KE_n5448) );
  MX4X1 top_core_KE_U5016 ( .A(top_core_KE_key_mem_4__18_), .B(
        top_core_KE_key_mem_5__18_), .C(top_core_KE_key_mem_6__18_), .D(
        top_core_KE_key_mem_7__18_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5046) );
  MX4X1 top_core_KE_U5114 ( .A(top_core_KE_key_mem_4__32_), .B(
        top_core_KE_key_mem_5__32_), .C(top_core_KE_key_mem_6__32_), .D(
        top_core_KE_key_mem_7__32_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5130) );
  MX4X1 top_core_KE_U5394 ( .A(top_core_KE_key_mem_4__72_), .B(
        top_core_KE_key_mem_5__72_), .C(top_core_KE_key_mem_6__72_), .D(
        top_core_KE_key_mem_7__72_), .S0(n4043), .S1(n3996), .Y(
        top_core_KE_n5370) );
  MX4X1 top_core_KE_U5058 ( .A(top_core_KE_key_mem_4__24_), .B(
        top_core_KE_key_mem_5__24_), .C(top_core_KE_key_mem_6__24_), .D(
        top_core_KE_key_mem_7__24_), .S0(n4049), .S1(n4000), .Y(
        top_core_KE_n5082) );
  MX4X1 top_core_KE_U5618 ( .A(top_core_KE_key_mem_4__104_), .B(
        top_core_KE_key_mem_5__104_), .C(top_core_KE_key_mem_6__104_), .D(
        top_core_KE_key_mem_7__104_), .S0(n4101), .S1(n4005), .Y(
        top_core_KE_n5562) );
  MX4X1 top_core_KE_U5282 ( .A(top_core_KE_key_mem_4__56_), .B(
        top_core_KE_key_mem_5__56_), .C(top_core_KE_key_mem_6__56_), .D(
        top_core_KE_key_mem_7__56_), .S0(n4039), .S1(n3993), .Y(
        top_core_KE_n5274) );
  MX4X1 top_core_KE_U5562 ( .A(top_core_KE_key_mem_4__96_), .B(
        top_core_KE_key_mem_5__96_), .C(top_core_KE_key_mem_6__96_), .D(
        top_core_KE_key_mem_7__96_), .S0(n4100), .S1(n4003), .Y(
        top_core_KE_n5514) );
  MX4X1 top_core_KE_U5534 ( .A(top_core_KE_key_mem_4__92_), .B(
        top_core_KE_key_mem_5__92_), .C(top_core_KE_key_mem_6__92_), .D(
        top_core_KE_key_mem_7__92_), .S0(top_core_EC_n864), .S1(n4009), .Y(
        top_core_KE_n5490) );
  MX4X1 top_core_KE_U5541 ( .A(top_core_KE_key_mem_4__93_), .B(
        top_core_KE_key_mem_5__93_), .C(top_core_KE_key_mem_6__93_), .D(
        top_core_KE_key_mem_7__93_), .S0(n4052), .S1(n4003), .Y(
        top_core_KE_n5496) );
  MX4X1 top_core_KE_U4974 ( .A(top_core_KE_key_mem_4__12_), .B(
        top_core_KE_key_mem_5__12_), .C(top_core_KE_key_mem_6__12_), .D(
        top_core_KE_key_mem_7__12_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5010) );
  MX4X1 top_core_KE_U4981 ( .A(top_core_KE_key_mem_4__13_), .B(
        top_core_KE_key_mem_5__13_), .C(top_core_KE_key_mem_6__13_), .D(
        top_core_KE_key_mem_7__13_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5016) );
  MX4X1 top_core_KE_U5233 ( .A(top_core_KE_key_mem_4__49_), .B(
        top_core_KE_key_mem_5__49_), .C(top_core_KE_key_mem_6__49_), .D(
        top_core_KE_key_mem_7__49_), .S0(n4038), .S1(n3991), .Y(
        top_core_KE_n5232) );
  MX4X1 top_core_KE_U5226 ( .A(top_core_KE_key_mem_4__48_), .B(
        top_core_KE_key_mem_5__48_), .C(top_core_KE_key_mem_6__48_), .D(
        top_core_KE_key_mem_7__48_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5226) );
  MX4X1 top_core_KE_U5674 ( .A(top_core_KE_key_mem_4__112_), .B(
        top_core_KE_key_mem_5__112_), .C(top_core_KE_key_mem_6__112_), .D(
        top_core_KE_key_mem_7__112_), .S0(n4052), .S1(n4006), .Y(
        top_core_KE_n5610) );
  MX4X1 top_core_KE_U4890 ( .A(top_core_KE_key_mem_4__0_), .B(
        top_core_KE_key_mem_5__0_), .C(top_core_KE_key_mem_6__0_), .D(
        top_core_KE_key_mem_7__0_), .S0(n4047), .S1(n3996), .Y(
        top_core_KE_n4938) );
  MX4X1 top_core_KE_U5758 ( .A(top_core_KE_key_mem_4__124_), .B(
        top_core_KE_key_mem_5__124_), .C(top_core_KE_key_mem_6__124_), .D(
        top_core_KE_key_mem_7__124_), .S0(n4055), .S1(n4008), .Y(
        top_core_KE_n5682) );
  MX4X1 top_core_KE_U5765 ( .A(top_core_KE_key_mem_4__125_), .B(
        top_core_KE_key_mem_5__125_), .C(top_core_KE_key_mem_6__125_), .D(
        top_core_KE_key_mem_7__125_), .S0(n4055), .S1(n4008), .Y(
        top_core_KE_n5688) );
  MX4X1 top_core_KE_U5457 ( .A(top_core_KE_key_mem_4__81_), .B(
        top_core_KE_key_mem_5__81_), .C(top_core_KE_key_mem_6__81_), .D(
        top_core_KE_key_mem_7__81_), .S0(n4056), .S1(n4009), .Y(
        top_core_KE_n5424) );
  MX4X1 top_core_KE_U5338 ( .A(top_core_KE_key_mem_4__64_), .B(
        top_core_KE_key_mem_5__64_), .C(top_core_KE_key_mem_6__64_), .D(
        top_core_KE_key_mem_7__64_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5322) );
  MX4X1 top_core_KE_U5198 ( .A(top_core_KE_key_mem_4__44_), .B(
        top_core_KE_key_mem_5__44_), .C(top_core_KE_key_mem_6__44_), .D(
        top_core_KE_key_mem_7__44_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5202) );
  MX4X1 top_core_KE_U5205 ( .A(top_core_KE_key_mem_4__45_), .B(
        top_core_KE_key_mem_5__45_), .C(top_core_KE_key_mem_6__45_), .D(
        top_core_KE_key_mem_7__45_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5208) );
  MX4X1 top_core_KE_U5009 ( .A(top_core_KE_key_mem_4__17_), .B(
        top_core_KE_key_mem_5__17_), .C(top_core_KE_key_mem_6__17_), .D(
        top_core_KE_key_mem_7__17_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5040) );
  MX4X1 top_core_KE_U5450 ( .A(top_core_KE_key_mem_4__80_), .B(
        top_core_KE_key_mem_5__80_), .C(top_core_KE_key_mem_6__80_), .D(
        top_core_KE_key_mem_7__80_), .S0(n4035), .S1(n4009), .Y(
        top_core_KE_n5418) );
  MX4X1 top_core_KE_U5002 ( .A(top_core_KE_key_mem_4__16_), .B(
        top_core_KE_key_mem_5__16_), .C(top_core_KE_key_mem_6__16_), .D(
        top_core_KE_key_mem_7__16_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5034) );
  MX4X1 top_core_KE_U5569 ( .A(top_core_KE_key_mem_4__97_), .B(
        top_core_KE_key_mem_5__97_), .C(top_core_KE_key_mem_6__97_), .D(
        top_core_KE_key_mem_7__97_), .S0(n4031), .S1(n4003), .Y(
        top_core_KE_n5520) );
  MX4X1 top_core_KE_U5128 ( .A(top_core_KE_key_mem_4__34_), .B(
        top_core_KE_key_mem_5__34_), .C(top_core_KE_key_mem_6__34_), .D(
        top_core_KE_key_mem_7__34_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5142) );
  MX4X1 top_core_KE_U5401 ( .A(top_core_KE_key_mem_4__73_), .B(
        top_core_KE_key_mem_5__73_), .C(top_core_KE_key_mem_6__73_), .D(
        top_core_KE_key_mem_7__73_), .S0(n4057), .S1(n4009), .Y(
        top_core_KE_n5376) );
  MX4X1 top_core_KE_U5408 ( .A(top_core_KE_key_mem_4__74_), .B(
        top_core_KE_key_mem_5__74_), .C(top_core_KE_key_mem_6__74_), .D(
        top_core_KE_key_mem_7__74_), .S0(n4039), .S1(n4010), .Y(
        top_core_KE_n5382) );
  MX4X1 top_core_KE_U5065 ( .A(top_core_KE_key_mem_4__25_), .B(
        top_core_KE_key_mem_5__25_), .C(top_core_KE_key_mem_6__25_), .D(
        top_core_KE_key_mem_7__25_), .S0(n4049), .S1(n4000), .Y(
        top_core_KE_n5088) );
  MX4X1 top_core_KE_U5072 ( .A(top_core_KE_key_mem_4__26_), .B(
        top_core_KE_key_mem_5__26_), .C(top_core_KE_key_mem_6__26_), .D(
        top_core_KE_key_mem_7__26_), .S0(n4049), .S1(n4001), .Y(
        top_core_KE_n5094) );
  MX4X1 top_core_KE_U4897 ( .A(top_core_KE_key_mem_4__1_), .B(
        top_core_KE_key_mem_5__1_), .C(top_core_KE_key_mem_6__1_), .D(
        top_core_KE_key_mem_7__1_), .S0(n4043), .S1(n3996), .Y(
        top_core_KE_n4944) );
  MX4X1 top_core_KE_U5625 ( .A(top_core_KE_key_mem_4__105_), .B(
        top_core_KE_key_mem_5__105_), .C(top_core_KE_key_mem_6__105_), .D(
        top_core_KE_key_mem_7__105_), .S0(n4049), .S1(n4005), .Y(
        top_core_KE_n5568) );
  MX4X1 top_core_KE_U5632 ( .A(top_core_KE_key_mem_4__106_), .B(
        top_core_KE_key_mem_5__106_), .C(top_core_KE_key_mem_6__106_), .D(
        top_core_KE_key_mem_7__106_), .S0(n4100), .S1(n4005), .Y(
        top_core_KE_n5574) );
  MX4X1 top_core_KE_U5289 ( .A(top_core_KE_key_mem_4__57_), .B(
        top_core_KE_key_mem_5__57_), .C(top_core_KE_key_mem_6__57_), .D(
        top_core_KE_key_mem_7__57_), .S0(n4039), .S1(n3993), .Y(
        top_core_KE_n5280) );
  MX4X1 top_core_KE_U5296 ( .A(top_core_KE_key_mem_4__58_), .B(
        top_core_KE_key_mem_5__58_), .C(top_core_KE_key_mem_6__58_), .D(
        top_core_KE_key_mem_7__58_), .S0(n4040), .S1(n3993), .Y(
        top_core_KE_n5286) );
  MX4X1 top_core_KE_U5121 ( .A(top_core_KE_key_mem_4__33_), .B(
        top_core_KE_key_mem_5__33_), .C(top_core_KE_key_mem_6__33_), .D(
        top_core_KE_key_mem_7__33_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5136) );
  MX4X1 top_core_KE_U5576 ( .A(top_core_KE_key_mem_4__98_), .B(
        top_core_KE_key_mem_5__98_), .C(top_core_KE_key_mem_6__98_), .D(
        top_core_KE_key_mem_7__98_), .S0(n4108), .S1(n4004), .Y(
        top_core_KE_n5526) );
  MX4X1 top_core_KE_U5520 ( .A(top_core_KE_key_mem_4__90_), .B(
        top_core_KE_key_mem_5__90_), .C(top_core_KE_key_mem_6__90_), .D(
        top_core_KE_key_mem_7__90_), .S0(top_core_EC_n864), .S1(n4010), .Y(
        top_core_KE_n5478) );
  MX4X1 top_core_KE_U4960 ( .A(top_core_KE_key_mem_4__10_), .B(
        top_core_KE_key_mem_5__10_), .C(top_core_KE_key_mem_6__10_), .D(
        top_core_KE_key_mem_7__10_), .S0(n4045), .S1(n3998), .Y(
        top_core_KE_n4998) );
  MX4X1 top_core_KE_U5681 ( .A(top_core_KE_key_mem_4__113_), .B(
        top_core_KE_key_mem_5__113_), .C(top_core_KE_key_mem_6__113_), .D(
        top_core_KE_key_mem_7__113_), .S0(n4052), .S1(n4006), .Y(
        top_core_KE_n5616) );
  MX4X1 top_core_KE_U5184 ( .A(top_core_KE_key_mem_4__42_), .B(
        top_core_KE_key_mem_5__42_), .C(top_core_KE_key_mem_6__42_), .D(
        top_core_KE_key_mem_7__42_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5190) );
  MX4X1 top_core_KE_U5345 ( .A(top_core_KE_key_mem_4__65_), .B(
        top_core_KE_key_mem_5__65_), .C(top_core_KE_key_mem_6__65_), .D(
        top_core_KE_key_mem_7__65_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5328) );
  MX4X1 top_core_KE_U5744 ( .A(top_core_KE_key_mem_4__122_), .B(
        top_core_KE_key_mem_5__122_), .C(top_core_KE_key_mem_6__122_), .D(
        top_core_KE_key_mem_7__122_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5670) );
  MX4X1 top_core_KE_U4904 ( .A(top_core_KE_key_mem_4__2_), .B(
        top_core_KE_key_mem_5__2_), .C(top_core_KE_key_mem_6__2_), .D(
        top_core_KE_key_mem_7__2_), .S0(n4044), .S1(n3996), .Y(
        top_core_KE_n4950) );
  MX4X1 top_core_KE_U5506 ( .A(top_core_KE_key_mem_4__88_), .B(
        top_core_KE_key_mem_5__88_), .C(top_core_KE_key_mem_6__88_), .D(
        top_core_KE_key_mem_7__88_), .S0(n4057), .S1(n4010), .Y(
        top_core_KE_n5466) );
  MX4X1 top_core_KE_U4946 ( .A(top_core_KE_key_mem_4__8_), .B(
        top_core_KE_key_mem_5__8_), .C(top_core_KE_key_mem_6__8_), .D(
        top_core_KE_key_mem_7__8_), .S0(n4045), .S1(n3997), .Y(
        top_core_KE_n4986) );
  MX4X1 top_core_KE_U5240 ( .A(top_core_KE_key_mem_4__50_), .B(
        top_core_KE_key_mem_5__50_), .C(top_core_KE_key_mem_6__50_), .D(
        top_core_KE_key_mem_7__50_), .S0(n4038), .S1(n3991), .Y(
        top_core_KE_n5238) );
  MX4X1 top_core_KE_U5170 ( .A(top_core_KE_key_mem_4__40_), .B(
        top_core_KE_key_mem_5__40_), .C(top_core_KE_key_mem_6__40_), .D(
        top_core_KE_key_mem_7__40_), .S0(n4035), .S1(n3990), .Y(
        top_core_KE_n5178) );
  MX4X1 top_core_KE_U5513 ( .A(top_core_KE_key_mem_4__89_), .B(
        top_core_KE_key_mem_5__89_), .C(top_core_KE_key_mem_6__89_), .D(
        top_core_KE_key_mem_7__89_), .S0(top_core_EC_n864), .S1(n4010), .Y(
        top_core_KE_n5472) );
  MX4X1 top_core_KE_U4953 ( .A(top_core_KE_key_mem_4__9_), .B(
        top_core_KE_key_mem_5__9_), .C(top_core_KE_key_mem_6__9_), .D(
        top_core_KE_key_mem_7__9_), .S0(n4045), .S1(n3997), .Y(
        top_core_KE_n4992) );
  MX4X1 top_core_KE_U5177 ( .A(top_core_KE_key_mem_4__41_), .B(
        top_core_KE_key_mem_5__41_), .C(top_core_KE_key_mem_6__41_), .D(
        top_core_KE_key_mem_7__41_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5184) );
  MX4X1 top_core_KE_U5737 ( .A(top_core_KE_key_mem_4__121_), .B(
        top_core_KE_key_mem_5__121_), .C(top_core_KE_key_mem_6__121_), .D(
        top_core_KE_key_mem_7__121_), .S0(n4054), .S1(n4008), .Y(
        top_core_KE_n5664) );
  MX4X1 top_core_KE_U5464 ( .A(top_core_KE_key_mem_4__82_), .B(
        top_core_KE_key_mem_5__82_), .C(top_core_KE_key_mem_6__82_), .D(
        top_core_KE_key_mem_7__82_), .S0(n4056), .S1(n4010), .Y(
        top_core_KE_n5430) );
  MX4X1 top_core_KE_U5730 ( .A(top_core_KE_key_mem_4__120_), .B(
        top_core_KE_key_mem_5__120_), .C(top_core_KE_key_mem_6__120_), .D(
        top_core_KE_key_mem_7__120_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5658) );
  MX4X1 top_core_KE_U5780 ( .A(top_core_KE_key_mem_0__127_), .B(
        top_core_KE_key_mem_1__127_), .C(top_core_KE_key_mem_2__127_), .D(
        top_core_KE_key_mem_3__127_), .S0(n4038), .S1(n4008), .Y(
        top_core_KE_n5701) );
  MX4X1 top_core_KE_U5778 ( .A(top_core_KE_key_mem_8__127_), .B(
        top_core_KE_key_mem_9__127_), .C(top_core_KE_key_mem_10__127_), .D(
        top_core_KE_key_mem_11__127_), .S0(n4055), .S1(n4008), .Y(
        top_core_KE_n5699) );
  MX2X1 top_core_KE_U5777 ( .A(top_core_KE_n5696), .B(top_core_KE_n5697), .S0(
        n4015), .Y(top_core_KE_n5698) );
  MX4X1 top_core_KE_U5781 ( .A(top_core_KE_n5701), .B(top_core_KE_n5699), .C(
        top_core_KE_n5700), .D(top_core_KE_n5698), .S0(n3972), .S1(n3984), .Y(
        top_core_Key[127]) );
  MX4X1 top_core_KE_U5773 ( .A(top_core_KE_key_mem_0__126_), .B(
        top_core_KE_key_mem_1__126_), .C(top_core_KE_key_mem_2__126_), .D(
        top_core_KE_key_mem_3__126_), .S0(n4055), .S1(n4008), .Y(
        top_core_KE_n5695) );
  MX4X1 top_core_KE_U5771 ( .A(top_core_KE_key_mem_8__126_), .B(
        top_core_KE_key_mem_9__126_), .C(top_core_KE_key_mem_10__126_), .D(
        top_core_KE_key_mem_11__126_), .S0(n4055), .S1(n4008), .Y(
        top_core_KE_n5693) );
  MX2X1 top_core_KE_U5770 ( .A(top_core_KE_n5690), .B(top_core_KE_n5691), .S0(
        n4015), .Y(top_core_KE_n5692) );
  MX4X1 top_core_KE_U5774 ( .A(top_core_KE_n5695), .B(top_core_KE_n5693), .C(
        top_core_KE_n5694), .D(top_core_KE_n5692), .S0(n3972), .S1(n3984), .Y(
        top_core_Key[126]) );
  MX4X1 top_core_KE_U5759 ( .A(top_core_KE_key_mem_0__124_), .B(
        top_core_KE_key_mem_1__124_), .C(top_core_KE_key_mem_2__124_), .D(
        top_core_KE_key_mem_3__124_), .S0(n4055), .S1(n4008), .Y(
        top_core_KE_n5683) );
  MX4X1 top_core_KE_U5757 ( .A(top_core_KE_key_mem_8__124_), .B(
        top_core_KE_key_mem_9__124_), .C(top_core_KE_key_mem_10__124_), .D(
        top_core_KE_key_mem_11__124_), .S0(n4055), .S1(n4007), .Y(
        top_core_KE_n5681) );
  MX2X1 top_core_KE_U5756 ( .A(top_core_KE_n5678), .B(top_core_KE_n5679), .S0(
        n4014), .Y(top_core_KE_n5680) );
  MX4X1 top_core_KE_U5760 ( .A(top_core_KE_n5683), .B(top_core_KE_n5681), .C(
        top_core_KE_n5682), .D(top_core_KE_n5680), .S0(n3972), .S1(n3984), .Y(
        top_core_Key[124]) );
  MX4X1 top_core_KE_U5766 ( .A(top_core_KE_key_mem_0__125_), .B(
        top_core_KE_key_mem_1__125_), .C(top_core_KE_key_mem_2__125_), .D(
        top_core_KE_key_mem_3__125_), .S0(n4055), .S1(n4008), .Y(
        top_core_KE_n5689) );
  MX4X1 top_core_KE_U5764 ( .A(top_core_KE_key_mem_8__125_), .B(
        top_core_KE_key_mem_9__125_), .C(top_core_KE_key_mem_10__125_), .D(
        top_core_KE_key_mem_11__125_), .S0(n4055), .S1(n4008), .Y(
        top_core_KE_n5687) );
  MX2X1 top_core_KE_U5763 ( .A(top_core_KE_n5684), .B(top_core_KE_n5685), .S0(
        n4015), .Y(top_core_KE_n5686) );
  MX4X1 top_core_KE_U5767 ( .A(top_core_KE_n5689), .B(top_core_KE_n5687), .C(
        top_core_KE_n5688), .D(top_core_KE_n5686), .S0(n3972), .S1(n3984), .Y(
        top_core_Key[125]) );
  MX4X1 top_core_KE_U4940 ( .A(top_core_KE_key_mem_0__7_), .B(
        top_core_KE_key_mem_1__7_), .C(top_core_KE_key_mem_2__7_), .D(
        top_core_KE_key_mem_3__7_), .S0(n4045), .S1(n3997), .Y(
        top_core_KE_n4981) );
  MX4X1 top_core_KE_U4938 ( .A(top_core_KE_key_mem_8__7_), .B(
        top_core_KE_key_mem_9__7_), .C(top_core_KE_key_mem_10__7_), .D(
        top_core_KE_key_mem_11__7_), .S0(n4045), .S1(n3997), .Y(
        top_core_KE_n4979) );
  MX2X1 top_core_KE_U4937 ( .A(top_core_KE_n4976), .B(top_core_KE_n4977), .S0(
        n4014), .Y(top_core_KE_n4978) );
  MX4X1 top_core_KE_U4941 ( .A(top_core_KE_n4981), .B(top_core_KE_n4979), .C(
        top_core_KE_n4980), .D(top_core_KE_n4978), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[7]) );
  MX4X1 top_core_KE_U4912 ( .A(top_core_KE_key_mem_0__3_), .B(
        top_core_KE_key_mem_1__3_), .C(top_core_KE_key_mem_2__3_), .D(
        top_core_KE_key_mem_3__3_), .S0(n4044), .S1(n3996), .Y(
        top_core_KE_n4957) );
  MX4X1 top_core_KE_U4910 ( .A(top_core_KE_key_mem_8__3_), .B(
        top_core_KE_key_mem_9__3_), .C(top_core_KE_key_mem_10__3_), .D(
        top_core_KE_key_mem_11__3_), .S0(n4044), .S1(n3996), .Y(
        top_core_KE_n4955) );
  MX2X1 top_core_KE_U4909 ( .A(top_core_KE_n4952), .B(top_core_KE_n4953), .S0(
        n4015), .Y(top_core_KE_n4954) );
  MX4X1 top_core_KE_U4913 ( .A(top_core_KE_n4957), .B(top_core_KE_n4955), .C(
        top_core_KE_n4956), .D(top_core_KE_n4954), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[3]) );
  MX4X1 top_core_KE_U4968 ( .A(top_core_KE_key_mem_0__11_), .B(
        top_core_KE_key_mem_1__11_), .C(top_core_KE_key_mem_2__11_), .D(
        top_core_KE_key_mem_3__11_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5005) );
  MX4X1 top_core_KE_U4966 ( .A(top_core_KE_key_mem_8__11_), .B(
        top_core_KE_key_mem_9__11_), .C(top_core_KE_key_mem_10__11_), .D(
        top_core_KE_key_mem_11__11_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5003) );
  MX2X1 top_core_KE_U4965 ( .A(top_core_KE_n5000), .B(top_core_KE_n5001), .S0(
        n4013), .Y(top_core_KE_n5002) );
  MX4X1 top_core_KE_U4969 ( .A(top_core_KE_n5005), .B(top_core_KE_n5003), .C(
        top_core_KE_n5004), .D(top_core_KE_n5002), .S0(n3964), .S1(n3976), .Y(
        top_core_Key[11]) );
  MX4X1 top_core_KE_U4933 ( .A(top_core_KE_key_mem_0__6_), .B(
        top_core_KE_key_mem_1__6_), .C(top_core_KE_key_mem_2__6_), .D(
        top_core_KE_key_mem_3__6_), .S0(n4045), .S1(n3997), .Y(
        top_core_KE_n4975) );
  MX4X1 top_core_KE_U4931 ( .A(top_core_KE_key_mem_8__6_), .B(
        top_core_KE_key_mem_9__6_), .C(top_core_KE_key_mem_10__6_), .D(
        top_core_KE_key_mem_11__6_), .S0(n4044), .S1(n3997), .Y(
        top_core_KE_n4973) );
  MX2X1 top_core_KE_U4930 ( .A(top_core_KE_n4970), .B(top_core_KE_n4971), .S0(
        n4014), .Y(top_core_KE_n4972) );
  MX4X1 top_core_KE_U4934 ( .A(top_core_KE_n4975), .B(top_core_KE_n4973), .C(
        top_core_KE_n4974), .D(top_core_KE_n4972), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[6]) );
  MX4X1 top_core_KE_U4926 ( .A(top_core_KE_key_mem_0__5_), .B(
        top_core_KE_key_mem_1__5_), .C(top_core_KE_key_mem_2__5_), .D(
        top_core_KE_key_mem_3__5_), .S0(n4044), .S1(n3997), .Y(
        top_core_KE_n4969) );
  MX4X1 top_core_KE_U4924 ( .A(top_core_KE_key_mem_8__5_), .B(
        top_core_KE_key_mem_9__5_), .C(top_core_KE_key_mem_10__5_), .D(
        top_core_KE_key_mem_11__5_), .S0(n4044), .S1(n3997), .Y(
        top_core_KE_n4967) );
  MX2X1 top_core_KE_U4923 ( .A(top_core_KE_n4964), .B(top_core_KE_n4965), .S0(
        n4014), .Y(top_core_KE_n4966) );
  MX4X1 top_core_KE_U4927 ( .A(top_core_KE_n4969), .B(top_core_KE_n4967), .C(
        top_core_KE_n4968), .D(top_core_KE_n4966), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[5]) );
  MX4X1 top_core_KE_U4919 ( .A(top_core_KE_key_mem_0__4_), .B(
        top_core_KE_key_mem_1__4_), .C(top_core_KE_key_mem_2__4_), .D(
        top_core_KE_key_mem_3__4_), .S0(n4044), .S1(n3997), .Y(
        top_core_KE_n4963) );
  MX4X1 top_core_KE_U4917 ( .A(top_core_KE_key_mem_8__4_), .B(
        top_core_KE_key_mem_9__4_), .C(top_core_KE_key_mem_10__4_), .D(
        top_core_KE_key_mem_11__4_), .S0(n4044), .S1(n3996), .Y(
        top_core_KE_n4961) );
  MX2X1 top_core_KE_U4916 ( .A(top_core_KE_n4958), .B(top_core_KE_n4959), .S0(
        n4014), .Y(top_core_KE_n4960) );
  MX4X1 top_core_KE_U4920 ( .A(top_core_KE_n4963), .B(top_core_KE_n4961), .C(
        top_core_KE_n4962), .D(top_core_KE_n4960), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[4]) );
  MX4X1 top_core_KE_U4891 ( .A(top_core_KE_key_mem_0__0_), .B(
        top_core_KE_key_mem_1__0_), .C(top_core_KE_key_mem_2__0_), .D(
        top_core_KE_key_mem_3__0_), .S0(n4043), .S1(n3996), .Y(
        top_core_KE_n4939) );
  MX4X1 top_core_KE_U4889 ( .A(top_core_KE_key_mem_8__0_), .B(
        top_core_KE_key_mem_9__0_), .C(top_core_KE_key_mem_10__0_), .D(
        top_core_KE_key_mem_11__0_), .S0(n4035), .S1(n3999), .Y(
        top_core_KE_n4937) );
  MX2X1 top_core_KE_U4888 ( .A(top_core_KE_n4934), .B(top_core_KE_n4935), .S0(
        n4015), .Y(top_core_KE_n4936) );
  MX4X1 top_core_KE_U4892 ( .A(top_core_KE_n4939), .B(top_core_KE_n4937), .C(
        top_core_KE_n4938), .D(top_core_KE_n4936), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[0]) );
  MX4X1 top_core_KE_U4898 ( .A(top_core_KE_key_mem_0__1_), .B(
        top_core_KE_key_mem_1__1_), .C(top_core_KE_key_mem_2__1_), .D(
        top_core_KE_key_mem_3__1_), .S0(n4043), .S1(n3996), .Y(
        top_core_KE_n4945) );
  MX4X1 top_core_KE_U4896 ( .A(top_core_KE_key_mem_8__1_), .B(
        top_core_KE_key_mem_9__1_), .C(top_core_KE_key_mem_10__1_), .D(
        top_core_KE_key_mem_11__1_), .S0(n4043), .S1(n3996), .Y(
        top_core_KE_n4943) );
  MX2X1 top_core_KE_U4895 ( .A(top_core_KE_n4940), .B(top_core_KE_n4941), .S0(
        n4015), .Y(top_core_KE_n4942) );
  MX4X1 top_core_KE_U4899 ( .A(top_core_KE_n4945), .B(top_core_KE_n4943), .C(
        top_core_KE_n4944), .D(top_core_KE_n4942), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[1]) );
  MX4X1 top_core_KE_U4961 ( .A(top_core_KE_key_mem_0__10_), .B(
        top_core_KE_key_mem_1__10_), .C(top_core_KE_key_mem_2__10_), .D(
        top_core_KE_key_mem_3__10_), .S0(n4045), .S1(n3998), .Y(
        top_core_KE_n4999) );
  MX4X1 top_core_KE_U4959 ( .A(top_core_KE_key_mem_8__10_), .B(
        top_core_KE_key_mem_9__10_), .C(top_core_KE_key_mem_10__10_), .D(
        top_core_KE_key_mem_11__10_), .S0(n4045), .S1(n3998), .Y(
        top_core_KE_n4997) );
  MX2X1 top_core_KE_U4958 ( .A(top_core_KE_n4994), .B(top_core_KE_n4995), .S0(
        n4013), .Y(top_core_KE_n4996) );
  MX4X1 top_core_KE_U4962 ( .A(top_core_KE_n4999), .B(top_core_KE_n4997), .C(
        top_core_KE_n4998), .D(top_core_KE_n4996), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[10]) );
  MX4X1 top_core_KE_U4905 ( .A(top_core_KE_key_mem_0__2_), .B(
        top_core_KE_key_mem_1__2_), .C(top_core_KE_key_mem_2__2_), .D(
        top_core_KE_key_mem_3__2_), .S0(n4044), .S1(n3996), .Y(
        top_core_KE_n4951) );
  MX4X1 top_core_KE_U4903 ( .A(top_core_KE_key_mem_8__2_), .B(
        top_core_KE_key_mem_9__2_), .C(top_core_KE_key_mem_10__2_), .D(
        top_core_KE_key_mem_11__2_), .S0(n4043), .S1(n3996), .Y(
        top_core_KE_n4949) );
  MX2X1 top_core_KE_U4902 ( .A(top_core_KE_n4946), .B(top_core_KE_n4947), .S0(
        n4015), .Y(top_core_KE_n4948) );
  MX4X1 top_core_KE_U4906 ( .A(top_core_KE_n4951), .B(top_core_KE_n4949), .C(
        top_core_KE_n4950), .D(top_core_KE_n4948), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[2]) );
  MX4X1 top_core_KE_U4947 ( .A(top_core_KE_key_mem_0__8_), .B(
        top_core_KE_key_mem_1__8_), .C(top_core_KE_key_mem_2__8_), .D(
        top_core_KE_key_mem_3__8_), .S0(n4045), .S1(n3997), .Y(
        top_core_KE_n4987) );
  MX4X1 top_core_KE_U4945 ( .A(top_core_KE_key_mem_8__8_), .B(
        top_core_KE_key_mem_9__8_), .C(top_core_KE_key_mem_10__8_), .D(
        top_core_KE_key_mem_11__8_), .S0(n4045), .S1(n3997), .Y(
        top_core_KE_n4985) );
  MX2X1 top_core_KE_U4944 ( .A(top_core_KE_n4982), .B(top_core_KE_n4983), .S0(
        n4014), .Y(top_core_KE_n4984) );
  MX4X1 top_core_KE_U4948 ( .A(top_core_KE_n4987), .B(top_core_KE_n4985), .C(
        top_core_KE_n4986), .D(top_core_KE_n4984), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[8]) );
  MX4X1 top_core_KE_U4954 ( .A(top_core_KE_key_mem_0__9_), .B(
        top_core_KE_key_mem_1__9_), .C(top_core_KE_key_mem_2__9_), .D(
        top_core_KE_key_mem_3__9_), .S0(n4045), .S1(n3998), .Y(
        top_core_KE_n4993) );
  MX4X1 top_core_KE_U4952 ( .A(top_core_KE_key_mem_8__9_), .B(
        top_core_KE_key_mem_9__9_), .C(top_core_KE_key_mem_10__9_), .D(
        top_core_KE_key_mem_11__9_), .S0(n4045), .S1(n3997), .Y(
        top_core_KE_n4991) );
  MX2X1 top_core_KE_U4951 ( .A(top_core_KE_n4988), .B(top_core_KE_n4989), .S0(
        n4014), .Y(top_core_KE_n4990) );
  MX4X1 top_core_KE_U4955 ( .A(top_core_KE_n4993), .B(top_core_KE_n4991), .C(
        top_core_KE_n4992), .D(top_core_KE_n4990), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[9]) );
  MX4X1 top_core_KE_U5612 ( .A(top_core_KE_key_mem_0__103_), .B(
        top_core_KE_key_mem_1__103_), .C(top_core_KE_key_mem_2__103_), .D(
        top_core_KE_key_mem_3__103_), .S0(n4107), .S1(n4005), .Y(
        top_core_KE_n5557) );
  MX4X1 top_core_KE_U5610 ( .A(top_core_KE_key_mem_8__103_), .B(
        top_core_KE_key_mem_9__103_), .C(top_core_KE_key_mem_10__103_), .D(
        top_core_KE_key_mem_11__103_), .S0(n4044), .S1(n4004), .Y(
        top_core_KE_n5555) );
  MX2X1 top_core_KE_U5609 ( .A(top_core_KE_n5552), .B(top_core_KE_n5553), .S0(
        n4018), .Y(top_core_KE_n5554) );
  MX4X1 top_core_KE_U5613 ( .A(top_core_KE_n5557), .B(top_core_KE_n5555), .C(
        top_core_KE_n5556), .D(top_core_KE_n5554), .S0(n3971), .S1(n3982), .Y(
        top_core_Key[103]) );
  MX4X1 top_core_KE_U5164 ( .A(top_core_KE_key_mem_0__39_), .B(
        top_core_KE_key_mem_1__39_), .C(top_core_KE_key_mem_2__39_), .D(
        top_core_KE_key_mem_3__39_), .S0(n4035), .S1(n3989), .Y(
        top_core_KE_n5173) );
  MX4X1 top_core_KE_U5162 ( .A(top_core_KE_key_mem_8__39_), .B(
        top_core_KE_key_mem_9__39_), .C(top_core_KE_key_mem_10__39_), .D(
        top_core_KE_key_mem_11__39_), .S0(n4035), .S1(n3989), .Y(
        top_core_KE_n5171) );
  MX2X1 top_core_KE_U5161 ( .A(top_core_KE_n5168), .B(top_core_KE_n5169), .S0(
        n4019), .Y(top_core_KE_n5170) );
  MX4X1 top_core_KE_U5165 ( .A(top_core_KE_n5173), .B(top_core_KE_n5171), .C(
        top_core_KE_n5172), .D(top_core_KE_n5170), .S0(n3966), .S1(n3978), .Y(
        top_core_Key[39]) );
  MX4X1 top_core_KE_U5444 ( .A(top_core_KE_key_mem_0__79_), .B(
        top_core_KE_key_mem_1__79_), .C(top_core_KE_key_mem_2__79_), .D(
        top_core_KE_key_mem_3__79_), .S0(top_core_Addr[0]), .S1(n4010), .Y(
        top_core_KE_n5413) );
  MX4X1 top_core_KE_U5442 ( .A(top_core_KE_key_mem_8__79_), .B(
        top_core_KE_key_mem_9__79_), .C(top_core_KE_key_mem_10__79_), .D(
        top_core_KE_key_mem_11__79_), .S0(top_core_EC_n864), .S1(n4012), .Y(
        top_core_KE_n5411) );
  MX2X1 top_core_KE_U5441 ( .A(top_core_KE_n5408), .B(top_core_KE_n5409), .S0(
        n4013), .Y(top_core_KE_n5410) );
  MX4X1 top_core_KE_U5445 ( .A(top_core_KE_n5413), .B(top_core_KE_n5411), .C(
        top_core_KE_n5412), .D(top_core_KE_n5410), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[79]) );
  MX4X1 top_core_KE_U5276 ( .A(top_core_KE_key_mem_0__55_), .B(
        top_core_KE_key_mem_1__55_), .C(top_core_KE_key_mem_2__55_), .D(
        top_core_KE_key_mem_3__55_), .S0(n4039), .S1(n3993), .Y(
        top_core_KE_n5269) );
  MX4X1 top_core_KE_U5274 ( .A(top_core_KE_key_mem_8__55_), .B(
        top_core_KE_key_mem_9__55_), .C(top_core_KE_key_mem_10__55_), .D(
        top_core_KE_key_mem_11__55_), .S0(n4039), .S1(n3992), .Y(
        top_core_KE_n5267) );
  MX2X1 top_core_KE_U5273 ( .A(top_core_KE_n5264), .B(top_core_KE_n5265), .S0(
        n4017), .Y(top_core_KE_n5266) );
  MX4X1 top_core_KE_U5277 ( .A(top_core_KE_n5269), .B(top_core_KE_n5267), .C(
        top_core_KE_n5268), .D(top_core_KE_n5266), .S0(n3967), .S1(n3979), .Y(
        top_core_Key[55]) );
  MX4X1 top_core_KE_U5724 ( .A(top_core_KE_key_mem_0__119_), .B(
        top_core_KE_key_mem_1__119_), .C(top_core_KE_key_mem_2__119_), .D(
        top_core_KE_key_mem_3__119_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5653) );
  MX4X1 top_core_KE_U5722 ( .A(top_core_KE_key_mem_8__119_), .B(
        top_core_KE_key_mem_9__119_), .C(top_core_KE_key_mem_10__119_), .D(
        top_core_KE_key_mem_11__119_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5651) );
  MX2X1 top_core_KE_U5721 ( .A(top_core_KE_n5648), .B(top_core_KE_n5649), .S0(
        n4013), .Y(top_core_KE_n5650) );
  MX4X1 top_core_KE_U5725 ( .A(top_core_KE_n5653), .B(top_core_KE_n5651), .C(
        top_core_KE_n5652), .D(top_core_KE_n5650), .S0(n3972), .S1(n3983), .Y(
        top_core_Key[119]) );
  MX4X1 top_core_KE_U5108 ( .A(top_core_KE_key_mem_0__31_), .B(
        top_core_KE_key_mem_1__31_), .C(top_core_KE_key_mem_2__31_), .D(
        top_core_KE_key_mem_3__31_), .S0(n4050), .S1(n4002), .Y(
        top_core_KE_n5125) );
  MX4X1 top_core_KE_U5106 ( .A(top_core_KE_key_mem_8__31_), .B(
        top_core_KE_key_mem_9__31_), .C(top_core_KE_key_mem_10__31_), .D(
        top_core_KE_key_mem_11__31_), .S0(n4050), .S1(n4002), .Y(
        top_core_KE_n5123) );
  MX2X1 top_core_KE_U5105 ( .A(top_core_KE_n5120), .B(top_core_KE_n5121), .S0(
        n4018), .Y(top_core_KE_n5122) );
  MX4X1 top_core_KE_U5109 ( .A(top_core_KE_n5125), .B(top_core_KE_n5123), .C(
        top_core_KE_n5124), .D(top_core_KE_n5122), .S0(n3965), .S1(n3978), .Y(
        top_core_Key[31]) );
  MX4X1 top_core_KE_U5388 ( .A(top_core_KE_key_mem_0__71_), .B(
        top_core_KE_key_mem_1__71_), .C(top_core_KE_key_mem_2__71_), .D(
        top_core_KE_key_mem_3__71_), .S0(n4043), .S1(n3996), .Y(
        top_core_KE_n5365) );
  MX4X1 top_core_KE_U5386 ( .A(top_core_KE_key_mem_8__71_), .B(
        top_core_KE_key_mem_9__71_), .C(top_core_KE_key_mem_10__71_), .D(
        top_core_KE_key_mem_11__71_), .S0(n4043), .S1(n3995), .Y(
        top_core_KE_n5363) );
  MX2X1 top_core_KE_U5385 ( .A(top_core_KE_n5360), .B(top_core_KE_n5361), .S0(
        n4015), .Y(top_core_KE_n5362) );
  MX4X1 top_core_KE_U5389 ( .A(top_core_KE_n5365), .B(top_core_KE_n5363), .C(
        top_core_KE_n5364), .D(top_core_KE_n5362), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[71]) );
  MX4X1 top_core_KE_U5668 ( .A(top_core_KE_key_mem_0__111_), .B(
        top_core_KE_key_mem_1__111_), .C(top_core_KE_key_mem_2__111_), .D(
        top_core_KE_key_mem_3__111_), .S0(n4052), .S1(n4006), .Y(
        top_core_KE_n5605) );
  MX4X1 top_core_KE_U5666 ( .A(top_core_KE_key_mem_8__111_), .B(
        top_core_KE_key_mem_9__111_), .C(top_core_KE_key_mem_10__111_), .D(
        top_core_KE_key_mem_11__111_), .S0(n4052), .S1(n4006), .Y(
        top_core_KE_n5603) );
  MX2X1 top_core_KE_U5665 ( .A(top_core_KE_n5600), .B(top_core_KE_n5601), .S0(
        n4016), .Y(top_core_KE_n5602) );
  MX4X1 top_core_KE_U5669 ( .A(top_core_KE_n5605), .B(top_core_KE_n5603), .C(
        top_core_KE_n5604), .D(top_core_KE_n5602), .S0(n3971), .S1(n3983), .Y(
        top_core_Key[111]) );
  MX4X1 top_core_KE_U5500 ( .A(top_core_KE_key_mem_0__87_), .B(
        top_core_KE_key_mem_1__87_), .C(top_core_KE_key_mem_2__87_), .D(
        top_core_KE_key_mem_3__87_), .S0(n4057), .S1(n4011), .Y(
        top_core_KE_n5461) );
  MX4X1 top_core_KE_U5498 ( .A(top_core_KE_key_mem_8__87_), .B(
        top_core_KE_key_mem_9__87_), .C(top_core_KE_key_mem_10__87_), .D(
        top_core_KE_key_mem_11__87_), .S0(n4057), .S1(n4011), .Y(
        top_core_KE_n5459) );
  MX2X1 top_core_KE_U5497 ( .A(top_core_KE_n5456), .B(top_core_KE_n5457), .S0(
        n4018), .Y(top_core_KE_n5458) );
  MX4X1 top_core_KE_U5501 ( .A(top_core_KE_n5461), .B(top_core_KE_n5459), .C(
        top_core_KE_n5460), .D(top_core_KE_n5458), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[87]) );
  MX4X1 top_core_KE_U5052 ( .A(top_core_KE_key_mem_0__23_), .B(
        top_core_KE_key_mem_1__23_), .C(top_core_KE_key_mem_2__23_), .D(
        top_core_KE_key_mem_3__23_), .S0(n4049), .S1(n4000), .Y(
        top_core_KE_n5077) );
  MX4X1 top_core_KE_U5050 ( .A(top_core_KE_key_mem_8__23_), .B(
        top_core_KE_key_mem_9__23_), .C(top_core_KE_key_mem_10__23_), .D(
        top_core_KE_key_mem_11__23_), .S0(n4048), .S1(n4000), .Y(
        top_core_KE_n5075) );
  MX2X1 top_core_KE_U5049 ( .A(top_core_KE_n5072), .B(top_core_KE_n5073), .S0(
        n4016), .Y(top_core_KE_n5074) );
  MX4X1 top_core_KE_U5053 ( .A(top_core_KE_n5077), .B(top_core_KE_n5075), .C(
        top_core_KE_n5076), .D(top_core_KE_n5074), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[23]) );
  MX4X1 top_core_KE_U5332 ( .A(top_core_KE_key_mem_0__63_), .B(
        top_core_KE_key_mem_1__63_), .C(top_core_KE_key_mem_2__63_), .D(
        top_core_KE_key_mem_3__63_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5317) );
  MX4X1 top_core_KE_U5330 ( .A(top_core_KE_key_mem_8__63_), .B(
        top_core_KE_key_mem_9__63_), .C(top_core_KE_key_mem_10__63_), .D(
        top_core_KE_key_mem_11__63_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5315) );
  MX2X1 top_core_KE_U5329 ( .A(top_core_KE_n5312), .B(top_core_KE_n5313), .S0(
        n4013), .Y(top_core_KE_n5314) );
  MX4X1 top_core_KE_U5333 ( .A(top_core_KE_n5317), .B(top_core_KE_n5315), .C(
        top_core_KE_n5316), .D(top_core_KE_n5314), .S0(n3967), .S1(n3980), .Y(
        top_core_Key[63]) );
  MX4X1 top_core_KE_U5556 ( .A(top_core_KE_key_mem_0__95_), .B(
        top_core_KE_key_mem_1__95_), .C(top_core_KE_key_mem_2__95_), .D(
        top_core_KE_key_mem_3__95_), .S0(n4032), .S1(n4003), .Y(
        top_core_KE_n5509) );
  MX4X1 top_core_KE_U5554 ( .A(top_core_KE_key_mem_8__95_), .B(
        top_core_KE_key_mem_9__95_), .C(top_core_KE_key_mem_10__95_), .D(
        top_core_KE_key_mem_11__95_), .S0(n4100), .S1(n4003), .Y(
        top_core_KE_n5507) );
  MX2X1 top_core_KE_U5553 ( .A(top_core_KE_n5504), .B(top_core_KE_n5505), .S0(
        n4020), .Y(top_core_KE_n5506) );
  MX4X1 top_core_KE_U5557 ( .A(top_core_KE_n5509), .B(top_core_KE_n5507), .C(
        top_core_KE_n5508), .D(top_core_KE_n5506), .S0(n3970), .S1(n3982), .Y(
        top_core_Key[95]) );
  MX4X1 top_core_KE_U4996 ( .A(top_core_KE_key_mem_0__15_), .B(
        top_core_KE_key_mem_1__15_), .C(top_core_KE_key_mem_2__15_), .D(
        top_core_KE_key_mem_3__15_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5029) );
  MX4X1 top_core_KE_U4994 ( .A(top_core_KE_key_mem_8__15_), .B(
        top_core_KE_key_mem_9__15_), .C(top_core_KE_key_mem_10__15_), .D(
        top_core_KE_key_mem_11__15_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5027) );
  MX2X1 top_core_KE_U4993 ( .A(top_core_KE_n5024), .B(top_core_KE_n5025), .S0(
        n4012), .Y(top_core_KE_n5026) );
  MX4X1 top_core_KE_U4997 ( .A(top_core_KE_n5029), .B(top_core_KE_n5027), .C(
        top_core_KE_n5028), .D(top_core_KE_n5026), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[15]) );
  MX4X1 top_core_KE_U5220 ( .A(top_core_KE_key_mem_0__47_), .B(
        top_core_KE_key_mem_1__47_), .C(top_core_KE_key_mem_2__47_), .D(
        top_core_KE_key_mem_3__47_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5221) );
  MX4X1 top_core_KE_U5218 ( .A(top_core_KE_key_mem_8__47_), .B(
        top_core_KE_key_mem_9__47_), .C(top_core_KE_key_mem_10__47_), .D(
        top_core_KE_key_mem_11__47_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5219) );
  MX2X1 top_core_KE_U5217 ( .A(top_core_KE_n5216), .B(top_core_KE_n5217), .S0(
        n4020), .Y(top_core_KE_n5218) );
  MX4X1 top_core_KE_U5221 ( .A(top_core_KE_n5221), .B(top_core_KE_n5219), .C(
        top_core_KE_n5220), .D(top_core_KE_n5218), .S0(n3966), .S1(n3979), .Y(
        top_core_Key[47]) );
  MX4X1 top_core_KE_U5136 ( .A(top_core_KE_key_mem_0__35_), .B(
        top_core_KE_key_mem_1__35_), .C(top_core_KE_key_mem_2__35_), .D(
        top_core_KE_key_mem_3__35_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5149) );
  MX4X1 top_core_KE_U5134 ( .A(top_core_KE_key_mem_8__35_), .B(
        top_core_KE_key_mem_9__35_), .C(top_core_KE_key_mem_10__35_), .D(
        top_core_KE_key_mem_11__35_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5147) );
  MX2X1 top_core_KE_U5133 ( .A(top_core_KE_n5144), .B(top_core_KE_n5145), .S0(
        n4018), .Y(top_core_KE_n5146) );
  MX4X1 top_core_KE_U5137 ( .A(top_core_KE_n5149), .B(top_core_KE_n5147), .C(
        top_core_KE_n5148), .D(top_core_KE_n5146), .S0(n3965), .S1(n3978), .Y(
        top_core_Key[35]) );
  MX4X1 top_core_KE_U5416 ( .A(top_core_KE_key_mem_0__75_), .B(
        top_core_KE_key_mem_1__75_), .C(top_core_KE_key_mem_2__75_), .D(
        top_core_KE_key_mem_3__75_), .S0(n4036), .S1(n4011), .Y(
        top_core_KE_n5389) );
  MX4X1 top_core_KE_U5414 ( .A(top_core_KE_key_mem_8__75_), .B(
        top_core_KE_key_mem_9__75_), .C(top_core_KE_key_mem_10__75_), .D(
        top_core_KE_key_mem_11__75_), .S0(n4037), .S1(n4010), .Y(
        top_core_KE_n5387) );
  MX2X1 top_core_KE_U5413 ( .A(top_core_KE_n5384), .B(top_core_KE_n5385), .S0(
        n4015), .Y(top_core_KE_n5386) );
  MX4X1 top_core_KE_U5417 ( .A(top_core_KE_n5389), .B(top_core_KE_n5387), .C(
        top_core_KE_n5388), .D(top_core_KE_n5386), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[75]) );
  MX4X1 top_core_KE_U5696 ( .A(top_core_KE_key_mem_0__115_), .B(
        top_core_KE_key_mem_1__115_), .C(top_core_KE_key_mem_2__115_), .D(
        top_core_KE_key_mem_3__115_), .S0(n4053), .S1(n4030), .Y(
        top_core_KE_n5629) );
  MX4X1 top_core_KE_U5694 ( .A(top_core_KE_key_mem_8__115_), .B(
        top_core_KE_key_mem_9__115_), .C(top_core_KE_key_mem_10__115_), .D(
        top_core_KE_key_mem_11__115_), .S0(n4053), .S1(n4020), .Y(
        top_core_KE_n5627) );
  MX2X1 top_core_KE_U5693 ( .A(top_core_KE_n5624), .B(top_core_KE_n5625), .S0(
        n4013), .Y(top_core_KE_n5626) );
  MX4X1 top_core_KE_U5697 ( .A(top_core_KE_n5629), .B(top_core_KE_n5627), .C(
        top_core_KE_n5628), .D(top_core_KE_n5626), .S0(n3972), .S1(n3983), .Y(
        top_core_Key[115]) );
  MX4X1 top_core_KE_U5080 ( .A(top_core_KE_key_mem_0__27_), .B(
        top_core_KE_key_mem_1__27_), .C(top_core_KE_key_mem_2__27_), .D(
        top_core_KE_key_mem_3__27_), .S0(n4049), .S1(n4001), .Y(
        top_core_KE_n5101) );
  MX4X1 top_core_KE_U5078 ( .A(top_core_KE_key_mem_8__27_), .B(
        top_core_KE_key_mem_9__27_), .C(top_core_KE_key_mem_10__27_), .D(
        top_core_KE_key_mem_11__27_), .S0(n4049), .S1(n4001), .Y(
        top_core_KE_n5099) );
  MX2X1 top_core_KE_U5077 ( .A(top_core_KE_n5096), .B(top_core_KE_n5097), .S0(
        n4017), .Y(top_core_KE_n5098) );
  MX4X1 top_core_KE_U5081 ( .A(top_core_KE_n5101), .B(top_core_KE_n5099), .C(
        top_core_KE_n5100), .D(top_core_KE_n5098), .S0(n3965), .S1(n3977), .Y(
        top_core_Key[27]) );
  MX4X1 top_core_KE_U5360 ( .A(top_core_KE_key_mem_0__67_), .B(
        top_core_KE_key_mem_1__67_), .C(top_core_KE_key_mem_2__67_), .D(
        top_core_KE_key_mem_3__67_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5341) );
  MX4X1 top_core_KE_U5358 ( .A(top_core_KE_key_mem_8__67_), .B(
        top_core_KE_key_mem_9__67_), .C(top_core_KE_key_mem_10__67_), .D(
        top_core_KE_key_mem_11__67_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5339) );
  MX2X1 top_core_KE_U5357 ( .A(top_core_KE_n5336), .B(top_core_KE_n5337), .S0(
        n4014), .Y(top_core_KE_n5338) );
  MX4X1 top_core_KE_U5361 ( .A(top_core_KE_n5341), .B(top_core_KE_n5339), .C(
        top_core_KE_n5340), .D(top_core_KE_n5338), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[67]) );
  MX4X1 top_core_KE_U5640 ( .A(top_core_KE_key_mem_0__107_), .B(
        top_core_KE_key_mem_1__107_), .C(top_core_KE_key_mem_2__107_), .D(
        top_core_KE_key_mem_3__107_), .S0(n4105), .S1(n4005), .Y(
        top_core_KE_n5581) );
  MX4X1 top_core_KE_U5638 ( .A(top_core_KE_key_mem_8__107_), .B(
        top_core_KE_key_mem_9__107_), .C(top_core_KE_key_mem_10__107_), .D(
        top_core_KE_key_mem_11__107_), .S0(n4099), .S1(n4005), .Y(
        top_core_KE_n5579) );
  MX2X1 top_core_KE_U5637 ( .A(top_core_KE_n5576), .B(top_core_KE_n5577), .S0(
        n4017), .Y(top_core_KE_n5578) );
  MX4X1 top_core_KE_U5641 ( .A(top_core_KE_n5581), .B(top_core_KE_n5579), .C(
        top_core_KE_n5580), .D(top_core_KE_n5578), .S0(n3971), .S1(n3982), .Y(
        top_core_Key[107]) );
  MX4X1 top_core_KE_U5024 ( .A(top_core_KE_key_mem_0__19_), .B(
        top_core_KE_key_mem_1__19_), .C(top_core_KE_key_mem_2__19_), .D(
        top_core_KE_key_mem_3__19_), .S0(n4048), .S1(n3999), .Y(
        top_core_KE_n5053) );
  MX4X1 top_core_KE_U5022 ( .A(top_core_KE_key_mem_8__19_), .B(
        top_core_KE_key_mem_9__19_), .C(top_core_KE_key_mem_10__19_), .D(
        top_core_KE_key_mem_11__19_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5051) );
  MX2X1 top_core_KE_U5021 ( .A(top_core_KE_n5048), .B(top_core_KE_n5049), .S0(
        n4016), .Y(top_core_KE_n5050) );
  MX4X1 top_core_KE_U5025 ( .A(top_core_KE_n5053), .B(top_core_KE_n5051), .C(
        top_core_KE_n5052), .D(top_core_KE_n5050), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[19]) );
  MX4X1 top_core_KE_U5304 ( .A(top_core_KE_key_mem_0__59_), .B(
        top_core_KE_key_mem_1__59_), .C(top_core_KE_key_mem_2__59_), .D(
        top_core_KE_key_mem_3__59_), .S0(n4040), .S1(n3993), .Y(
        top_core_KE_n5293) );
  MX4X1 top_core_KE_U5302 ( .A(top_core_KE_key_mem_8__59_), .B(
        top_core_KE_key_mem_9__59_), .C(top_core_KE_key_mem_10__59_), .D(
        top_core_KE_key_mem_11__59_), .S0(n4040), .S1(n3993), .Y(
        top_core_KE_n5291) );
  MX2X1 top_core_KE_U5301 ( .A(top_core_KE_n5288), .B(top_core_KE_n5289), .S0(
        n4016), .Y(top_core_KE_n5290) );
  MX4X1 top_core_KE_U5305 ( .A(top_core_KE_n5293), .B(top_core_KE_n5291), .C(
        top_core_KE_n5292), .D(top_core_KE_n5290), .S0(n3967), .S1(n3979), .Y(
        top_core_Key[59]) );
  MX4X1 top_core_KE_U5584 ( .A(top_core_KE_key_mem_0__99_), .B(
        top_core_KE_key_mem_1__99_), .C(top_core_KE_key_mem_2__99_), .D(
        top_core_KE_key_mem_3__99_), .S0(n4110), .S1(n4004), .Y(
        top_core_KE_n5533) );
  MX4X1 top_core_KE_U5582 ( .A(top_core_KE_key_mem_8__99_), .B(
        top_core_KE_key_mem_9__99_), .C(top_core_KE_key_mem_10__99_), .D(
        top_core_KE_key_mem_11__99_), .S0(n4110), .S1(n4004), .Y(
        top_core_KE_n5531) );
  MX2X1 top_core_KE_U5581 ( .A(top_core_KE_n5528), .B(top_core_KE_n5529), .S0(
        n4019), .Y(top_core_KE_n5530) );
  MX4X1 top_core_KE_U5585 ( .A(top_core_KE_n5533), .B(top_core_KE_n5531), .C(
        top_core_KE_n5532), .D(top_core_KE_n5530), .S0(n3970), .S1(n3982), .Y(
        top_core_Key[99]) );
  MX4X1 top_core_KE_U5248 ( .A(top_core_KE_key_mem_0__51_), .B(
        top_core_KE_key_mem_1__51_), .C(top_core_KE_key_mem_2__51_), .D(
        top_core_KE_key_mem_3__51_), .S0(n4038), .S1(n3992), .Y(
        top_core_KE_n5245) );
  MX4X1 top_core_KE_U5246 ( .A(top_core_KE_key_mem_8__51_), .B(
        top_core_KE_key_mem_9__51_), .C(top_core_KE_key_mem_10__51_), .D(
        top_core_KE_key_mem_11__51_), .S0(n4038), .S1(n3992), .Y(
        top_core_KE_n5243) );
  MX2X1 top_core_KE_U5245 ( .A(top_core_KE_n5240), .B(top_core_KE_n5241), .S0(
        n4019), .Y(top_core_KE_n5242) );
  MX4X1 top_core_KE_U5249 ( .A(top_core_KE_n5245), .B(top_core_KE_n5243), .C(
        top_core_KE_n5244), .D(top_core_KE_n5242), .S0(n3967), .S1(n3979), .Y(
        top_core_Key[51]) );
  MX4X1 top_core_KE_U5472 ( .A(top_core_KE_key_mem_0__83_), .B(
        top_core_KE_key_mem_1__83_), .C(top_core_KE_key_mem_2__83_), .D(
        top_core_KE_key_mem_3__83_), .S0(n4056), .S1(n4011), .Y(
        top_core_KE_n5437) );
  MX4X1 top_core_KE_U5470 ( .A(top_core_KE_key_mem_8__83_), .B(
        top_core_KE_key_mem_9__83_), .C(top_core_KE_key_mem_10__83_), .D(
        top_core_KE_key_mem_11__83_), .S0(n4056), .S1(n4011), .Y(
        top_core_KE_n5435) );
  MX2X1 top_core_KE_U5469 ( .A(top_core_KE_n5432), .B(top_core_KE_n5433), .S0(
        n4016), .Y(top_core_KE_n5434) );
  MX4X1 top_core_KE_U5473 ( .A(top_core_KE_n5437), .B(top_core_KE_n5435), .C(
        top_core_KE_n5436), .D(top_core_KE_n5434), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[83]) );
  MX4X1 top_core_KE_U5605 ( .A(top_core_KE_key_mem_0__102_), .B(
        top_core_KE_key_mem_1__102_), .C(top_core_KE_key_mem_2__102_), .D(
        top_core_KE_key_mem_3__102_), .S0(n4048), .S1(n4004), .Y(
        top_core_KE_n5551) );
  MX4X1 top_core_KE_U5603 ( .A(top_core_KE_key_mem_8__102_), .B(
        top_core_KE_key_mem_9__102_), .C(top_core_KE_key_mem_10__102_), .D(
        top_core_KE_key_mem_11__102_), .S0(n4033), .S1(n4004), .Y(
        top_core_KE_n5549) );
  MX2X1 top_core_KE_U5602 ( .A(top_core_KE_n5546), .B(top_core_KE_n5547), .S0(
        n4018), .Y(top_core_KE_n5548) );
  MX4X1 top_core_KE_U5606 ( .A(top_core_KE_n5551), .B(top_core_KE_n5549), .C(
        top_core_KE_n5550), .D(top_core_KE_n5548), .S0(n3971), .S1(n3982), .Y(
        top_core_Key[102]) );
  MX4X1 top_core_KE_U5157 ( .A(top_core_KE_key_mem_0__38_), .B(
        top_core_KE_key_mem_1__38_), .C(top_core_KE_key_mem_2__38_), .D(
        top_core_KE_key_mem_3__38_), .S0(n4035), .S1(n3989), .Y(
        top_core_KE_n5167) );
  MX4X1 top_core_KE_U5155 ( .A(top_core_KE_key_mem_8__38_), .B(
        top_core_KE_key_mem_9__38_), .C(top_core_KE_key_mem_10__38_), .D(
        top_core_KE_key_mem_11__38_), .S0(n4035), .S1(n3989), .Y(
        top_core_KE_n5165) );
  MX2X1 top_core_KE_U5154 ( .A(top_core_KE_n5162), .B(top_core_KE_n5163), .S0(
        n4019), .Y(top_core_KE_n5164) );
  MX4X1 top_core_KE_U5158 ( .A(top_core_KE_n5167), .B(top_core_KE_n5165), .C(
        top_core_KE_n5166), .D(top_core_KE_n5164), .S0(n3966), .S1(n3978), .Y(
        top_core_Key[38]) );
  MX4X1 top_core_KE_U5437 ( .A(top_core_KE_key_mem_0__78_), .B(
        top_core_KE_key_mem_1__78_), .C(top_core_KE_key_mem_2__78_), .D(
        top_core_KE_key_mem_3__78_), .S0(n4099), .S1(n4011), .Y(
        top_core_KE_n5407) );
  MX4X1 top_core_KE_U5435 ( .A(top_core_KE_key_mem_8__78_), .B(
        top_core_KE_key_mem_9__78_), .C(top_core_KE_key_mem_10__78_), .D(
        top_core_KE_key_mem_11__78_), .S0(n4031), .S1(n4011), .Y(
        top_core_KE_n5405) );
  MX2X1 top_core_KE_U5434 ( .A(top_core_KE_n5402), .B(top_core_KE_n5403), .S0(
        n4013), .Y(top_core_KE_n5404) );
  MX4X1 top_core_KE_U5438 ( .A(top_core_KE_n5407), .B(top_core_KE_n5405), .C(
        top_core_KE_n5406), .D(top_core_KE_n5404), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[78]) );
  MX4X1 top_core_KE_U5101 ( .A(top_core_KE_key_mem_0__30_), .B(
        top_core_KE_key_mem_1__30_), .C(top_core_KE_key_mem_2__30_), .D(
        top_core_KE_key_mem_3__30_), .S0(n4050), .S1(n4001), .Y(
        top_core_KE_n5119) );
  MX4X1 top_core_KE_U5099 ( .A(top_core_KE_key_mem_8__30_), .B(
        top_core_KE_key_mem_9__30_), .C(top_core_KE_key_mem_10__30_), .D(
        top_core_KE_key_mem_11__30_), .S0(n4050), .S1(n4001), .Y(
        top_core_KE_n5117) );
  MX2X1 top_core_KE_U5098 ( .A(top_core_KE_n5114), .B(top_core_KE_n5115), .S0(
        n4018), .Y(top_core_KE_n5116) );
  MX4X1 top_core_KE_U5102 ( .A(top_core_KE_n5119), .B(top_core_KE_n5117), .C(
        top_core_KE_n5118), .D(top_core_KE_n5116), .S0(n3968), .S1(n3978), .Y(
        top_core_Key[30]) );
  MX4X1 top_core_KE_U5661 ( .A(top_core_KE_key_mem_0__110_), .B(
        top_core_KE_key_mem_1__110_), .C(top_core_KE_key_mem_2__110_), .D(
        top_core_KE_key_mem_3__110_), .S0(n4052), .S1(n4006), .Y(
        top_core_KE_n5599) );
  MX4X1 top_core_KE_U5659 ( .A(top_core_KE_key_mem_8__110_), .B(
        top_core_KE_key_mem_9__110_), .C(top_core_KE_key_mem_10__110_), .D(
        top_core_KE_key_mem_11__110_), .S0(n4109), .S1(n4006), .Y(
        top_core_KE_n5597) );
  MX2X1 top_core_KE_U5658 ( .A(top_core_KE_n5594), .B(top_core_KE_n5595), .S0(
        n4016), .Y(top_core_KE_n5596) );
  MX4X1 top_core_KE_U5662 ( .A(top_core_KE_n5599), .B(top_core_KE_n5597), .C(
        top_core_KE_n5598), .D(top_core_KE_n5596), .S0(n3971), .S1(n3983), .Y(
        top_core_Key[110]) );
  MX4X1 top_core_KE_U5325 ( .A(top_core_KE_key_mem_0__62_), .B(
        top_core_KE_key_mem_1__62_), .C(top_core_KE_key_mem_2__62_), .D(
        top_core_KE_key_mem_3__62_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5311) );
  MX4X1 top_core_KE_U5323 ( .A(top_core_KE_key_mem_8__62_), .B(
        top_core_KE_key_mem_9__62_), .C(top_core_KE_key_mem_10__62_), .D(
        top_core_KE_key_mem_11__62_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5309) );
  MX2X1 top_core_KE_U5322 ( .A(top_core_KE_n5306), .B(top_core_KE_n5307), .S0(
        n4012), .Y(top_core_KE_n5308) );
  MX4X1 top_core_KE_U5326 ( .A(top_core_KE_n5311), .B(top_core_KE_n5309), .C(
        top_core_KE_n5310), .D(top_core_KE_n5308), .S0(n3967), .S1(n3980), .Y(
        top_core_Key[62]) );
  MX4X1 top_core_KE_U5528 ( .A(top_core_KE_key_mem_0__91_), .B(
        top_core_KE_key_mem_1__91_), .C(top_core_KE_key_mem_2__91_), .D(
        top_core_KE_key_mem_3__91_), .S0(top_core_EC_n864), .S1(n4009), .Y(
        top_core_KE_n5485) );
  MX4X1 top_core_KE_U5526 ( .A(top_core_KE_key_mem_8__91_), .B(
        top_core_KE_key_mem_9__91_), .C(top_core_KE_key_mem_10__91_), .D(
        top_core_KE_key_mem_11__91_), .S0(n4057), .S1(n4009), .Y(
        top_core_KE_n5483) );
  MX2X1 top_core_KE_U5525 ( .A(top_core_KE_n5480), .B(top_core_KE_n5481), .S0(
        n4019), .Y(top_core_KE_n5482) );
  MX4X1 top_core_KE_U5529 ( .A(top_core_KE_n5485), .B(top_core_KE_n5483), .C(
        top_core_KE_n5484), .D(top_core_KE_n5482), .S0(n3970), .S1(n3981), .Y(
        top_core_Key[91]) );
  MX4X1 top_core_KE_U5717 ( .A(top_core_KE_key_mem_0__118_), .B(
        top_core_KE_key_mem_1__118_), .C(top_core_KE_key_mem_2__118_), .D(
        top_core_KE_key_mem_3__118_), .S0(n4053), .S1(n4029), .Y(
        top_core_KE_n5647) );
  MX4X1 top_core_KE_U5715 ( .A(top_core_KE_key_mem_8__118_), .B(
        top_core_KE_key_mem_9__118_), .C(top_core_KE_key_mem_10__118_), .D(
        top_core_KE_key_mem_11__118_), .S0(n4053), .S1(n3988), .Y(
        top_core_KE_n5645) );
  MX2X1 top_core_KE_U5714 ( .A(top_core_KE_n5642), .B(top_core_KE_n5643), .S0(
        n4013), .Y(top_core_KE_n5644) );
  MX4X1 top_core_KE_U5718 ( .A(top_core_KE_n5647), .B(top_core_KE_n5645), .C(
        top_core_KE_n5646), .D(top_core_KE_n5644), .S0(n3972), .S1(n3983), .Y(
        top_core_Key[118]) );
  MX4X1 top_core_KE_U5381 ( .A(top_core_KE_key_mem_0__70_), .B(
        top_core_KE_key_mem_1__70_), .C(top_core_KE_key_mem_2__70_), .D(
        top_core_KE_key_mem_3__70_), .S0(n4043), .S1(n3995), .Y(
        top_core_KE_n5359) );
  MX4X1 top_core_KE_U5379 ( .A(top_core_KE_key_mem_8__70_), .B(
        top_core_KE_key_mem_9__70_), .C(top_core_KE_key_mem_10__70_), .D(
        top_core_KE_key_mem_11__70_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5357) );
  MX2X1 top_core_KE_U5378 ( .A(top_core_KE_n5354), .B(top_core_KE_n5355), .S0(
        n4015), .Y(top_core_KE_n5356) );
  MX4X1 top_core_KE_U5382 ( .A(top_core_KE_n5359), .B(top_core_KE_n5357), .C(
        top_core_KE_n5358), .D(top_core_KE_n5356), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[70]) );
  MX4X1 top_core_KE_U5752 ( .A(top_core_KE_key_mem_0__123_), .B(
        top_core_KE_key_mem_1__123_), .C(top_core_KE_key_mem_2__123_), .D(
        top_core_KE_key_mem_3__123_), .S0(n4055), .S1(n4007), .Y(
        top_core_KE_n5677) );
  MX4X1 top_core_KE_U5750 ( .A(top_core_KE_key_mem_8__123_), .B(
        top_core_KE_key_mem_9__123_), .C(top_core_KE_key_mem_10__123_), .D(
        top_core_KE_key_mem_11__123_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5675) );
  MX2X1 top_core_KE_U5749 ( .A(top_core_KE_n5672), .B(top_core_KE_n5673), .S0(
        n4014), .Y(top_core_KE_n5674) );
  MX4X1 top_core_KE_U5753 ( .A(top_core_KE_n5677), .B(top_core_KE_n5675), .C(
        top_core_KE_n5676), .D(top_core_KE_n5674), .S0(n3972), .S1(n3983), .Y(
        top_core_Key[123]) );
  MX4X1 top_core_KE_U5192 ( .A(top_core_KE_key_mem_0__43_), .B(
        top_core_KE_key_mem_1__43_), .C(top_core_KE_key_mem_2__43_), .D(
        top_core_KE_key_mem_3__43_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5197) );
  MX4X1 top_core_KE_U5190 ( .A(top_core_KE_key_mem_8__43_), .B(
        top_core_KE_key_mem_9__43_), .C(top_core_KE_key_mem_10__43_), .D(
        top_core_KE_key_mem_11__43_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5195) );
  MX2X1 top_core_KE_U5189 ( .A(top_core_KE_n5192), .B(top_core_KE_n5193), .S0(
        n4020), .Y(top_core_KE_n5194) );
  MX4X1 top_core_KE_U5193 ( .A(top_core_KE_n5197), .B(top_core_KE_n5195), .C(
        top_core_KE_n5196), .D(top_core_KE_n5194), .S0(n3966), .S1(n3978), .Y(
        top_core_Key[43]) );
  MX4X1 top_core_KE_U5045 ( .A(top_core_KE_key_mem_0__22_), .B(
        top_core_KE_key_mem_1__22_), .C(top_core_KE_key_mem_2__22_), .D(
        top_core_KE_key_mem_3__22_), .S0(n4048), .S1(n4000), .Y(
        top_core_KE_n5071) );
  MX4X1 top_core_KE_U5043 ( .A(top_core_KE_key_mem_8__22_), .B(
        top_core_KE_key_mem_9__22_), .C(top_core_KE_key_mem_10__22_), .D(
        top_core_KE_key_mem_11__22_), .S0(n4048), .S1(n4000), .Y(
        top_core_KE_n5069) );
  MX2X1 top_core_KE_U5042 ( .A(top_core_KE_n5066), .B(top_core_KE_n5067), .S0(
        n4016), .Y(top_core_KE_n5068) );
  MX4X1 top_core_KE_U5046 ( .A(top_core_KE_n5071), .B(top_core_KE_n5069), .C(
        top_core_KE_n5070), .D(top_core_KE_n5068), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[22]) );
  MX4X1 top_core_KE_U5269 ( .A(top_core_KE_key_mem_0__54_), .B(
        top_core_KE_key_mem_1__54_), .C(top_core_KE_key_mem_2__54_), .D(
        top_core_KE_key_mem_3__54_), .S0(n4039), .S1(n3992), .Y(
        top_core_KE_n5263) );
  MX4X1 top_core_KE_U5267 ( .A(top_core_KE_key_mem_8__54_), .B(
        top_core_KE_key_mem_9__54_), .C(top_core_KE_key_mem_10__54_), .D(
        top_core_KE_key_mem_11__54_), .S0(n4039), .S1(n3992), .Y(
        top_core_KE_n5261) );
  MX2X1 top_core_KE_U5266 ( .A(top_core_KE_n5258), .B(top_core_KE_n5259), .S0(
        n4018), .Y(top_core_KE_n5260) );
  MX4X1 top_core_KE_U5270 ( .A(top_core_KE_n5263), .B(top_core_KE_n5261), .C(
        top_core_KE_n5262), .D(top_core_KE_n5260), .S0(n3967), .S1(n3979), .Y(
        top_core_Key[54]) );
  MX4X1 top_core_KE_U5703 ( .A(top_core_KE_key_mem_0__116_), .B(
        top_core_KE_key_mem_1__116_), .C(top_core_KE_key_mem_2__116_), .D(
        top_core_KE_key_mem_3__116_), .S0(n4053), .S1(top_core_Addr[1]), .Y(
        top_core_KE_n5635) );
  MX4X1 top_core_KE_U5701 ( .A(top_core_KE_key_mem_8__116_), .B(
        top_core_KE_key_mem_9__116_), .C(top_core_KE_key_mem_10__116_), .D(
        top_core_KE_key_mem_11__116_), .S0(n4053), .S1(n4030), .Y(
        top_core_KE_n5633) );
  MX2X1 top_core_KE_U5700 ( .A(top_core_KE_n5630), .B(top_core_KE_n5631), .S0(
        n4012), .Y(top_core_KE_n5632) );
  MX4X1 top_core_KE_U5704 ( .A(top_core_KE_n5635), .B(top_core_KE_n5633), .C(
        top_core_KE_n5634), .D(top_core_KE_n5632), .S0(n3972), .S1(n3983), .Y(
        top_core_Key[116]) );
  MX4X1 top_core_KE_U5150 ( .A(top_core_KE_key_mem_0__37_), .B(
        top_core_KE_key_mem_1__37_), .C(top_core_KE_key_mem_2__37_), .D(
        top_core_KE_key_mem_3__37_), .S0(n4035), .S1(n3989), .Y(
        top_core_KE_n5161) );
  MX4X1 top_core_KE_U5148 ( .A(top_core_KE_key_mem_8__37_), .B(
        top_core_KE_key_mem_9__37_), .C(top_core_KE_key_mem_10__37_), .D(
        top_core_KE_key_mem_11__37_), .S0(n4035), .S1(n3989), .Y(
        top_core_KE_n5159) );
  MX2X1 top_core_KE_U5147 ( .A(top_core_KE_n5156), .B(top_core_KE_n5157), .S0(
        n4019), .Y(top_core_KE_n5158) );
  MX4X1 top_core_KE_U5151 ( .A(top_core_KE_n5161), .B(top_core_KE_n5159), .C(
        top_core_KE_n5160), .D(top_core_KE_n5158), .S0(n3965), .S1(n3978), .Y(
        top_core_Key[37]) );
  MX4X1 top_core_KE_U5591 ( .A(top_core_KE_key_mem_0__100_), .B(
        top_core_KE_key_mem_1__100_), .C(top_core_KE_key_mem_2__100_), .D(
        top_core_KE_key_mem_3__100_), .S0(n4104), .S1(n4004), .Y(
        top_core_KE_n5539) );
  MX4X1 top_core_KE_U5589 ( .A(top_core_KE_key_mem_8__100_), .B(
        top_core_KE_key_mem_9__100_), .C(top_core_KE_key_mem_10__100_), .D(
        top_core_KE_key_mem_11__100_), .S0(n4098), .S1(n4004), .Y(
        top_core_KE_n5537) );
  MX2X1 top_core_KE_U5588 ( .A(top_core_KE_n5534), .B(top_core_KE_n5535), .S0(
        n4019), .Y(top_core_KE_n5536) );
  MX4X1 top_core_KE_U5592 ( .A(top_core_KE_n5539), .B(top_core_KE_n5537), .C(
        top_core_KE_n5538), .D(top_core_KE_n5536), .S0(n3970), .S1(n3982), .Y(
        top_core_Key[100]) );
  MX4X1 top_core_KE_U5598 ( .A(top_core_KE_key_mem_0__101_), .B(
        top_core_KE_key_mem_1__101_), .C(top_core_KE_key_mem_2__101_), .D(
        top_core_KE_key_mem_3__101_), .S0(n4101), .S1(n4004), .Y(
        top_core_KE_n5545) );
  MX4X1 top_core_KE_U5596 ( .A(top_core_KE_key_mem_8__101_), .B(
        top_core_KE_key_mem_9__101_), .C(top_core_KE_key_mem_10__101_), .D(
        top_core_KE_key_mem_11__101_), .S0(n4104), .S1(n4004), .Y(
        top_core_KE_n5543) );
  MX2X1 top_core_KE_U5595 ( .A(top_core_KE_n5540), .B(top_core_KE_n5541), .S0(
        n4018), .Y(top_core_KE_n5542) );
  MX4X1 top_core_KE_U5599 ( .A(top_core_KE_n5545), .B(top_core_KE_n5543), .C(
        top_core_KE_n5544), .D(top_core_KE_n5542), .S0(n3970), .S1(n3982), .Y(
        top_core_Key[101]) );
  MX4X1 top_core_KE_U5367 ( .A(top_core_KE_key_mem_0__68_), .B(
        top_core_KE_key_mem_1__68_), .C(top_core_KE_key_mem_2__68_), .D(
        top_core_KE_key_mem_3__68_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5347) );
  MX4X1 top_core_KE_U5365 ( .A(top_core_KE_key_mem_8__68_), .B(
        top_core_KE_key_mem_9__68_), .C(top_core_KE_key_mem_10__68_), .D(
        top_core_KE_key_mem_11__68_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5345) );
  MX2X1 top_core_KE_U5364 ( .A(top_core_KE_n5342), .B(top_core_KE_n5343), .S0(
        n4014), .Y(top_core_KE_n5344) );
  MX4X1 top_core_KE_U5368 ( .A(top_core_KE_n5347), .B(top_core_KE_n5345), .C(
        top_core_KE_n5346), .D(top_core_KE_n5344), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[68]) );
  MX4X1 top_core_KE_U5493 ( .A(top_core_KE_key_mem_0__86_), .B(
        top_core_KE_key_mem_1__86_), .C(top_core_KE_key_mem_2__86_), .D(
        top_core_KE_key_mem_3__86_), .S0(n4057), .S1(n4010), .Y(
        top_core_KE_n5455) );
  MX4X1 top_core_KE_U5491 ( .A(top_core_KE_key_mem_8__86_), .B(
        top_core_KE_key_mem_9__86_), .C(top_core_KE_key_mem_10__86_), .D(
        top_core_KE_key_mem_11__86_), .S0(n4057), .S1(n4012), .Y(
        top_core_KE_n5453) );
  MX2X1 top_core_KE_U5490 ( .A(top_core_KE_n5450), .B(top_core_KE_n5451), .S0(
        n4017), .Y(top_core_KE_n5452) );
  MX4X1 top_core_KE_U5494 ( .A(top_core_KE_n5455), .B(top_core_KE_n5453), .C(
        top_core_KE_n5454), .D(top_core_KE_n5452), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[86]) );
  MX4X1 top_core_KE_U5143 ( .A(top_core_KE_key_mem_0__36_), .B(
        top_core_KE_key_mem_1__36_), .C(top_core_KE_key_mem_2__36_), .D(
        top_core_KE_key_mem_3__36_), .S0(n4039), .S1(n3992), .Y(
        top_core_KE_n5155) );
  MX4X1 top_core_KE_U5141 ( .A(top_core_KE_key_mem_8__36_), .B(
        top_core_KE_key_mem_9__36_), .C(top_core_KE_key_mem_10__36_), .D(
        top_core_KE_key_mem_11__36_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5153) );
  MX2X1 top_core_KE_U5140 ( .A(top_core_KE_n5150), .B(top_core_KE_n5151), .S0(
        n4018), .Y(top_core_KE_n5152) );
  MX4X1 top_core_KE_U5144 ( .A(top_core_KE_n5155), .B(top_core_KE_n5153), .C(
        top_core_KE_n5154), .D(top_core_KE_n5152), .S0(n3965), .S1(n3978), .Y(
        top_core_Key[36]) );
  MX4X1 top_core_KE_U5430 ( .A(top_core_KE_key_mem_0__77_), .B(
        top_core_KE_key_mem_1__77_), .C(top_core_KE_key_mem_2__77_), .D(
        top_core_KE_key_mem_3__77_), .S0(n4108), .S1(n4012), .Y(
        top_core_KE_n5401) );
  MX4X1 top_core_KE_U5428 ( .A(top_core_KE_key_mem_8__77_), .B(
        top_core_KE_key_mem_9__77_), .C(top_core_KE_key_mem_10__77_), .D(
        top_core_KE_key_mem_11__77_), .S0(n4032), .S1(n4012), .Y(
        top_core_KE_n5399) );
  MX2X1 top_core_KE_U5427 ( .A(top_core_KE_n5396), .B(top_core_KE_n5397), .S0(
        n4014), .Y(top_core_KE_n5398) );
  MX4X1 top_core_KE_U5431 ( .A(top_core_KE_n5401), .B(top_core_KE_n5399), .C(
        top_core_KE_n5400), .D(top_core_KE_n5398), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[77]) );
  MX4X1 top_core_KE_U5423 ( .A(top_core_KE_key_mem_0__76_), .B(
        top_core_KE_key_mem_1__76_), .C(top_core_KE_key_mem_2__76_), .D(
        top_core_KE_key_mem_3__76_), .S0(n4103), .S1(n4011), .Y(
        top_core_KE_n5395) );
  MX4X1 top_core_KE_U5421 ( .A(top_core_KE_key_mem_8__76_), .B(
        top_core_KE_key_mem_9__76_), .C(top_core_KE_key_mem_10__76_), .D(
        top_core_KE_key_mem_11__76_), .S0(n4057), .S1(n4011), .Y(
        top_core_KE_n5393) );
  MX2X1 top_core_KE_U5420 ( .A(top_core_KE_n5390), .B(top_core_KE_n5391), .S0(
        n4014), .Y(top_core_KE_n5392) );
  MX4X1 top_core_KE_U5424 ( .A(top_core_KE_n5395), .B(top_core_KE_n5393), .C(
        top_core_KE_n5394), .D(top_core_KE_n5392), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[76]) );
  MX4X1 top_core_KE_U5094 ( .A(top_core_KE_key_mem_0__29_), .B(
        top_core_KE_key_mem_1__29_), .C(top_core_KE_key_mem_2__29_), .D(
        top_core_KE_key_mem_3__29_), .S0(n4050), .S1(n4001), .Y(
        top_core_KE_n5113) );
  MX4X1 top_core_KE_U5092 ( .A(top_core_KE_key_mem_8__29_), .B(
        top_core_KE_key_mem_9__29_), .C(top_core_KE_key_mem_10__29_), .D(
        top_core_KE_key_mem_11__29_), .S0(n4050), .S1(n4001), .Y(
        top_core_KE_n5111) );
  MX2X1 top_core_KE_U5091 ( .A(top_core_KE_n5108), .B(top_core_KE_n5109), .S0(
        n4017), .Y(top_core_KE_n5110) );
  MX4X1 top_core_KE_U5095 ( .A(top_core_KE_n5113), .B(top_core_KE_n5111), .C(
        top_core_KE_n5112), .D(top_core_KE_n5110), .S0(n3965), .S1(n3978), .Y(
        top_core_Key[29]) );
  MX4X1 top_core_KE_U5087 ( .A(top_core_KE_key_mem_0__28_), .B(
        top_core_KE_key_mem_1__28_), .C(top_core_KE_key_mem_2__28_), .D(
        top_core_KE_key_mem_3__28_), .S0(n4050), .S1(n4001), .Y(
        top_core_KE_n5107) );
  MX4X1 top_core_KE_U5085 ( .A(top_core_KE_key_mem_8__28_), .B(
        top_core_KE_key_mem_9__28_), .C(top_core_KE_key_mem_10__28_), .D(
        top_core_KE_key_mem_11__28_), .S0(n4050), .S1(n4001), .Y(
        top_core_KE_n5105) );
  MX2X1 top_core_KE_U5084 ( .A(top_core_KE_n5102), .B(top_core_KE_n5103), .S0(
        n4017), .Y(top_core_KE_n5104) );
  MX4X1 top_core_KE_U5088 ( .A(top_core_KE_n5107), .B(top_core_KE_n5105), .C(
        top_core_KE_n5106), .D(top_core_KE_n5104), .S0(n3965), .S1(n3980), .Y(
        top_core_Key[28]) );
  MX4X1 top_core_KE_U5654 ( .A(top_core_KE_key_mem_0__109_), .B(
        top_core_KE_key_mem_1__109_), .C(top_core_KE_key_mem_2__109_), .D(
        top_core_KE_key_mem_3__109_), .S0(n4108), .S1(n4006), .Y(
        top_core_KE_n5593) );
  MX4X1 top_core_KE_U5652 ( .A(top_core_KE_key_mem_8__109_), .B(
        top_core_KE_key_mem_9__109_), .C(top_core_KE_key_mem_10__109_), .D(
        top_core_KE_key_mem_11__109_), .S0(n4109), .S1(n4006), .Y(
        top_core_KE_n5591) );
  MX2X1 top_core_KE_U5651 ( .A(top_core_KE_n5588), .B(top_core_KE_n5589), .S0(
        n4017), .Y(top_core_KE_n5590) );
  MX4X1 top_core_KE_U5655 ( .A(top_core_KE_n5593), .B(top_core_KE_n5591), .C(
        top_core_KE_n5592), .D(top_core_KE_n5590), .S0(n3971), .S1(n3983), .Y(
        top_core_Key[109]) );
  MX4X1 top_core_KE_U5647 ( .A(top_core_KE_key_mem_0__108_), .B(
        top_core_KE_key_mem_1__108_), .C(top_core_KE_key_mem_2__108_), .D(
        top_core_KE_key_mem_3__108_), .S0(n4110), .S1(n4006), .Y(
        top_core_KE_n5587) );
  MX4X1 top_core_KE_U5645 ( .A(top_core_KE_key_mem_8__108_), .B(
        top_core_KE_key_mem_9__108_), .C(top_core_KE_key_mem_10__108_), .D(
        top_core_KE_key_mem_11__108_), .S0(n4110), .S1(n4005), .Y(
        top_core_KE_n5585) );
  MX2X1 top_core_KE_U5644 ( .A(top_core_KE_n5582), .B(top_core_KE_n5583), .S0(
        n4017), .Y(top_core_KE_n5584) );
  MX4X1 top_core_KE_U5648 ( .A(top_core_KE_n5587), .B(top_core_KE_n5585), .C(
        top_core_KE_n5586), .D(top_core_KE_n5584), .S0(n3971), .S1(n3983), .Y(
        top_core_Key[108]) );
  MX4X1 top_core_KE_U5318 ( .A(top_core_KE_key_mem_0__61_), .B(
        top_core_KE_key_mem_1__61_), .C(top_core_KE_key_mem_2__61_), .D(
        top_core_KE_key_mem_3__61_), .S0(n4040), .S1(n3994), .Y(
        top_core_KE_n5305) );
  MX4X1 top_core_KE_U5316 ( .A(top_core_KE_key_mem_8__61_), .B(
        top_core_KE_key_mem_9__61_), .C(top_core_KE_key_mem_10__61_), .D(
        top_core_KE_key_mem_11__61_), .S0(n4040), .S1(n3994), .Y(
        top_core_KE_n5303) );
  MX2X1 top_core_KE_U5315 ( .A(top_core_KE_n5300), .B(top_core_KE_n5301), .S0(
        n4016), .Y(top_core_KE_n5302) );
  MX4X1 top_core_KE_U5319 ( .A(top_core_KE_n5305), .B(top_core_KE_n5303), .C(
        top_core_KE_n5304), .D(top_core_KE_n5302), .S0(n3967), .S1(n3980), .Y(
        top_core_Key[61]) );
  MX4X1 top_core_KE_U5311 ( .A(top_core_KE_key_mem_0__60_), .B(
        top_core_KE_key_mem_1__60_), .C(top_core_KE_key_mem_2__60_), .D(
        top_core_KE_key_mem_3__60_), .S0(n4040), .S1(n3993), .Y(
        top_core_KE_n5299) );
  MX4X1 top_core_KE_U5309 ( .A(top_core_KE_key_mem_8__60_), .B(
        top_core_KE_key_mem_9__60_), .C(top_core_KE_key_mem_10__60_), .D(
        top_core_KE_key_mem_11__60_), .S0(n4040), .S1(n3993), .Y(
        top_core_KE_n5297) );
  MX2X1 top_core_KE_U5308 ( .A(top_core_KE_n5294), .B(top_core_KE_n5295), .S0(
        n4016), .Y(top_core_KE_n5296) );
  MX4X1 top_core_KE_U5312 ( .A(top_core_KE_n5299), .B(top_core_KE_n5297), .C(
        top_core_KE_n5298), .D(top_core_KE_n5296), .S0(n3967), .S1(n3979), .Y(
        top_core_Key[60]) );
  MX4X1 top_core_KE_U5549 ( .A(top_core_KE_key_mem_0__94_), .B(
        top_core_KE_key_mem_1__94_), .C(top_core_KE_key_mem_2__94_), .D(
        top_core_KE_key_mem_3__94_), .S0(n4103), .S1(n4003), .Y(
        top_core_KE_n5503) );
  MX4X1 top_core_KE_U5547 ( .A(top_core_KE_key_mem_8__94_), .B(
        top_core_KE_key_mem_9__94_), .C(top_core_KE_key_mem_10__94_), .D(
        top_core_KE_key_mem_11__94_), .S0(n4108), .S1(n4003), .Y(
        top_core_KE_n5501) );
  MX2X1 top_core_KE_U5546 ( .A(top_core_KE_n5498), .B(top_core_KE_n5499), .S0(
        n4020), .Y(top_core_KE_n5500) );
  MX4X1 top_core_KE_U5550 ( .A(top_core_KE_n5503), .B(top_core_KE_n5501), .C(
        top_core_KE_n5502), .D(top_core_KE_n5500), .S0(n3970), .S1(n3982), .Y(
        top_core_Key[94]) );
  MX4X1 top_core_KE_U4989 ( .A(top_core_KE_key_mem_0__14_), .B(
        top_core_KE_key_mem_1__14_), .C(top_core_KE_key_mem_2__14_), .D(
        top_core_KE_key_mem_3__14_), .S0(n4046), .S1(n4003), .Y(
        top_core_KE_n5023) );
  MX4X1 top_core_KE_U4987 ( .A(top_core_KE_key_mem_8__14_), .B(
        top_core_KE_key_mem_9__14_), .C(top_core_KE_key_mem_10__14_), .D(
        top_core_KE_key_mem_11__14_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5021) );
  MX2X1 top_core_KE_U4986 ( .A(top_core_KE_n5018), .B(top_core_KE_n5019), .S0(
        n4012), .Y(top_core_KE_n5020) );
  MX4X1 top_core_KE_U4990 ( .A(top_core_KE_n5023), .B(top_core_KE_n5021), .C(
        top_core_KE_n5022), .D(top_core_KE_n5020), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[14]) );
  MX4X1 top_core_KE_U5710 ( .A(top_core_KE_key_mem_0__117_), .B(
        top_core_KE_key_mem_1__117_), .C(top_core_KE_key_mem_2__117_), .D(
        top_core_KE_key_mem_3__117_), .S0(n4053), .S1(n4029), .Y(
        top_core_KE_n5641) );
  MX4X1 top_core_KE_U5708 ( .A(top_core_KE_key_mem_8__117_), .B(
        top_core_KE_key_mem_9__117_), .C(top_core_KE_key_mem_10__117_), .D(
        top_core_KE_key_mem_11__117_), .S0(n4053), .S1(n3988), .Y(
        top_core_KE_n5639) );
  MX2X1 top_core_KE_U5707 ( .A(top_core_KE_n5636), .B(top_core_KE_n5637), .S0(
        n4013), .Y(top_core_KE_n5638) );
  MX4X1 top_core_KE_U5711 ( .A(top_core_KE_n5641), .B(top_core_KE_n5639), .C(
        top_core_KE_n5640), .D(top_core_KE_n5638), .S0(n3972), .S1(n3983), .Y(
        top_core_Key[117]) );
  MX4X1 top_core_KE_U5374 ( .A(top_core_KE_key_mem_0__69_), .B(
        top_core_KE_key_mem_1__69_), .C(top_core_KE_key_mem_2__69_), .D(
        top_core_KE_key_mem_3__69_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5353) );
  MX4X1 top_core_KE_U5372 ( .A(top_core_KE_key_mem_8__69_), .B(
        top_core_KE_key_mem_9__69_), .C(top_core_KE_key_mem_10__69_), .D(
        top_core_KE_key_mem_11__69_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5351) );
  MX2X1 top_core_KE_U5371 ( .A(top_core_KE_n5348), .B(top_core_KE_n5349), .S0(
        n4014), .Y(top_core_KE_n5350) );
  MX4X1 top_core_KE_U5375 ( .A(top_core_KE_n5353), .B(top_core_KE_n5351), .C(
        top_core_KE_n5352), .D(top_core_KE_n5350), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[69]) );
  MX4X1 top_core_KE_U5213 ( .A(top_core_KE_key_mem_0__46_), .B(
        top_core_KE_key_mem_1__46_), .C(top_core_KE_key_mem_2__46_), .D(
        top_core_KE_key_mem_3__46_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5215) );
  MX4X1 top_core_KE_U5211 ( .A(top_core_KE_key_mem_8__46_), .B(
        top_core_KE_key_mem_9__46_), .C(top_core_KE_key_mem_10__46_), .D(
        top_core_KE_key_mem_11__46_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5213) );
  MX2X1 top_core_KE_U5210 ( .A(top_core_KE_n5210), .B(top_core_KE_n5211), .S0(
        n4020), .Y(top_core_KE_n5212) );
  MX4X1 top_core_KE_U5214 ( .A(top_core_KE_n5215), .B(top_core_KE_n5213), .C(
        top_core_KE_n5214), .D(top_core_KE_n5212), .S0(n3966), .S1(n3979), .Y(
        top_core_Key[46]) );
  MX4X1 top_core_KE_U5031 ( .A(top_core_KE_key_mem_0__20_), .B(
        top_core_KE_key_mem_1__20_), .C(top_core_KE_key_mem_2__20_), .D(
        top_core_KE_key_mem_3__20_), .S0(n4048), .S1(n4000), .Y(
        top_core_KE_n5059) );
  MX4X1 top_core_KE_U5029 ( .A(top_core_KE_key_mem_8__20_), .B(
        top_core_KE_key_mem_9__20_), .C(top_core_KE_key_mem_10__20_), .D(
        top_core_KE_key_mem_11__20_), .S0(n4048), .S1(n3999), .Y(
        top_core_KE_n5057) );
  MX2X1 top_core_KE_U5028 ( .A(top_core_KE_n5054), .B(top_core_KE_n5055), .S0(
        n4016), .Y(top_core_KE_n5056) );
  MX4X1 top_core_KE_U5032 ( .A(top_core_KE_n5059), .B(top_core_KE_n5057), .C(
        top_core_KE_n5058), .D(top_core_KE_n5056), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[20]) );
  MX4X1 top_core_KE_U5038 ( .A(top_core_KE_key_mem_0__21_), .B(
        top_core_KE_key_mem_1__21_), .C(top_core_KE_key_mem_2__21_), .D(
        top_core_KE_key_mem_3__21_), .S0(n4048), .S1(n4000), .Y(
        top_core_KE_n5065) );
  MX4X1 top_core_KE_U5036 ( .A(top_core_KE_key_mem_8__21_), .B(
        top_core_KE_key_mem_9__21_), .C(top_core_KE_key_mem_10__21_), .D(
        top_core_KE_key_mem_11__21_), .S0(n4048), .S1(n4000), .Y(
        top_core_KE_n5063) );
  MX2X1 top_core_KE_U5035 ( .A(top_core_KE_n5060), .B(top_core_KE_n5061), .S0(
        n4016), .Y(top_core_KE_n5062) );
  MX4X1 top_core_KE_U5039 ( .A(top_core_KE_n5065), .B(top_core_KE_n5063), .C(
        top_core_KE_n5064), .D(top_core_KE_n5062), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[21]) );
  MX4X1 top_core_KE_U5255 ( .A(top_core_KE_key_mem_0__52_), .B(
        top_core_KE_key_mem_1__52_), .C(top_core_KE_key_mem_2__52_), .D(
        top_core_KE_key_mem_3__52_), .S0(n4038), .S1(n3992), .Y(
        top_core_KE_n5251) );
  MX4X1 top_core_KE_U5253 ( .A(top_core_KE_key_mem_8__52_), .B(
        top_core_KE_key_mem_9__52_), .C(top_core_KE_key_mem_10__52_), .D(
        top_core_KE_key_mem_11__52_), .S0(n4038), .S1(n3992), .Y(
        top_core_KE_n5249) );
  MX2X1 top_core_KE_U5252 ( .A(top_core_KE_n5246), .B(top_core_KE_n5247), .S0(
        n4018), .Y(top_core_KE_n5248) );
  MX4X1 top_core_KE_U5256 ( .A(top_core_KE_n5251), .B(top_core_KE_n5249), .C(
        top_core_KE_n5250), .D(top_core_KE_n5248), .S0(n3967), .S1(n3979), .Y(
        top_core_Key[52]) );
  MX4X1 top_core_KE_U5262 ( .A(top_core_KE_key_mem_0__53_), .B(
        top_core_KE_key_mem_1__53_), .C(top_core_KE_key_mem_2__53_), .D(
        top_core_KE_key_mem_3__53_), .S0(n4039), .S1(n3992), .Y(
        top_core_KE_n5257) );
  MX4X1 top_core_KE_U5260 ( .A(top_core_KE_key_mem_8__53_), .B(
        top_core_KE_key_mem_9__53_), .C(top_core_KE_key_mem_10__53_), .D(
        top_core_KE_key_mem_11__53_), .S0(n4038), .S1(n3992), .Y(
        top_core_KE_n5255) );
  MX2X1 top_core_KE_U5259 ( .A(top_core_KE_n5252), .B(top_core_KE_n5253), .S0(
        n4018), .Y(top_core_KE_n5254) );
  MX4X1 top_core_KE_U5263 ( .A(top_core_KE_n5257), .B(top_core_KE_n5255), .C(
        top_core_KE_n5256), .D(top_core_KE_n5254), .S0(n3967), .S1(n3979), .Y(
        top_core_Key[53]) );
  MX4X1 top_core_KE_U5689 ( .A(top_core_KE_key_mem_0__114_), .B(
        top_core_KE_key_mem_1__114_), .C(top_core_KE_key_mem_2__114_), .D(
        top_core_KE_key_mem_3__114_), .S0(n4053), .S1(top_core_Addr[1]), .Y(
        top_core_KE_n5623) );
  MX4X1 top_core_KE_U5687 ( .A(top_core_KE_key_mem_8__114_), .B(
        top_core_KE_key_mem_9__114_), .C(top_core_KE_key_mem_10__114_), .D(
        top_core_KE_key_mem_11__114_), .S0(n4052), .S1(n4030), .Y(
        top_core_KE_n5621) );
  MX2X1 top_core_KE_U5686 ( .A(top_core_KE_n5618), .B(top_core_KE_n5619), .S0(
        n4015), .Y(top_core_KE_n5620) );
  MX4X1 top_core_KE_U5690 ( .A(top_core_KE_n5623), .B(top_core_KE_n5621), .C(
        top_core_KE_n5622), .D(top_core_KE_n5620), .S0(n3971), .S1(n3983), .Y(
        top_core_Key[114]) );
  MX4X1 top_core_KE_U5353 ( .A(top_core_KE_key_mem_0__66_), .B(
        top_core_KE_key_mem_1__66_), .C(top_core_KE_key_mem_2__66_), .D(
        top_core_KE_key_mem_3__66_), .S0(n4042), .S1(n3995), .Y(
        top_core_KE_n5335) );
  MX4X1 top_core_KE_U5351 ( .A(top_core_KE_key_mem_8__66_), .B(
        top_core_KE_key_mem_9__66_), .C(top_core_KE_key_mem_10__66_), .D(
        top_core_KE_key_mem_11__66_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5333) );
  MX2X1 top_core_KE_U5350 ( .A(top_core_KE_n5330), .B(top_core_KE_n5331), .S0(
        n4013), .Y(top_core_KE_n5332) );
  MX4X1 top_core_KE_U5354 ( .A(top_core_KE_n5335), .B(top_core_KE_n5333), .C(
        top_core_KE_n5334), .D(top_core_KE_n5332), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[66]) );
  MX4X1 top_core_KE_U5479 ( .A(top_core_KE_key_mem_0__84_), .B(
        top_core_KE_key_mem_1__84_), .C(top_core_KE_key_mem_2__84_), .D(
        top_core_KE_key_mem_3__84_), .S0(n4056), .S1(n4012), .Y(
        top_core_KE_n5443) );
  MX4X1 top_core_KE_U5477 ( .A(top_core_KE_key_mem_8__84_), .B(
        top_core_KE_key_mem_9__84_), .C(top_core_KE_key_mem_10__84_), .D(
        top_core_KE_key_mem_11__84_), .S0(n4056), .S1(n4011), .Y(
        top_core_KE_n5441) );
  MX2X1 top_core_KE_U5476 ( .A(top_core_KE_n5438), .B(top_core_KE_n5439), .S0(
        n4017), .Y(top_core_KE_n5440) );
  MX4X1 top_core_KE_U5480 ( .A(top_core_KE_n5443), .B(top_core_KE_n5441), .C(
        top_core_KE_n5442), .D(top_core_KE_n5440), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[84]) );
  MX4X1 top_core_KE_U5486 ( .A(top_core_KE_key_mem_0__85_), .B(
        top_core_KE_key_mem_1__85_), .C(top_core_KE_key_mem_2__85_), .D(
        top_core_KE_key_mem_3__85_), .S0(n4057), .S1(n4012), .Y(
        top_core_KE_n5449) );
  MX4X1 top_core_KE_U5484 ( .A(top_core_KE_key_mem_8__85_), .B(
        top_core_KE_key_mem_9__85_), .C(top_core_KE_key_mem_10__85_), .D(
        top_core_KE_key_mem_11__85_), .S0(n4056), .S1(n4012), .Y(
        top_core_KE_n5447) );
  MX2X1 top_core_KE_U5483 ( .A(top_core_KE_n5444), .B(top_core_KE_n5445), .S0(
        n4017), .Y(top_core_KE_n5446) );
  MX4X1 top_core_KE_U5487 ( .A(top_core_KE_n5449), .B(top_core_KE_n5447), .C(
        top_core_KE_n5448), .D(top_core_KE_n5446), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[85]) );
  MX4X1 top_core_KE_U5017 ( .A(top_core_KE_key_mem_0__18_), .B(
        top_core_KE_key_mem_1__18_), .C(top_core_KE_key_mem_2__18_), .D(
        top_core_KE_key_mem_3__18_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5047) );
  MX4X1 top_core_KE_U5015 ( .A(top_core_KE_key_mem_8__18_), .B(
        top_core_KE_key_mem_9__18_), .C(top_core_KE_key_mem_10__18_), .D(
        top_core_KE_key_mem_11__18_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5045) );
  MX2X1 top_core_KE_U5014 ( .A(top_core_KE_n5042), .B(top_core_KE_n5043), .S0(
        n4015), .Y(top_core_KE_n5044) );
  MX4X1 top_core_KE_U5018 ( .A(top_core_KE_n5047), .B(top_core_KE_n5045), .C(
        top_core_KE_n5046), .D(top_core_KE_n5044), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[18]) );
  MX4X1 top_core_KE_U5115 ( .A(top_core_KE_key_mem_0__32_), .B(
        top_core_KE_key_mem_1__32_), .C(top_core_KE_key_mem_2__32_), .D(
        top_core_KE_key_mem_3__32_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5131) );
  MX4X1 top_core_KE_U5113 ( .A(top_core_KE_key_mem_8__32_), .B(
        top_core_KE_key_mem_9__32_), .C(top_core_KE_key_mem_10__32_), .D(
        top_core_KE_key_mem_11__32_), .S0(n4050), .S1(n4002), .Y(
        top_core_KE_n5129) );
  MX2X1 top_core_KE_U5112 ( .A(top_core_KE_n5126), .B(top_core_KE_n5127), .S0(
        n4018), .Y(top_core_KE_n5128) );
  MX4X1 top_core_KE_U5116 ( .A(top_core_KE_n5131), .B(top_core_KE_n5129), .C(
        top_core_KE_n5130), .D(top_core_KE_n5128), .S0(n3965), .S1(n3978), .Y(
        top_core_Key[32]) );
  MX4X1 top_core_KE_U5395 ( .A(top_core_KE_key_mem_0__72_), .B(
        top_core_KE_key_mem_1__72_), .C(top_core_KE_key_mem_2__72_), .D(
        top_core_KE_key_mem_3__72_), .S0(n4043), .S1(n3996), .Y(
        top_core_KE_n5371) );
  MX4X1 top_core_KE_U5393 ( .A(top_core_KE_key_mem_8__72_), .B(
        top_core_KE_key_mem_9__72_), .C(top_core_KE_key_mem_10__72_), .D(
        top_core_KE_key_mem_11__72_), .S0(n4043), .S1(n3996), .Y(
        top_core_KE_n5369) );
  MX2X1 top_core_KE_U5392 ( .A(top_core_KE_n5366), .B(top_core_KE_n5367), .S0(
        n4015), .Y(top_core_KE_n5368) );
  MX4X1 top_core_KE_U5396 ( .A(top_core_KE_n5371), .B(top_core_KE_n5369), .C(
        top_core_KE_n5370), .D(top_core_KE_n5368), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[72]) );
  MX4X1 top_core_KE_U5059 ( .A(top_core_KE_key_mem_0__24_), .B(
        top_core_KE_key_mem_1__24_), .C(top_core_KE_key_mem_2__24_), .D(
        top_core_KE_key_mem_3__24_), .S0(n4049), .S1(n4000), .Y(
        top_core_KE_n5083) );
  MX4X1 top_core_KE_U5057 ( .A(top_core_KE_key_mem_8__24_), .B(
        top_core_KE_key_mem_9__24_), .C(top_core_KE_key_mem_10__24_), .D(
        top_core_KE_key_mem_11__24_), .S0(n4049), .S1(n4000), .Y(
        top_core_KE_n5081) );
  MX2X1 top_core_KE_U5056 ( .A(top_core_KE_n5078), .B(top_core_KE_n5079), .S0(
        n4016), .Y(top_core_KE_n5080) );
  MX4X1 top_core_KE_U5060 ( .A(top_core_KE_n5083), .B(top_core_KE_n5081), .C(
        top_core_KE_n5082), .D(top_core_KE_n5080), .S0(n3965), .S1(n3977), .Y(
        top_core_Key[24]) );
  MX4X1 top_core_KE_U5619 ( .A(top_core_KE_key_mem_0__104_), .B(
        top_core_KE_key_mem_1__104_), .C(top_core_KE_key_mem_2__104_), .D(
        top_core_KE_key_mem_3__104_), .S0(n4099), .S1(n4005), .Y(
        top_core_KE_n5563) );
  MX4X1 top_core_KE_U5617 ( .A(top_core_KE_key_mem_8__104_), .B(
        top_core_KE_key_mem_9__104_), .C(top_core_KE_key_mem_10__104_), .D(
        top_core_KE_key_mem_11__104_), .S0(top_core_Addr[0]), .S1(n4005), .Y(
        top_core_KE_n5561) );
  MX2X1 top_core_KE_U5616 ( .A(top_core_KE_n5558), .B(top_core_KE_n5559), .S0(
        n4018), .Y(top_core_KE_n5560) );
  MX4X1 top_core_KE_U5620 ( .A(top_core_KE_n5563), .B(top_core_KE_n5561), .C(
        top_core_KE_n5562), .D(top_core_KE_n5560), .S0(n3971), .S1(n3982), .Y(
        top_core_Key[104]) );
  MX4X1 top_core_KE_U5283 ( .A(top_core_KE_key_mem_0__56_), .B(
        top_core_KE_key_mem_1__56_), .C(top_core_KE_key_mem_2__56_), .D(
        top_core_KE_key_mem_3__56_), .S0(n4039), .S1(n3993), .Y(
        top_core_KE_n5275) );
  MX4X1 top_core_KE_U5281 ( .A(top_core_KE_key_mem_8__56_), .B(
        top_core_KE_key_mem_9__56_), .C(top_core_KE_key_mem_10__56_), .D(
        top_core_KE_key_mem_11__56_), .S0(n4039), .S1(n3993), .Y(
        top_core_KE_n5273) );
  MX2X1 top_core_KE_U5280 ( .A(top_core_KE_n5270), .B(top_core_KE_n5271), .S0(
        n4017), .Y(top_core_KE_n5272) );
  MX4X1 top_core_KE_U5284 ( .A(top_core_KE_n5275), .B(top_core_KE_n5273), .C(
        top_core_KE_n5274), .D(top_core_KE_n5272), .S0(n3967), .S1(n3979), .Y(
        top_core_Key[56]) );
  MX4X1 top_core_KE_U5563 ( .A(top_core_KE_key_mem_0__96_), .B(
        top_core_KE_key_mem_1__96_), .C(top_core_KE_key_mem_2__96_), .D(
        top_core_KE_key_mem_3__96_), .S0(n4106), .S1(n4003), .Y(
        top_core_KE_n5515) );
  MX4X1 top_core_KE_U5561 ( .A(top_core_KE_key_mem_8__96_), .B(
        top_core_KE_key_mem_9__96_), .C(top_core_KE_key_mem_10__96_), .D(
        top_core_KE_key_mem_11__96_), .S0(n4102), .S1(n4003), .Y(
        top_core_KE_n5513) );
  MX2X1 top_core_KE_U5560 ( .A(top_core_KE_n5510), .B(top_core_KE_n5511), .S0(
        n4019), .Y(top_core_KE_n5512) );
  MX4X1 top_core_KE_U5564 ( .A(top_core_KE_n5515), .B(top_core_KE_n5513), .C(
        top_core_KE_n5514), .D(top_core_KE_n5512), .S0(n3970), .S1(n3982), .Y(
        top_core_Key[96]) );
  MX4X1 top_core_KE_U5535 ( .A(top_core_KE_key_mem_0__92_), .B(
        top_core_KE_key_mem_1__92_), .C(top_core_KE_key_mem_2__92_), .D(
        top_core_KE_key_mem_3__92_), .S0(n4057), .S1(n4008), .Y(
        top_core_KE_n5491) );
  MX4X1 top_core_KE_U5533 ( .A(top_core_KE_key_mem_8__92_), .B(
        top_core_KE_key_mem_9__92_), .C(top_core_KE_key_mem_10__92_), .D(
        top_core_KE_key_mem_11__92_), .S0(top_core_EC_n864), .S1(n4009), .Y(
        top_core_KE_n5489) );
  MX2X1 top_core_KE_U5532 ( .A(top_core_KE_n5486), .B(top_core_KE_n5487), .S0(
        n4020), .Y(top_core_KE_n5488) );
  MX4X1 top_core_KE_U5536 ( .A(top_core_KE_n5491), .B(top_core_KE_n5489), .C(
        top_core_KE_n5490), .D(top_core_KE_n5488), .S0(n3970), .S1(n3982), .Y(
        top_core_Key[92]) );
  MX4X1 top_core_KE_U5542 ( .A(top_core_KE_key_mem_0__93_), .B(
        top_core_KE_key_mem_1__93_), .C(top_core_KE_key_mem_2__93_), .D(
        top_core_KE_key_mem_3__93_), .S0(n4105), .S1(n4003), .Y(
        top_core_KE_n5497) );
  MX4X1 top_core_KE_U5540 ( .A(top_core_KE_key_mem_8__93_), .B(
        top_core_KE_key_mem_9__93_), .C(top_core_KE_key_mem_10__93_), .D(
        top_core_KE_key_mem_11__93_), .S0(top_core_EC_n864), .S1(n4006), .Y(
        top_core_KE_n5495) );
  MX2X1 top_core_KE_U5539 ( .A(top_core_KE_n5492), .B(top_core_KE_n5493), .S0(
        n4012), .Y(top_core_KE_n5494) );
  MX4X1 top_core_KE_U5543 ( .A(top_core_KE_n5497), .B(top_core_KE_n5495), .C(
        top_core_KE_n5496), .D(top_core_KE_n5494), .S0(n3970), .S1(n3982), .Y(
        top_core_Key[93]) );
  MX4X1 top_core_KE_U4975 ( .A(top_core_KE_key_mem_0__12_), .B(
        top_core_KE_key_mem_1__12_), .C(top_core_KE_key_mem_2__12_), .D(
        top_core_KE_key_mem_3__12_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5011) );
  MX4X1 top_core_KE_U4973 ( .A(top_core_KE_key_mem_8__12_), .B(
        top_core_KE_key_mem_9__12_), .C(top_core_KE_key_mem_10__12_), .D(
        top_core_KE_key_mem_11__12_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5009) );
  MX2X1 top_core_KE_U4972 ( .A(top_core_KE_n5006), .B(top_core_KE_n5007), .S0(
        n4013), .Y(top_core_KE_n5008) );
  MX4X1 top_core_KE_U4976 ( .A(top_core_KE_n5011), .B(top_core_KE_n5009), .C(
        top_core_KE_n5010), .D(top_core_KE_n5008), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[12]) );
  MX4X1 top_core_KE_U4982 ( .A(top_core_KE_key_mem_0__13_), .B(
        top_core_KE_key_mem_1__13_), .C(top_core_KE_key_mem_2__13_), .D(
        top_core_KE_key_mem_3__13_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5017) );
  MX4X1 top_core_KE_U4980 ( .A(top_core_KE_key_mem_8__13_), .B(
        top_core_KE_key_mem_9__13_), .C(top_core_KE_key_mem_10__13_), .D(
        top_core_KE_key_mem_11__13_), .S0(n4046), .S1(n3998), .Y(
        top_core_KE_n5015) );
  MX2X1 top_core_KE_U4979 ( .A(top_core_KE_n5012), .B(top_core_KE_n5013), .S0(
        n4013), .Y(top_core_KE_n5014) );
  MX4X1 top_core_KE_U4983 ( .A(top_core_KE_n5017), .B(top_core_KE_n5015), .C(
        top_core_KE_n5016), .D(top_core_KE_n5014), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[13]) );
  MX4X1 top_core_KE_U5234 ( .A(top_core_KE_key_mem_0__49_), .B(
        top_core_KE_key_mem_1__49_), .C(top_core_KE_key_mem_2__49_), .D(
        top_core_KE_key_mem_3__49_), .S0(n4038), .S1(n3991), .Y(
        top_core_KE_n5233) );
  MX4X1 top_core_KE_U5232 ( .A(top_core_KE_key_mem_8__49_), .B(
        top_core_KE_key_mem_9__49_), .C(top_core_KE_key_mem_10__49_), .D(
        top_core_KE_key_mem_11__49_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5231) );
  MX2X1 top_core_KE_U5231 ( .A(top_core_KE_n5228), .B(top_core_KE_n5229), .S0(
        n4019), .Y(top_core_KE_n5230) );
  MX4X1 top_core_KE_U5235 ( .A(top_core_KE_n5233), .B(top_core_KE_n5231), .C(
        top_core_KE_n5232), .D(top_core_KE_n5230), .S0(n3966), .S1(n3979), .Y(
        top_core_Key[49]) );
  MX4X1 top_core_KE_U5227 ( .A(top_core_KE_key_mem_0__48_), .B(
        top_core_KE_key_mem_1__48_), .C(top_core_KE_key_mem_2__48_), .D(
        top_core_KE_key_mem_3__48_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5227) );
  MX4X1 top_core_KE_U5225 ( .A(top_core_KE_key_mem_8__48_), .B(
        top_core_KE_key_mem_9__48_), .C(top_core_KE_key_mem_10__48_), .D(
        top_core_KE_key_mem_11__48_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5225) );
  MX2X1 top_core_KE_U5224 ( .A(top_core_KE_n5222), .B(top_core_KE_n5223), .S0(
        n4020), .Y(top_core_KE_n5224) );
  MX4X1 top_core_KE_U5228 ( .A(top_core_KE_n5227), .B(top_core_KE_n5225), .C(
        top_core_KE_n5226), .D(top_core_KE_n5224), .S0(n3966), .S1(n3979), .Y(
        top_core_Key[48]) );
  MX4X1 top_core_KE_U5675 ( .A(top_core_KE_key_mem_0__112_), .B(
        top_core_KE_key_mem_1__112_), .C(top_core_KE_key_mem_2__112_), .D(
        top_core_KE_key_mem_3__112_), .S0(n4052), .S1(n4006), .Y(
        top_core_KE_n5611) );
  MX4X1 top_core_KE_U5673 ( .A(top_core_KE_key_mem_8__112_), .B(
        top_core_KE_key_mem_9__112_), .C(top_core_KE_key_mem_10__112_), .D(
        top_core_KE_key_mem_11__112_), .S0(n4052), .S1(n4006), .Y(
        top_core_KE_n5609) );
  MX2X1 top_core_KE_U5672 ( .A(top_core_KE_n5606), .B(top_core_KE_n5607), .S0(
        n4016), .Y(top_core_KE_n5608) );
  MX4X1 top_core_KE_U5676 ( .A(top_core_KE_n5611), .B(top_core_KE_n5609), .C(
        top_core_KE_n5610), .D(top_core_KE_n5608), .S0(n3971), .S1(n3983), .Y(
        top_core_Key[112]) );
  MX4X1 top_core_KE_U5458 ( .A(top_core_KE_key_mem_0__81_), .B(
        top_core_KE_key_mem_1__81_), .C(top_core_KE_key_mem_2__81_), .D(
        top_core_KE_key_mem_3__81_), .S0(n4056), .S1(n4009), .Y(
        top_core_KE_n5425) );
  MX4X1 top_core_KE_U5456 ( .A(top_core_KE_key_mem_8__81_), .B(
        top_core_KE_key_mem_9__81_), .C(top_core_KE_key_mem_10__81_), .D(
        top_core_KE_key_mem_11__81_), .S0(n4102), .S1(n4009), .Y(
        top_core_KE_n5423) );
  MX2X1 top_core_KE_U5455 ( .A(top_core_KE_n5420), .B(top_core_KE_n5421), .S0(
        n4013), .Y(top_core_KE_n5422) );
  MX4X1 top_core_KE_U5459 ( .A(top_core_KE_n5425), .B(top_core_KE_n5423), .C(
        top_core_KE_n5424), .D(top_core_KE_n5422), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[81]) );
  MX4X1 top_core_KE_U5339 ( .A(top_core_KE_key_mem_0__64_), .B(
        top_core_KE_key_mem_1__64_), .C(top_core_KE_key_mem_2__64_), .D(
        top_core_KE_key_mem_3__64_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5323) );
  MX4X1 top_core_KE_U5337 ( .A(top_core_KE_key_mem_8__64_), .B(
        top_core_KE_key_mem_9__64_), .C(top_core_KE_key_mem_10__64_), .D(
        top_core_KE_key_mem_11__64_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5321) );
  MX2X1 top_core_KE_U5336 ( .A(top_core_KE_n5318), .B(top_core_KE_n5319), .S0(
        n4013), .Y(top_core_KE_n5320) );
  MX4X1 top_core_KE_U5340 ( .A(top_core_KE_n5323), .B(top_core_KE_n5321), .C(
        top_core_KE_n5322), .D(top_core_KE_n5320), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[64]) );
  MX4X1 top_core_KE_U5199 ( .A(top_core_KE_key_mem_0__44_), .B(
        top_core_KE_key_mem_1__44_), .C(top_core_KE_key_mem_2__44_), .D(
        top_core_KE_key_mem_3__44_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5203) );
  MX4X1 top_core_KE_U5197 ( .A(top_core_KE_key_mem_8__44_), .B(
        top_core_KE_key_mem_9__44_), .C(top_core_KE_key_mem_10__44_), .D(
        top_core_KE_key_mem_11__44_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5201) );
  MX2X1 top_core_KE_U5196 ( .A(top_core_KE_n5198), .B(top_core_KE_n5199), .S0(
        n4020), .Y(top_core_KE_n5200) );
  MX4X1 top_core_KE_U5200 ( .A(top_core_KE_n5203), .B(top_core_KE_n5201), .C(
        top_core_KE_n5202), .D(top_core_KE_n5200), .S0(n3966), .S1(n3978), .Y(
        top_core_Key[44]) );
  MX4X1 top_core_KE_U5206 ( .A(top_core_KE_key_mem_0__45_), .B(
        top_core_KE_key_mem_1__45_), .C(top_core_KE_key_mem_2__45_), .D(
        top_core_KE_key_mem_3__45_), .S0(n4037), .S1(n3991), .Y(
        top_core_KE_n5209) );
  MX4X1 top_core_KE_U5204 ( .A(top_core_KE_key_mem_8__45_), .B(
        top_core_KE_key_mem_9__45_), .C(top_core_KE_key_mem_10__45_), .D(
        top_core_KE_key_mem_11__45_), .S0(n4037), .S1(n3990), .Y(
        top_core_KE_n5207) );
  MX2X1 top_core_KE_U5203 ( .A(top_core_KE_n5204), .B(top_core_KE_n5205), .S0(
        n4020), .Y(top_core_KE_n5206) );
  MX4X1 top_core_KE_U5207 ( .A(top_core_KE_n5209), .B(top_core_KE_n5207), .C(
        top_core_KE_n5208), .D(top_core_KE_n5206), .S0(n3966), .S1(n3979), .Y(
        top_core_Key[45]) );
  MX4X1 top_core_KE_U5010 ( .A(top_core_KE_key_mem_0__17_), .B(
        top_core_KE_key_mem_1__17_), .C(top_core_KE_key_mem_2__17_), .D(
        top_core_KE_key_mem_3__17_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5041) );
  MX4X1 top_core_KE_U5008 ( .A(top_core_KE_key_mem_8__17_), .B(
        top_core_KE_key_mem_9__17_), .C(top_core_KE_key_mem_10__17_), .D(
        top_core_KE_key_mem_11__17_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5039) );
  MX2X1 top_core_KE_U5007 ( .A(top_core_KE_n5036), .B(top_core_KE_n5037), .S0(
        n4012), .Y(top_core_KE_n5038) );
  MX4X1 top_core_KE_U5011 ( .A(top_core_KE_n5041), .B(top_core_KE_n5039), .C(
        top_core_KE_n5040), .D(top_core_KE_n5038), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[17]) );
  MX4X1 top_core_KE_U5451 ( .A(top_core_KE_key_mem_0__80_), .B(
        top_core_KE_key_mem_1__80_), .C(top_core_KE_key_mem_2__80_), .D(
        top_core_KE_key_mem_3__80_), .S0(n4106), .S1(n4009), .Y(
        top_core_KE_n5419) );
  MX4X1 top_core_KE_U5449 ( .A(top_core_KE_key_mem_8__80_), .B(
        top_core_KE_key_mem_9__80_), .C(top_core_KE_key_mem_10__80_), .D(
        top_core_KE_key_mem_11__80_), .S0(n4056), .S1(n4010), .Y(
        top_core_KE_n5417) );
  MX2X1 top_core_KE_U5448 ( .A(top_core_KE_n5414), .B(top_core_KE_n5415), .S0(
        n4013), .Y(top_core_KE_n5416) );
  MX4X1 top_core_KE_U5452 ( .A(top_core_KE_n5419), .B(top_core_KE_n5417), .C(
        top_core_KE_n5418), .D(top_core_KE_n5416), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[80]) );
  MX4X1 top_core_KE_U5003 ( .A(top_core_KE_key_mem_0__16_), .B(
        top_core_KE_key_mem_1__16_), .C(top_core_KE_key_mem_2__16_), .D(
        top_core_KE_key_mem_3__16_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5035) );
  MX4X1 top_core_KE_U5001 ( .A(top_core_KE_key_mem_8__16_), .B(
        top_core_KE_key_mem_9__16_), .C(top_core_KE_key_mem_10__16_), .D(
        top_core_KE_key_mem_11__16_), .S0(n4047), .S1(n3999), .Y(
        top_core_KE_n5033) );
  MX2X1 top_core_KE_U5000 ( .A(top_core_KE_n5030), .B(top_core_KE_n5031), .S0(
        n4012), .Y(top_core_KE_n5032) );
  MX4X1 top_core_KE_U5004 ( .A(top_core_KE_n5035), .B(top_core_KE_n5033), .C(
        top_core_KE_n5034), .D(top_core_KE_n5032), .S0(n3964), .S1(n3977), .Y(
        top_core_Key[16]) );
  MX4X1 top_core_KE_U5570 ( .A(top_core_KE_key_mem_0__97_), .B(
        top_core_KE_key_mem_1__97_), .C(top_core_KE_key_mem_2__97_), .D(
        top_core_KE_key_mem_3__97_), .S0(n4097), .S1(n4003), .Y(
        top_core_KE_n5521) );
  MX4X1 top_core_KE_U5568 ( .A(top_core_KE_key_mem_8__97_), .B(
        top_core_KE_key_mem_9__97_), .C(top_core_KE_key_mem_10__97_), .D(
        top_core_KE_key_mem_11__97_), .S0(n4098), .S1(n4003), .Y(
        top_core_KE_n5519) );
  MX2X1 top_core_KE_U5567 ( .A(top_core_KE_n5516), .B(top_core_KE_n5517), .S0(
        n4019), .Y(top_core_KE_n5518) );
  MX4X1 top_core_KE_U5571 ( .A(top_core_KE_n5521), .B(top_core_KE_n5519), .C(
        top_core_KE_n5520), .D(top_core_KE_n5518), .S0(n3970), .S1(n3982), .Y(
        top_core_Key[97]) );
  MX4X1 top_core_KE_U5129 ( .A(top_core_KE_key_mem_0__34_), .B(
        top_core_KE_key_mem_1__34_), .C(top_core_KE_key_mem_2__34_), .D(
        top_core_KE_key_mem_3__34_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5143) );
  MX4X1 top_core_KE_U5127 ( .A(top_core_KE_key_mem_8__34_), .B(
        top_core_KE_key_mem_9__34_), .C(top_core_KE_key_mem_10__34_), .D(
        top_core_KE_key_mem_11__34_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5141) );
  MX2X1 top_core_KE_U5126 ( .A(top_core_KE_n5138), .B(top_core_KE_n5139), .S0(
        n4018), .Y(top_core_KE_n5140) );
  MX4X1 top_core_KE_U5130 ( .A(top_core_KE_n5143), .B(top_core_KE_n5141), .C(
        top_core_KE_n5142), .D(top_core_KE_n5140), .S0(n3965), .S1(n3978), .Y(
        top_core_Key[34]) );
  MX4X1 top_core_KE_U5402 ( .A(top_core_KE_key_mem_0__73_), .B(
        top_core_KE_key_mem_1__73_), .C(top_core_KE_key_mem_2__73_), .D(
        top_core_KE_key_mem_3__73_), .S0(n4054), .S1(n4009), .Y(
        top_core_KE_n5377) );
  MX4X1 top_core_KE_U5400 ( .A(top_core_KE_key_mem_8__73_), .B(
        top_core_KE_key_mem_9__73_), .C(top_core_KE_key_mem_10__73_), .D(
        top_core_KE_key_mem_11__73_), .S0(n4043), .S1(n4008), .Y(
        top_core_KE_n5375) );
  MX2X1 top_core_KE_U5399 ( .A(top_core_KE_n5372), .B(top_core_KE_n5373), .S0(
        n4015), .Y(top_core_KE_n5374) );
  MX4X1 top_core_KE_U5403 ( .A(top_core_KE_n5377), .B(top_core_KE_n5375), .C(
        top_core_KE_n5376), .D(top_core_KE_n5374), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[73]) );
  MX4X1 top_core_KE_U5409 ( .A(top_core_KE_key_mem_0__74_), .B(
        top_core_KE_key_mem_1__74_), .C(top_core_KE_key_mem_2__74_), .D(
        top_core_KE_key_mem_3__74_), .S0(n4052), .S1(n4010), .Y(
        top_core_KE_n5383) );
  MX4X1 top_core_KE_U5407 ( .A(top_core_KE_key_mem_8__74_), .B(
        top_core_KE_key_mem_9__74_), .C(top_core_KE_key_mem_10__74_), .D(
        top_core_KE_key_mem_11__74_), .S0(n4055), .S1(n4009), .Y(
        top_core_KE_n5381) );
  MX2X1 top_core_KE_U5406 ( .A(top_core_KE_n5378), .B(top_core_KE_n5379), .S0(
        n4015), .Y(top_core_KE_n5380) );
  MX4X1 top_core_KE_U5410 ( .A(top_core_KE_n5383), .B(top_core_KE_n5381), .C(
        top_core_KE_n5382), .D(top_core_KE_n5380), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[74]) );
  MX4X1 top_core_KE_U5066 ( .A(top_core_KE_key_mem_0__25_), .B(
        top_core_KE_key_mem_1__25_), .C(top_core_KE_key_mem_2__25_), .D(
        top_core_KE_key_mem_3__25_), .S0(n4049), .S1(n4001), .Y(
        top_core_KE_n5089) );
  MX4X1 top_core_KE_U5064 ( .A(top_core_KE_key_mem_8__25_), .B(
        top_core_KE_key_mem_9__25_), .C(top_core_KE_key_mem_10__25_), .D(
        top_core_KE_key_mem_11__25_), .S0(n4049), .S1(n4000), .Y(
        top_core_KE_n5087) );
  MX2X1 top_core_KE_U5063 ( .A(top_core_KE_n5084), .B(top_core_KE_n5085), .S0(
        n4017), .Y(top_core_KE_n5086) );
  MX4X1 top_core_KE_U5067 ( .A(top_core_KE_n5089), .B(top_core_KE_n5087), .C(
        top_core_KE_n5088), .D(top_core_KE_n5086), .S0(n3965), .S1(n3977), .Y(
        top_core_Key[25]) );
  MX4X1 top_core_KE_U5073 ( .A(top_core_KE_key_mem_0__26_), .B(
        top_core_KE_key_mem_1__26_), .C(top_core_KE_key_mem_2__26_), .D(
        top_core_KE_key_mem_3__26_), .S0(n4049), .S1(n4001), .Y(
        top_core_KE_n5095) );
  MX4X1 top_core_KE_U5071 ( .A(top_core_KE_key_mem_8__26_), .B(
        top_core_KE_key_mem_9__26_), .C(top_core_KE_key_mem_10__26_), .D(
        top_core_KE_key_mem_11__26_), .S0(n4049), .S1(n4001), .Y(
        top_core_KE_n5093) );
  MX2X1 top_core_KE_U5070 ( .A(top_core_KE_n5090), .B(top_core_KE_n5091), .S0(
        n4017), .Y(top_core_KE_n5092) );
  MX4X1 top_core_KE_U5074 ( .A(top_core_KE_n5095), .B(top_core_KE_n5093), .C(
        top_core_KE_n5094), .D(top_core_KE_n5092), .S0(n3965), .S1(n3977), .Y(
        top_core_Key[26]) );
  MX4X1 top_core_KE_U5626 ( .A(top_core_KE_key_mem_0__105_), .B(
        top_core_KE_key_mem_1__105_), .C(top_core_KE_key_mem_2__105_), .D(
        top_core_KE_key_mem_3__105_), .S0(n4032), .S1(n4005), .Y(
        top_core_KE_n5569) );
  MX4X1 top_core_KE_U5624 ( .A(top_core_KE_key_mem_8__105_), .B(
        top_core_KE_key_mem_9__105_), .C(top_core_KE_key_mem_10__105_), .D(
        top_core_KE_key_mem_11__105_), .S0(n4031), .S1(n4005), .Y(
        top_core_KE_n5567) );
  MX2X1 top_core_KE_U5623 ( .A(top_core_KE_n5564), .B(top_core_KE_n5565), .S0(
        n4017), .Y(top_core_KE_n5566) );
  MX4X1 top_core_KE_U5627 ( .A(top_core_KE_n5569), .B(top_core_KE_n5567), .C(
        top_core_KE_n5568), .D(top_core_KE_n5566), .S0(n3971), .S1(n3982), .Y(
        top_core_Key[105]) );
  MX4X1 top_core_KE_U5633 ( .A(top_core_KE_key_mem_0__106_), .B(
        top_core_KE_key_mem_1__106_), .C(top_core_KE_key_mem_2__106_), .D(
        top_core_KE_key_mem_3__106_), .S0(n4101), .S1(n4005), .Y(
        top_core_KE_n5575) );
  MX4X1 top_core_KE_U5631 ( .A(top_core_KE_key_mem_8__106_), .B(
        top_core_KE_key_mem_9__106_), .C(top_core_KE_key_mem_10__106_), .D(
        top_core_KE_key_mem_11__106_), .S0(top_core_Addr[0]), .S1(n4005), .Y(
        top_core_KE_n5573) );
  MX2X1 top_core_KE_U5630 ( .A(top_core_KE_n5570), .B(top_core_KE_n5571), .S0(
        n4017), .Y(top_core_KE_n5572) );
  MX4X1 top_core_KE_U5634 ( .A(top_core_KE_n5575), .B(top_core_KE_n5573), .C(
        top_core_KE_n5574), .D(top_core_KE_n5572), .S0(n3971), .S1(n3982), .Y(
        top_core_Key[106]) );
  MX4X1 top_core_KE_U5290 ( .A(top_core_KE_key_mem_0__57_), .B(
        top_core_KE_key_mem_1__57_), .C(top_core_KE_key_mem_2__57_), .D(
        top_core_KE_key_mem_3__57_), .S0(n4040), .S1(n3993), .Y(
        top_core_KE_n5281) );
  MX4X1 top_core_KE_U5288 ( .A(top_core_KE_key_mem_8__57_), .B(
        top_core_KE_key_mem_9__57_), .C(top_core_KE_key_mem_10__57_), .D(
        top_core_KE_key_mem_11__57_), .S0(n4039), .S1(n3993), .Y(
        top_core_KE_n5279) );
  MX2X1 top_core_KE_U5287 ( .A(top_core_KE_n5276), .B(top_core_KE_n5277), .S0(
        n4017), .Y(top_core_KE_n5278) );
  MX4X1 top_core_KE_U5291 ( .A(top_core_KE_n5281), .B(top_core_KE_n5279), .C(
        top_core_KE_n5280), .D(top_core_KE_n5278), .S0(n3967), .S1(n3979), .Y(
        top_core_Key[57]) );
  MX4X1 top_core_KE_U5297 ( .A(top_core_KE_key_mem_0__58_), .B(
        top_core_KE_key_mem_1__58_), .C(top_core_KE_key_mem_2__58_), .D(
        top_core_KE_key_mem_3__58_), .S0(n4040), .S1(n3993), .Y(
        top_core_KE_n5287) );
  MX4X1 top_core_KE_U5295 ( .A(top_core_KE_key_mem_8__58_), .B(
        top_core_KE_key_mem_9__58_), .C(top_core_KE_key_mem_10__58_), .D(
        top_core_KE_key_mem_11__58_), .S0(n4040), .S1(n3993), .Y(
        top_core_KE_n5285) );
  MX2X1 top_core_KE_U5294 ( .A(top_core_KE_n5282), .B(top_core_KE_n5283), .S0(
        n4016), .Y(top_core_KE_n5284) );
  MX4X1 top_core_KE_U5298 ( .A(top_core_KE_n5287), .B(top_core_KE_n5285), .C(
        top_core_KE_n5286), .D(top_core_KE_n5284), .S0(n3967), .S1(n3979), .Y(
        top_core_Key[58]) );
  MX4X1 top_core_KE_U5122 ( .A(top_core_KE_key_mem_0__33_), .B(
        top_core_KE_key_mem_1__33_), .C(top_core_KE_key_mem_2__33_), .D(
        top_core_KE_key_mem_3__33_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5137) );
  MX4X1 top_core_KE_U5120 ( .A(top_core_KE_key_mem_8__33_), .B(
        top_core_KE_key_mem_9__33_), .C(top_core_KE_key_mem_10__33_), .D(
        top_core_KE_key_mem_11__33_), .S0(n4051), .S1(n4002), .Y(
        top_core_KE_n5135) );
  MX2X1 top_core_KE_U5119 ( .A(top_core_KE_n5132), .B(top_core_KE_n5133), .S0(
        n4018), .Y(top_core_KE_n5134) );
  MX4X1 top_core_KE_U5123 ( .A(top_core_KE_n5137), .B(top_core_KE_n5135), .C(
        top_core_KE_n5136), .D(top_core_KE_n5134), .S0(n3965), .S1(n3978), .Y(
        top_core_Key[33]) );
  MX4X1 top_core_KE_U5577 ( .A(top_core_KE_key_mem_0__98_), .B(
        top_core_KE_key_mem_1__98_), .C(top_core_KE_key_mem_2__98_), .D(
        top_core_KE_key_mem_3__98_), .S0(n4099), .S1(n4004), .Y(
        top_core_KE_n5527) );
  MX4X1 top_core_KE_U5575 ( .A(top_core_KE_key_mem_8__98_), .B(
        top_core_KE_key_mem_9__98_), .C(top_core_KE_key_mem_10__98_), .D(
        top_core_KE_key_mem_11__98_), .S0(n4043), .S1(n4004), .Y(
        top_core_KE_n5525) );
  MX2X1 top_core_KE_U5574 ( .A(top_core_KE_n5522), .B(top_core_KE_n5523), .S0(
        n4019), .Y(top_core_KE_n5524) );
  MX4X1 top_core_KE_U5578 ( .A(top_core_KE_n5527), .B(top_core_KE_n5525), .C(
        top_core_KE_n5526), .D(top_core_KE_n5524), .S0(n3970), .S1(n3982), .Y(
        top_core_Key[98]) );
  MX4X1 top_core_KE_U5521 ( .A(top_core_KE_key_mem_0__90_), .B(
        top_core_KE_key_mem_1__90_), .C(top_core_KE_key_mem_2__90_), .D(
        top_core_KE_key_mem_3__90_), .S0(top_core_EC_n864), .S1(n4009), .Y(
        top_core_KE_n5479) );
  MX4X1 top_core_KE_U5519 ( .A(top_core_KE_key_mem_8__90_), .B(
        top_core_KE_key_mem_9__90_), .C(top_core_KE_key_mem_10__90_), .D(
        top_core_KE_key_mem_11__90_), .S0(top_core_EC_n864), .S1(n4010), .Y(
        top_core_KE_n5477) );
  MX2X1 top_core_KE_U5518 ( .A(top_core_KE_n5474), .B(top_core_KE_n5475), .S0(
        n4019), .Y(top_core_KE_n5476) );
  MX4X1 top_core_KE_U5522 ( .A(top_core_KE_n5479), .B(top_core_KE_n5477), .C(
        top_core_KE_n5478), .D(top_core_KE_n5476), .S0(n3970), .S1(n3981), .Y(
        top_core_Key[90]) );
  MX4X1 top_core_KE_U5682 ( .A(top_core_KE_key_mem_0__113_), .B(
        top_core_KE_key_mem_1__113_), .C(top_core_KE_key_mem_2__113_), .D(
        top_core_KE_key_mem_3__113_), .S0(n4052), .S1(n4030), .Y(
        top_core_KE_n5617) );
  MX4X1 top_core_KE_U5680 ( .A(top_core_KE_key_mem_8__113_), .B(
        top_core_KE_key_mem_9__113_), .C(top_core_KE_key_mem_10__113_), .D(
        top_core_KE_key_mem_11__113_), .S0(n4052), .S1(n4006), .Y(
        top_core_KE_n5615) );
  MX2X1 top_core_KE_U5679 ( .A(top_core_KE_n5612), .B(top_core_KE_n5613), .S0(
        n4016), .Y(top_core_KE_n5614) );
  MX4X1 top_core_KE_U5683 ( .A(top_core_KE_n5617), .B(top_core_KE_n5615), .C(
        top_core_KE_n5616), .D(top_core_KE_n5614), .S0(n3971), .S1(n3983), .Y(
        top_core_Key[113]) );
  MX4X1 top_core_KE_U5185 ( .A(top_core_KE_key_mem_0__42_), .B(
        top_core_KE_key_mem_1__42_), .C(top_core_KE_key_mem_2__42_), .D(
        top_core_KE_key_mem_3__42_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5191) );
  MX4X1 top_core_KE_U5183 ( .A(top_core_KE_key_mem_8__42_), .B(
        top_core_KE_key_mem_9__42_), .C(top_core_KE_key_mem_10__42_), .D(
        top_core_KE_key_mem_11__42_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5189) );
  MX2X1 top_core_KE_U5182 ( .A(top_core_KE_n5186), .B(top_core_KE_n5187), .S0(
        n4020), .Y(top_core_KE_n5188) );
  MX4X1 top_core_KE_U5186 ( .A(top_core_KE_n5191), .B(top_core_KE_n5189), .C(
        top_core_KE_n5190), .D(top_core_KE_n5188), .S0(n3966), .S1(n3978), .Y(
        top_core_Key[42]) );
  MX4X1 top_core_KE_U5346 ( .A(top_core_KE_key_mem_0__65_), .B(
        top_core_KE_key_mem_1__65_), .C(top_core_KE_key_mem_2__65_), .D(
        top_core_KE_key_mem_3__65_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5329) );
  MX4X1 top_core_KE_U5344 ( .A(top_core_KE_key_mem_8__65_), .B(
        top_core_KE_key_mem_9__65_), .C(top_core_KE_key_mem_10__65_), .D(
        top_core_KE_key_mem_11__65_), .S0(n4041), .S1(n3994), .Y(
        top_core_KE_n5327) );
  MX2X1 top_core_KE_U5343 ( .A(top_core_KE_n5324), .B(top_core_KE_n5325), .S0(
        n4013), .Y(top_core_KE_n5326) );
  MX4X1 top_core_KE_U5347 ( .A(top_core_KE_n5329), .B(top_core_KE_n5327), .C(
        top_core_KE_n5328), .D(top_core_KE_n5326), .S0(n3968), .S1(n3980), .Y(
        top_core_Key[65]) );
  MX4X1 top_core_KE_U5745 ( .A(top_core_KE_key_mem_0__122_), .B(
        top_core_KE_key_mem_1__122_), .C(top_core_KE_key_mem_2__122_), .D(
        top_core_KE_key_mem_3__122_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5671) );
  MX4X1 top_core_KE_U5743 ( .A(top_core_KE_key_mem_8__122_), .B(
        top_core_KE_key_mem_9__122_), .C(top_core_KE_key_mem_10__122_), .D(
        top_core_KE_key_mem_11__122_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5669) );
  MX2X1 top_core_KE_U5742 ( .A(top_core_KE_n5666), .B(top_core_KE_n5667), .S0(
        n4014), .Y(top_core_KE_n5668) );
  MX4X1 top_core_KE_U5746 ( .A(top_core_KE_n5671), .B(top_core_KE_n5669), .C(
        top_core_KE_n5670), .D(top_core_KE_n5668), .S0(n3972), .S1(n3983), .Y(
        top_core_Key[122]) );
  MX4X1 top_core_KE_U5507 ( .A(top_core_KE_key_mem_0__88_), .B(
        top_core_KE_key_mem_1__88_), .C(top_core_KE_key_mem_2__88_), .D(
        top_core_KE_key_mem_3__88_), .S0(n4057), .S1(n4011), .Y(
        top_core_KE_n5467) );
  MX4X1 top_core_KE_U5505 ( .A(top_core_KE_key_mem_8__88_), .B(
        top_core_KE_key_mem_9__88_), .C(top_core_KE_key_mem_10__88_), .D(
        top_core_KE_key_mem_11__88_), .S0(n4057), .S1(n4009), .Y(
        top_core_KE_n5465) );
  MX2X1 top_core_KE_U5504 ( .A(top_core_KE_n5462), .B(top_core_KE_n5463), .S0(
        n4018), .Y(top_core_KE_n5464) );
  MX4X1 top_core_KE_U5508 ( .A(top_core_KE_n5467), .B(top_core_KE_n5465), .C(
        top_core_KE_n5466), .D(top_core_KE_n5464), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[88]) );
  MX4X1 top_core_KE_U5241 ( .A(top_core_KE_key_mem_0__50_), .B(
        top_core_KE_key_mem_1__50_), .C(top_core_KE_key_mem_2__50_), .D(
        top_core_KE_key_mem_3__50_), .S0(n4038), .S1(n3992), .Y(
        top_core_KE_n5239) );
  MX4X1 top_core_KE_U5239 ( .A(top_core_KE_key_mem_8__50_), .B(
        top_core_KE_key_mem_9__50_), .C(top_core_KE_key_mem_10__50_), .D(
        top_core_KE_key_mem_11__50_), .S0(n4038), .S1(n3991), .Y(
        top_core_KE_n5237) );
  MX2X1 top_core_KE_U5238 ( .A(top_core_KE_n5234), .B(top_core_KE_n5235), .S0(
        n4019), .Y(top_core_KE_n5236) );
  MX4X1 top_core_KE_U5242 ( .A(top_core_KE_n5239), .B(top_core_KE_n5237), .C(
        top_core_KE_n5238), .D(top_core_KE_n5236), .S0(n3966), .S1(n3979), .Y(
        top_core_Key[50]) );
  MX4X1 top_core_KE_U5171 ( .A(top_core_KE_key_mem_0__40_), .B(
        top_core_KE_key_mem_1__40_), .C(top_core_KE_key_mem_2__40_), .D(
        top_core_KE_key_mem_3__40_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5179) );
  MX4X1 top_core_KE_U5169 ( .A(top_core_KE_key_mem_8__40_), .B(
        top_core_KE_key_mem_9__40_), .C(top_core_KE_key_mem_10__40_), .D(
        top_core_KE_key_mem_11__40_), .S0(n4035), .S1(n3990), .Y(
        top_core_KE_n5177) );
  MX2X1 top_core_KE_U5168 ( .A(top_core_KE_n5174), .B(top_core_KE_n5175), .S0(
        n4019), .Y(top_core_KE_n5176) );
  MX4X1 top_core_KE_U5172 ( .A(top_core_KE_n5179), .B(top_core_KE_n5177), .C(
        top_core_KE_n5178), .D(top_core_KE_n5176), .S0(n3966), .S1(n3978), .Y(
        top_core_Key[40]) );
  MX4X1 top_core_KE_U5514 ( .A(top_core_KE_key_mem_0__89_), .B(
        top_core_KE_key_mem_1__89_), .C(top_core_KE_key_mem_2__89_), .D(
        top_core_KE_key_mem_3__89_), .S0(top_core_EC_n864), .S1(n4008), .Y(
        top_core_KE_n5473) );
  MX4X1 top_core_KE_U5512 ( .A(top_core_KE_key_mem_8__89_), .B(
        top_core_KE_key_mem_9__89_), .C(top_core_KE_key_mem_10__89_), .D(
        top_core_KE_key_mem_11__89_), .S0(top_core_EC_n864), .S1(n4010), .Y(
        top_core_KE_n5471) );
  MX2X1 top_core_KE_U5511 ( .A(top_core_KE_n5468), .B(top_core_KE_n5469), .S0(
        n4019), .Y(top_core_KE_n5470) );
  MX4X1 top_core_KE_U5515 ( .A(top_core_KE_n5473), .B(top_core_KE_n5471), .C(
        top_core_KE_n5472), .D(top_core_KE_n5470), .S0(n3970), .S1(n3981), .Y(
        top_core_Key[89]) );
  MX4X1 top_core_KE_U5178 ( .A(top_core_KE_key_mem_0__41_), .B(
        top_core_KE_key_mem_1__41_), .C(top_core_KE_key_mem_2__41_), .D(
        top_core_KE_key_mem_3__41_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5185) );
  MX4X1 top_core_KE_U5176 ( .A(top_core_KE_key_mem_8__41_), .B(
        top_core_KE_key_mem_9__41_), .C(top_core_KE_key_mem_10__41_), .D(
        top_core_KE_key_mem_11__41_), .S0(n4036), .S1(n3990), .Y(
        top_core_KE_n5183) );
  MX2X1 top_core_KE_U5175 ( .A(top_core_KE_n5180), .B(top_core_KE_n5181), .S0(
        n4019), .Y(top_core_KE_n5182) );
  MX4X1 top_core_KE_U5179 ( .A(top_core_KE_n5185), .B(top_core_KE_n5183), .C(
        top_core_KE_n5184), .D(top_core_KE_n5182), .S0(n3966), .S1(n3978), .Y(
        top_core_Key[41]) );
  MX4X1 top_core_KE_U5738 ( .A(top_core_KE_key_mem_0__121_), .B(
        top_core_KE_key_mem_1__121_), .C(top_core_KE_key_mem_2__121_), .D(
        top_core_KE_key_mem_3__121_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5665) );
  MX4X1 top_core_KE_U5736 ( .A(top_core_KE_key_mem_8__121_), .B(
        top_core_KE_key_mem_9__121_), .C(top_core_KE_key_mem_10__121_), .D(
        top_core_KE_key_mem_11__121_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5663) );
  MX2X1 top_core_KE_U5735 ( .A(top_core_KE_n5660), .B(top_core_KE_n5661), .S0(
        n4014), .Y(top_core_KE_n5662) );
  MX4X1 top_core_KE_U5739 ( .A(top_core_KE_n5665), .B(top_core_KE_n5663), .C(
        top_core_KE_n5664), .D(top_core_KE_n5662), .S0(n3972), .S1(n3983), .Y(
        top_core_Key[121]) );
  MX4X1 top_core_KE_U5465 ( .A(top_core_KE_key_mem_0__82_), .B(
        top_core_KE_key_mem_1__82_), .C(top_core_KE_key_mem_2__82_), .D(
        top_core_KE_key_mem_3__82_), .S0(n4056), .S1(n4010), .Y(
        top_core_KE_n5431) );
  MX4X1 top_core_KE_U5463 ( .A(top_core_KE_key_mem_8__82_), .B(
        top_core_KE_key_mem_9__82_), .C(top_core_KE_key_mem_10__82_), .D(
        top_core_KE_key_mem_11__82_), .S0(n4056), .S1(n4009), .Y(
        top_core_KE_n5429) );
  MX2X1 top_core_KE_U5462 ( .A(top_core_KE_n5426), .B(top_core_KE_n5427), .S0(
        n4016), .Y(top_core_KE_n5428) );
  MX4X1 top_core_KE_U5466 ( .A(top_core_KE_n5431), .B(top_core_KE_n5429), .C(
        top_core_KE_n5430), .D(top_core_KE_n5428), .S0(n3969), .S1(n3981), .Y(
        top_core_Key[82]) );
  MX4X1 top_core_KE_U5731 ( .A(top_core_KE_key_mem_0__120_), .B(
        top_core_KE_key_mem_1__120_), .C(top_core_KE_key_mem_2__120_), .D(
        top_core_KE_key_mem_3__120_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5659) );
  MX4X1 top_core_KE_U5729 ( .A(top_core_KE_key_mem_8__120_), .B(
        top_core_KE_key_mem_9__120_), .C(top_core_KE_key_mem_10__120_), .D(
        top_core_KE_key_mem_11__120_), .S0(n4054), .S1(n4007), .Y(
        top_core_KE_n5657) );
  MX2X1 top_core_KE_U5728 ( .A(top_core_KE_n5654), .B(top_core_KE_n5655), .S0(
        n4014), .Y(top_core_KE_n5656) );
  MX4X1 top_core_KE_U5732 ( .A(top_core_KE_n5659), .B(top_core_KE_n5657), .C(
        top_core_KE_n5658), .D(top_core_KE_n5656), .S0(n3972), .S1(n3983), .Y(
        top_core_Key[120]) );
  MX4X1 top_core_KE_U5785 ( .A(top_core_KE_key_mem_8__128_), .B(
        top_core_KE_key_mem_9__128_), .C(top_core_KE_key_mem_10__128_), .D(
        top_core_KE_key_mem_11__128_), .S0(n4045), .S1(n4008), .Y(
        top_core_KE_n5705) );
  MX2X1 top_core_KE_U5784 ( .A(top_core_KE_n5702), .B(top_core_KE_n5703), .S0(
        n4015), .Y(top_core_KE_n5704) );
  MX4X1 top_core_KE_U5788 ( .A(top_core_KE_n5707), .B(top_core_KE_n5705), .C(
        top_core_KE_n5706), .D(top_core_KE_n5704), .S0(n3963), .S1(n3976), .Y(
        top_core_Key[128]) );
  MX4X1 top_core_io_U1593 ( .A(top_core_io_n1192), .B(top_core_io_n1190), .C(
        top_core_io_n1191), .D(top_core_io_n1189), .S0(n4141), .S1(n_ADDR[2]), 
        .Y(top_core_io_n1193) );
  MX4X1 top_core_io_U1738 ( .A(top_core_io_CipherKey_w_39_), .B(
        top_core_io_CipherKey_w_47_), .C(top_core_io_CipherKey_w_55_), .D(
        top_core_io_CipherKey_w_63_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1331) );
  MX4X1 top_core_io_U1737 ( .A(top_core_io_CipherKey_w_71_), .B(
        top_core_io_CipherKey_w_79_), .C(top_core_io_CipherKey_w_87_), .D(
        top_core_io_CipherKey_w_95_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1330) );
  MX4X1 top_core_io_U1739 ( .A(top_core_io_CipherKey_w_7_), .B(
        top_core_io_CipherKey_w_15_), .C(top_core_io_CipherKey_w_23_), .D(
        top_core_io_CipherKey_w_31_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1332) );
  MX4X1 top_core_io_U1612 ( .A(top_core_io_CipherKey_w_33_), .B(
        top_core_io_CipherKey_w_41_), .C(top_core_io_CipherKey_w_49_), .D(
        top_core_io_CipherKey_w_57_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1211) );
  MX4X1 top_core_io_U1611 ( .A(top_core_io_CipherKey_w_65_), .B(
        top_core_io_CipherKey_w_73_), .C(top_core_io_CipherKey_w_81_), .D(
        top_core_io_CipherKey_w_89_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1210) );
  MX4X1 top_core_io_U1613 ( .A(top_core_io_CipherKey_w_1_), .B(
        top_core_io_CipherKey_w_9_), .C(top_core_io_CipherKey_w_17_), .D(
        top_core_io_CipherKey_w_25_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1212) );
  MX4X1 top_core_io_U1614 ( .A(top_core_io_n1212), .B(top_core_io_n1210), .C(
        top_core_io_n1211), .D(top_core_io_n1209), .S0(n4141), .S1(n_ADDR[2]), 
        .Y(top_core_io_n1213) );
  MX4X1 top_core_io_U1633 ( .A(top_core_io_CipherKey_w_34_), .B(
        top_core_io_CipherKey_w_42_), .C(top_core_io_CipherKey_w_50_), .D(
        top_core_io_CipherKey_w_58_), .S0(n4119), .S1(n4130), .Y(
        top_core_io_n1231) );
  MX4X1 top_core_io_U1632 ( .A(top_core_io_CipherKey_w_66_), .B(
        top_core_io_CipherKey_w_74_), .C(top_core_io_CipherKey_w_82_), .D(
        top_core_io_CipherKey_w_90_), .S0(n4119), .S1(n4130), .Y(
        top_core_io_n1230) );
  MX4X1 top_core_io_U1634 ( .A(top_core_io_CipherKey_w_2_), .B(
        top_core_io_CipherKey_w_10_), .C(top_core_io_CipherKey_w_18_), .D(
        top_core_io_CipherKey_w_26_), .S0(n4119), .S1(n4130), .Y(
        top_core_io_n1232) );
  MX4X1 top_core_io_U1635 ( .A(top_core_io_n1232), .B(top_core_io_n1230), .C(
        top_core_io_n1231), .D(top_core_io_n1229), .S0(n4141), .S1(n4139), .Y(
        top_core_io_n1233) );
  MX4X1 top_core_io_U1588 ( .A(top_core_io_n1187), .B(top_core_io_n1185), .C(
        top_core_io_n1186), .D(top_core_io_n1184), .S0(n4141), .S1(n_ADDR[2]), 
        .Y(top_core_io_n1188) );
  MX4X1 top_core_io_U1649 ( .A(top_core_io_CipherKey_w_163_), .B(
        top_core_io_CipherKey_w_171_), .C(top_core_io_CipherKey_w_179_), .D(
        top_core_io_CipherKey_w_187_), .S0(n4116), .S1(n4131), .Y(
        top_core_io_n1246) );
  MX4X1 top_core_io_U1648 ( .A(top_core_io_CipherKey_w_195_), .B(
        top_core_io_CipherKey_w_203_), .C(top_core_io_CipherKey_w_211_), .D(
        top_core_io_CipherKey_w_219_), .S0(n4120), .S1(n4131), .Y(
        top_core_io_n1245) );
  MX4X1 top_core_io_U1650 ( .A(top_core_io_CipherKey_w_131_), .B(
        top_core_io_CipherKey_w_139_), .C(top_core_io_CipherKey_w_147_), .D(
        top_core_io_CipherKey_w_155_), .S0(n4123), .S1(n4131), .Y(
        top_core_io_n1247) );
  MX4X1 top_core_io_U1651 ( .A(top_core_io_n1247), .B(top_core_io_n1245), .C(
        top_core_io_n1246), .D(top_core_io_n1244), .S0(n_ADDR[3]), .S1(n4139), 
        .Y(top_core_io_n1248) );
  MX4X1 top_core_io_U1670 ( .A(top_core_io_CipherKey_w_164_), .B(
        top_core_io_CipherKey_w_172_), .C(top_core_io_CipherKey_w_180_), .D(
        top_core_io_CipherKey_w_188_), .S0(n4120), .S1(n4131), .Y(
        top_core_io_n1266) );
  MX4X1 top_core_io_U1669 ( .A(top_core_io_CipherKey_w_196_), .B(
        top_core_io_CipherKey_w_204_), .C(top_core_io_CipherKey_w_212_), .D(
        top_core_io_CipherKey_w_220_), .S0(n4120), .S1(n_ADDR[1]), .Y(
        top_core_io_n1265) );
  MX4X1 top_core_io_U1671 ( .A(top_core_io_CipherKey_w_132_), .B(
        top_core_io_CipherKey_w_140_), .C(top_core_io_CipherKey_w_148_), .D(
        top_core_io_CipherKey_w_156_), .S0(n4120), .S1(n4132), .Y(
        top_core_io_n1267) );
  MX4X1 top_core_io_U1672 ( .A(top_core_io_n1267), .B(top_core_io_n1265), .C(
        top_core_io_n1266), .D(top_core_io_n1264), .S0(n4141), .S1(n4139), .Y(
        top_core_io_n1268) );
  MX4X1 top_core_io_U1691 ( .A(top_core_io_CipherKey_w_165_), .B(
        top_core_io_CipherKey_w_173_), .C(top_core_io_CipherKey_w_181_), .D(
        top_core_io_CipherKey_w_189_), .S0(n4121), .S1(n4133), .Y(
        top_core_io_n1286) );
  MX4X1 top_core_io_U1690 ( .A(top_core_io_CipherKey_w_197_), .B(
        top_core_io_CipherKey_w_205_), .C(top_core_io_CipherKey_w_213_), .D(
        top_core_io_CipherKey_w_221_), .S0(n4121), .S1(n4133), .Y(
        top_core_io_n1285) );
  MX4X1 top_core_io_U1692 ( .A(top_core_io_CipherKey_w_133_), .B(
        top_core_io_CipherKey_w_141_), .C(top_core_io_CipherKey_w_149_), .D(
        top_core_io_CipherKey_w_157_), .S0(n4121), .S1(n4133), .Y(
        top_core_io_n1287) );
  MX4X1 top_core_io_U1693 ( .A(top_core_io_n1287), .B(top_core_io_n1285), .C(
        top_core_io_n1286), .D(top_core_io_n1284), .S0(n4141), .S1(n4139), .Y(
        top_core_io_n1288) );
  MX4X1 top_core_io_U1712 ( .A(top_core_io_CipherKey_w_166_), .B(
        top_core_io_CipherKey_w_174_), .C(top_core_io_CipherKey_w_182_), .D(
        top_core_io_CipherKey_w_190_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1306) );
  MX4X1 top_core_io_U1711 ( .A(top_core_io_CipherKey_w_198_), .B(
        top_core_io_CipherKey_w_206_), .C(top_core_io_CipherKey_w_214_), .D(
        top_core_io_CipherKey_w_222_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1305) );
  MX4X1 top_core_io_U1713 ( .A(top_core_io_CipherKey_w_134_), .B(
        top_core_io_CipherKey_w_142_), .C(top_core_io_CipherKey_w_150_), .D(
        top_core_io_CipherKey_w_158_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1307) );
  MX4X1 top_core_io_U1733 ( .A(top_core_io_CipherKey_w_167_), .B(
        top_core_io_CipherKey_w_175_), .C(top_core_io_CipherKey_w_183_), .D(
        top_core_io_CipherKey_w_191_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1326) );
  MX4X1 top_core_io_U1732 ( .A(top_core_io_CipherKey_w_199_), .B(
        top_core_io_CipherKey_w_207_), .C(top_core_io_CipherKey_w_215_), .D(
        top_core_io_CipherKey_w_223_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1325) );
  MX4X1 top_core_io_U1734 ( .A(top_core_io_CipherKey_w_135_), .B(
        top_core_io_CipherKey_w_143_), .C(top_core_io_CipherKey_w_151_), .D(
        top_core_io_CipherKey_w_159_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1327) );
  MX4X1 top_core_io_U1742 ( .A(top_core_io_Data_reg_24__7_), .B(
        top_core_io_Data_reg_25__7_), .C(top_core_io_Data_reg_26__7_), .D(
        top_core_io_Data_reg_27__7_), .S0(n4124), .S1(n4135), .Y(
        top_core_io_n1335) );
  MX4X1 top_core_io_U1598 ( .A(top_core_io_n1197), .B(top_core_io_n1195), .C(
        top_core_io_n1196), .D(top_core_io_n1194), .S0(n4141), .S1(n_ADDR[2]), 
        .Y(top_core_io_n1198) );
  MX4X1 top_core_io_U1659 ( .A(top_core_io_Data_reg_20__3_), .B(
        top_core_io_Data_reg_21__3_), .C(top_core_io_Data_reg_22__3_), .D(
        top_core_io_Data_reg_23__3_), .S0(n4117), .S1(n4134), .Y(
        top_core_io_n1256) );
  MX4X1 top_core_io_U1658 ( .A(top_core_io_Data_reg_24__3_), .B(
        top_core_io_Data_reg_25__3_), .C(top_core_io_Data_reg_26__3_), .D(
        top_core_io_Data_reg_27__3_), .S0(n4122), .S1(n_ADDR[1]), .Y(
        top_core_io_n1255) );
  MX4X1 top_core_io_U1660 ( .A(top_core_io_Data_reg_16__3_), .B(
        top_core_io_Data_reg_17__3_), .C(top_core_io_Data_reg_18__3_), .D(
        top_core_io_Data_reg_19__3_), .S0(n4123), .S1(n4131), .Y(
        top_core_io_n1257) );
  MX4X1 top_core_io_U1661 ( .A(top_core_io_n1257), .B(top_core_io_n1255), .C(
        top_core_io_n1256), .D(top_core_io_n1254), .S0(n_ADDR[3]), .S1(n4139), 
        .Y(top_core_io_n1258) );
  MX4X1 top_core_io_U1680 ( .A(top_core_io_Data_reg_20__4_), .B(
        top_core_io_Data_reg_21__4_), .C(top_core_io_Data_reg_22__4_), .D(
        top_core_io_Data_reg_23__4_), .S0(n4121), .S1(n4132), .Y(
        top_core_io_n1276) );
  MX4X1 top_core_io_U1679 ( .A(top_core_io_Data_reg_24__4_), .B(
        top_core_io_Data_reg_25__4_), .C(top_core_io_Data_reg_26__4_), .D(
        top_core_io_Data_reg_27__4_), .S0(n4121), .S1(n4132), .Y(
        top_core_io_n1275) );
  MX4X1 top_core_io_U1681 ( .A(top_core_io_Data_reg_16__4_), .B(
        top_core_io_Data_reg_17__4_), .C(top_core_io_Data_reg_18__4_), .D(
        top_core_io_Data_reg_19__4_), .S0(n4121), .S1(n4132), .Y(
        top_core_io_n1277) );
  MX4X1 top_core_io_U1682 ( .A(top_core_io_n1277), .B(top_core_io_n1275), .C(
        top_core_io_n1276), .D(top_core_io_n1274), .S0(n_ADDR[3]), .S1(n4139), 
        .Y(top_core_io_n1278) );
  MX4X1 top_core_io_U1701 ( .A(top_core_io_Data_reg_20__5_), .B(
        top_core_io_Data_reg_21__5_), .C(top_core_io_Data_reg_22__5_), .D(
        top_core_io_Data_reg_23__5_), .S0(n4118), .S1(n4133), .Y(
        top_core_io_n1296) );
  MX4X1 top_core_io_U1700 ( .A(top_core_io_Data_reg_24__5_), .B(
        top_core_io_Data_reg_25__5_), .C(top_core_io_Data_reg_26__5_), .D(
        top_core_io_Data_reg_27__5_), .S0(n_ADDR[0]), .S1(n4133), .Y(
        top_core_io_n1295) );
  MX4X1 top_core_io_U1702 ( .A(top_core_io_Data_reg_16__5_), .B(
        top_core_io_Data_reg_17__5_), .C(top_core_io_Data_reg_18__5_), .D(
        top_core_io_Data_reg_19__5_), .S0(n_ADDR[0]), .S1(n4133), .Y(
        top_core_io_n1297) );
  MX4X1 top_core_io_U1703 ( .A(top_core_io_n1297), .B(top_core_io_n1295), .C(
        top_core_io_n1296), .D(top_core_io_n1294), .S0(n_ADDR[3]), .S1(n4138), 
        .Y(top_core_io_n1298) );
  MX4X1 top_core_io_U1722 ( .A(top_core_io_Data_reg_20__6_), .B(
        top_core_io_Data_reg_21__6_), .C(top_core_io_Data_reg_22__6_), .D(
        top_core_io_Data_reg_23__6_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1316) );
  MX4X1 top_core_io_U1721 ( .A(top_core_io_Data_reg_24__6_), .B(
        top_core_io_Data_reg_25__6_), .C(top_core_io_Data_reg_26__6_), .D(
        top_core_io_Data_reg_27__6_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1315) );
  MX4X1 top_core_io_U1723 ( .A(top_core_io_Data_reg_16__6_), .B(
        top_core_io_Data_reg_17__6_), .C(top_core_io_Data_reg_18__6_), .D(
        top_core_io_Data_reg_19__6_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1317) );
  MX4X1 top_core_io_U1657 ( .A(top_core_io_Data_reg_28__3_), .B(
        top_core_io_Data_reg_29__3_), .C(top_core_io_Data_reg_30__3_), .D(
        top_core_io_Data_reg_31__3_), .S0(n4121), .S1(n4130), .Y(
        top_core_io_n1254) );
  MX4X1 top_core_io_U1678 ( .A(top_core_io_Data_reg_28__4_), .B(
        top_core_io_Data_reg_29__4_), .C(top_core_io_Data_reg_30__4_), .D(
        top_core_io_Data_reg_31__4_), .S0(n4121), .S1(n4132), .Y(
        top_core_io_n1274) );
  MX4X1 top_core_io_U1699 ( .A(top_core_io_Data_reg_28__5_), .B(
        top_core_io_Data_reg_29__5_), .C(top_core_io_Data_reg_30__5_), .D(
        top_core_io_Data_reg_31__5_), .S0(n4119), .S1(n4133), .Y(
        top_core_io_n1294) );
  MX4X1 top_core_io_U1720 ( .A(top_core_io_Data_reg_28__6_), .B(
        top_core_io_Data_reg_29__6_), .C(top_core_io_Data_reg_30__6_), .D(
        top_core_io_Data_reg_31__6_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1314) );
  MX4X1 top_core_io_U1741 ( .A(top_core_io_Data_reg_28__7_), .B(
        top_core_io_Data_reg_29__7_), .C(top_core_io_Data_reg_30__7_), .D(
        top_core_io_Data_reg_31__7_), .S0(n4124), .S1(n4135), .Y(
        top_core_io_n1334) );
  MX4X1 top_core_io_U1600 ( .A(top_core_io_Plain_text_w_64_), .B(
        top_core_io_Plain_text_w_72_), .C(top_core_io_Plain_text_w_80_), .D(
        top_core_io_Plain_text_w_88_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1200) );
  MX4X1 top_core_io_U1663 ( .A(top_core_io_Plain_text_w_67_), .B(
        top_core_io_Plain_text_w_75_), .C(top_core_io_Plain_text_w_83_), .D(
        top_core_io_Plain_text_w_91_), .S0(n4120), .S1(n_ADDR[1]), .Y(
        top_core_io_n1260) );
  MX4X1 top_core_io_U1653 ( .A(top_core_io_CipherKey_w_67_), .B(
        top_core_io_CipherKey_w_75_), .C(top_core_io_CipherKey_w_83_), .D(
        top_core_io_CipherKey_w_91_), .S0(n4116), .S1(n4131), .Y(
        top_core_io_n1250) );
  MX4X1 top_core_io_U1684 ( .A(top_core_io_Plain_text_w_68_), .B(
        top_core_io_Plain_text_w_76_), .C(top_core_io_Plain_text_w_84_), .D(
        top_core_io_Plain_text_w_92_), .S0(n4121), .S1(n4132), .Y(
        top_core_io_n1280) );
  MX4X1 top_core_io_U1674 ( .A(top_core_io_CipherKey_w_68_), .B(
        top_core_io_CipherKey_w_76_), .C(top_core_io_CipherKey_w_84_), .D(
        top_core_io_CipherKey_w_92_), .S0(n4120), .S1(n4132), .Y(
        top_core_io_n1270) );
  MX4X1 top_core_io_U1705 ( .A(top_core_io_Plain_text_w_69_), .B(
        top_core_io_Plain_text_w_77_), .C(top_core_io_Plain_text_w_85_), .D(
        top_core_io_Plain_text_w_93_), .S0(n_ADDR[0]), .S1(n4133), .Y(
        top_core_io_n1300) );
  MX4X1 top_core_io_U1695 ( .A(top_core_io_CipherKey_w_69_), .B(
        top_core_io_CipherKey_w_77_), .C(top_core_io_CipherKey_w_85_), .D(
        top_core_io_CipherKey_w_93_), .S0(n_ADDR[0]), .S1(n4133), .Y(
        top_core_io_n1290) );
  MX4X1 top_core_io_U1726 ( .A(top_core_io_Plain_text_w_70_), .B(
        top_core_io_Plain_text_w_78_), .C(top_core_io_Plain_text_w_86_), .D(
        top_core_io_Plain_text_w_94_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1320) );
  MX4X1 top_core_io_U1716 ( .A(top_core_io_CipherKey_w_70_), .B(
        top_core_io_CipherKey_w_78_), .C(top_core_io_CipherKey_w_86_), .D(
        top_core_io_CipherKey_w_94_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1310) );
  MX4X1 top_core_io_U1747 ( .A(top_core_io_Plain_text_w_71_), .B(
        top_core_io_Plain_text_w_79_), .C(top_core_io_Plain_text_w_87_), .D(
        top_core_io_Plain_text_w_95_), .S0(n4124), .S1(n4133), .Y(
        top_core_io_n1340) );
  MX4X1 top_core_io_U1621 ( .A(top_core_io_Plain_text_w_65_), .B(
        top_core_io_Plain_text_w_73_), .C(top_core_io_Plain_text_w_81_), .D(
        top_core_io_Plain_text_w_89_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1220) );
  MX4X1 top_core_io_U1642 ( .A(top_core_io_Plain_text_w_66_), .B(
        top_core_io_Plain_text_w_74_), .C(top_core_io_Plain_text_w_82_), .D(
        top_core_io_Plain_text_w_90_), .S0(n4119), .S1(n4131), .Y(
        top_core_io_n1240) );
  MX4X1 top_core_io_U1744 ( .A(top_core_io_Data_reg_16__7_), .B(
        top_core_io_Data_reg_17__7_), .C(top_core_io_Data_reg_18__7_), .D(
        top_core_io_Data_reg_19__7_), .S0(n4124), .S1(n4132), .Y(
        top_core_io_n1337) );
  MX4X1 top_core_io_U1599 ( .A(top_core_io_Plain_text_w_96_), .B(
        top_core_io_Plain_text_w_104_), .C(top_core_io_Plain_text_w_112_), .D(
        top_core_io_Plain_text_w_120_), .S0(n4116), .S1(n4129), .Y(
        top_core_io_n1199) );
  MX4X1 top_core_io_U1584 ( .A(top_core_io_CipherKey_w_224_), .B(
        top_core_io_CipherKey_w_232_), .C(top_core_io_CipherKey_w_240_), .D(
        top_core_io_CipherKey_w_248_), .S0(n4120), .S1(n4134), .Y(
        top_core_io_n1184) );
  MX4X1 top_core_io_U1662 ( .A(top_core_io_Plain_text_w_99_), .B(
        top_core_io_Plain_text_w_107_), .C(top_core_io_Plain_text_w_115_), .D(
        top_core_io_Plain_text_w_123_), .S0(n4122), .S1(n4129), .Y(
        top_core_io_n1259) );
  MX4X1 top_core_io_U1652 ( .A(top_core_io_CipherKey_w_99_), .B(
        top_core_io_CipherKey_w_107_), .C(top_core_io_CipherKey_w_115_), .D(
        top_core_io_CipherKey_w_123_), .S0(n4121), .S1(n4131), .Y(
        top_core_io_n1249) );
  MX4X1 top_core_io_U1647 ( .A(top_core_io_CipherKey_w_227_), .B(
        top_core_io_CipherKey_w_235_), .C(top_core_io_CipherKey_w_243_), .D(
        top_core_io_CipherKey_w_251_), .S0(n4119), .S1(n4131), .Y(
        top_core_io_n1244) );
  MX4X1 top_core_io_U1683 ( .A(top_core_io_Plain_text_w_100_), .B(
        top_core_io_Plain_text_w_108_), .C(top_core_io_Plain_text_w_116_), .D(
        top_core_io_Plain_text_w_124_), .S0(n4121), .S1(n4132), .Y(
        top_core_io_n1279) );
  MX4X1 top_core_io_U1673 ( .A(top_core_io_CipherKey_w_100_), .B(
        top_core_io_CipherKey_w_108_), .C(top_core_io_CipherKey_w_116_), .D(
        top_core_io_CipherKey_w_124_), .S0(n4120), .S1(n4132), .Y(
        top_core_io_n1269) );
  MX4X1 top_core_io_U1668 ( .A(top_core_io_CipherKey_w_228_), .B(
        top_core_io_CipherKey_w_236_), .C(top_core_io_CipherKey_w_244_), .D(
        top_core_io_CipherKey_w_252_), .S0(n4120), .S1(n4129), .Y(
        top_core_io_n1264) );
  MX4X1 top_core_io_U1704 ( .A(top_core_io_Plain_text_w_101_), .B(
        top_core_io_Plain_text_w_109_), .C(top_core_io_Plain_text_w_117_), .D(
        top_core_io_Plain_text_w_125_), .S0(n4117), .S1(n4133), .Y(
        top_core_io_n1299) );
  MX4X1 top_core_io_U1694 ( .A(top_core_io_CipherKey_w_101_), .B(
        top_core_io_CipherKey_w_109_), .C(top_core_io_CipherKey_w_117_), .D(
        top_core_io_CipherKey_w_125_), .S0(n4119), .S1(n4133), .Y(
        top_core_io_n1289) );
  MX4X1 top_core_io_U1689 ( .A(top_core_io_CipherKey_w_229_), .B(
        top_core_io_CipherKey_w_237_), .C(top_core_io_CipherKey_w_245_), .D(
        top_core_io_CipherKey_w_253_), .S0(n4121), .S1(n4132), .Y(
        top_core_io_n1284) );
  MX4X1 top_core_io_U1725 ( .A(top_core_io_Plain_text_w_102_), .B(
        top_core_io_Plain_text_w_110_), .C(top_core_io_Plain_text_w_118_), .D(
        top_core_io_Plain_text_w_126_), .S0(n4123), .S1(n4134), .Y(
        top_core_io_n1319) );
  MX4X1 top_core_io_U1715 ( .A(top_core_io_CipherKey_w_102_), .B(
        top_core_io_CipherKey_w_110_), .C(top_core_io_CipherKey_w_118_), .D(
        top_core_io_CipherKey_w_126_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1309) );
  MX4X1 top_core_io_U1710 ( .A(top_core_io_CipherKey_w_230_), .B(
        top_core_io_CipherKey_w_238_), .C(top_core_io_CipherKey_w_246_), .D(
        top_core_io_CipherKey_w_254_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1304) );
  MX4X1 top_core_io_U1746 ( .A(top_core_io_Plain_text_w_103_), .B(
        top_core_io_Plain_text_w_111_), .C(top_core_io_Plain_text_w_119_), .D(
        top_core_io_Plain_text_w_127_), .S0(n4124), .S1(n4135), .Y(
        top_core_io_n1339) );
  MX4X1 top_core_io_U1736 ( .A(top_core_io_CipherKey_w_103_), .B(
        top_core_io_CipherKey_w_111_), .C(top_core_io_CipherKey_w_119_), .D(
        top_core_io_CipherKey_w_127_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1329) );
  MX4X1 top_core_io_U1731 ( .A(top_core_io_CipherKey_w_231_), .B(
        top_core_io_CipherKey_w_239_), .C(top_core_io_CipherKey_w_247_), .D(
        top_core_io_CipherKey_w_255_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1324) );
  MX4X1 top_core_io_U1620 ( .A(top_core_io_Plain_text_w_97_), .B(
        top_core_io_Plain_text_w_105_), .C(top_core_io_Plain_text_w_113_), .D(
        top_core_io_Plain_text_w_121_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1219) );
  MX4X1 top_core_io_U1610 ( .A(top_core_io_CipherKey_w_97_), .B(
        top_core_io_CipherKey_w_105_), .C(top_core_io_CipherKey_w_113_), .D(
        top_core_io_CipherKey_w_121_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1209) );
  MX4X1 top_core_io_U1641 ( .A(top_core_io_Plain_text_w_98_), .B(
        top_core_io_Plain_text_w_106_), .C(top_core_io_Plain_text_w_114_), .D(
        top_core_io_Plain_text_w_122_), .S0(n4119), .S1(n4131), .Y(
        top_core_io_n1239) );
  MX4X1 top_core_io_U1631 ( .A(top_core_io_CipherKey_w_98_), .B(
        top_core_io_CipherKey_w_106_), .C(top_core_io_CipherKey_w_114_), .D(
        top_core_io_CipherKey_w_122_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1229) );
  MX4X1 top_core_io_U1743 ( .A(top_core_io_Data_reg_20__7_), .B(
        top_core_io_Data_reg_21__7_), .C(top_core_io_Data_reg_22__7_), .D(
        top_core_io_Data_reg_23__7_), .S0(n4124), .S1(n4135), .Y(
        top_core_io_n1336) );
  MX4X1 top_core_io_U1602 ( .A(top_core_io_Plain_text_w_0_), .B(
        top_core_io_Plain_text_w_8_), .C(top_core_io_Plain_text_w_16_), .D(
        top_core_io_Plain_text_w_24_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1202) );
  MX4X1 top_core_io_U1665 ( .A(top_core_io_Plain_text_w_3_), .B(
        top_core_io_Plain_text_w_11_), .C(top_core_io_Plain_text_w_19_), .D(
        top_core_io_Plain_text_w_27_), .S0(n4120), .S1(n_ADDR[1]), .Y(
        top_core_io_n1262) );
  MX4X1 top_core_io_U1655 ( .A(top_core_io_CipherKey_w_3_), .B(
        top_core_io_CipherKey_w_11_), .C(top_core_io_CipherKey_w_19_), .D(
        top_core_io_CipherKey_w_27_), .S0(n4116), .S1(n_ADDR[1]), .Y(
        top_core_io_n1252) );
  MX4X1 top_core_io_U1686 ( .A(top_core_io_Plain_text_w_4_), .B(
        top_core_io_Plain_text_w_12_), .C(top_core_io_Plain_text_w_20_), .D(
        top_core_io_Plain_text_w_28_), .S0(n4121), .S1(n4132), .Y(
        top_core_io_n1282) );
  MX4X1 top_core_io_U1676 ( .A(top_core_io_CipherKey_w_4_), .B(
        top_core_io_CipherKey_w_12_), .C(top_core_io_CipherKey_w_20_), .D(
        top_core_io_CipherKey_w_28_), .S0(n4120), .S1(n4132), .Y(
        top_core_io_n1272) );
  MX4X1 top_core_io_U1707 ( .A(top_core_io_Plain_text_w_5_), .B(
        top_core_io_Plain_text_w_13_), .C(top_core_io_Plain_text_w_21_), .D(
        top_core_io_Plain_text_w_29_), .S0(n_ADDR[0]), .S1(n4134), .Y(
        top_core_io_n1302) );
  MX4X1 top_core_io_U1697 ( .A(top_core_io_CipherKey_w_5_), .B(
        top_core_io_CipherKey_w_13_), .C(top_core_io_CipherKey_w_21_), .D(
        top_core_io_CipherKey_w_29_), .S0(n_ADDR[0]), .S1(n4133), .Y(
        top_core_io_n1292) );
  MX4X1 top_core_io_U1728 ( .A(top_core_io_Plain_text_w_6_), .B(
        top_core_io_Plain_text_w_14_), .C(top_core_io_Plain_text_w_22_), .D(
        top_core_io_Plain_text_w_30_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1322) );
  MX4X1 top_core_io_U1718 ( .A(top_core_io_CipherKey_w_6_), .B(
        top_core_io_CipherKey_w_14_), .C(top_core_io_CipherKey_w_22_), .D(
        top_core_io_CipherKey_w_30_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1312) );
  MX4X1 top_core_io_U1749 ( .A(top_core_io_Plain_text_w_7_), .B(
        top_core_io_Plain_text_w_15_), .C(top_core_io_Plain_text_w_23_), .D(
        top_core_io_Plain_text_w_31_), .S0(n4124), .S1(n4133), .Y(
        top_core_io_n1342) );
  MX4X1 top_core_io_U1623 ( .A(top_core_io_Plain_text_w_1_), .B(
        top_core_io_Plain_text_w_9_), .C(top_core_io_Plain_text_w_17_), .D(
        top_core_io_Plain_text_w_25_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1222) );
  MX4X1 top_core_io_U1644 ( .A(top_core_io_Plain_text_w_2_), .B(
        top_core_io_Plain_text_w_10_), .C(top_core_io_Plain_text_w_18_), .D(
        top_core_io_Plain_text_w_26_), .S0(n4119), .S1(n4131), .Y(
        top_core_io_n1242) );
  MX4X1 top_core_io_U1601 ( .A(top_core_io_Plain_text_w_32_), .B(
        top_core_io_Plain_text_w_40_), .C(top_core_io_Plain_text_w_48_), .D(
        top_core_io_Plain_text_w_56_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1201) );
  MX4X1 top_core_io_U1664 ( .A(top_core_io_Plain_text_w_35_), .B(
        top_core_io_Plain_text_w_43_), .C(top_core_io_Plain_text_w_51_), .D(
        top_core_io_Plain_text_w_59_), .S0(n4120), .S1(n4130), .Y(
        top_core_io_n1261) );
  MX4X1 top_core_io_U1654 ( .A(top_core_io_CipherKey_w_35_), .B(
        top_core_io_CipherKey_w_43_), .C(top_core_io_CipherKey_w_51_), .D(
        top_core_io_CipherKey_w_59_), .S0(n4120), .S1(n_ADDR[1]), .Y(
        top_core_io_n1251) );
  MX4X1 top_core_io_U1685 ( .A(top_core_io_Plain_text_w_36_), .B(
        top_core_io_Plain_text_w_44_), .C(top_core_io_Plain_text_w_52_), .D(
        top_core_io_Plain_text_w_60_), .S0(n4121), .S1(n4132), .Y(
        top_core_io_n1281) );
  MX4X1 top_core_io_U1675 ( .A(top_core_io_CipherKey_w_36_), .B(
        top_core_io_CipherKey_w_44_), .C(top_core_io_CipherKey_w_52_), .D(
        top_core_io_CipherKey_w_60_), .S0(n4120), .S1(n4132), .Y(
        top_core_io_n1271) );
  MX4X1 top_core_io_U1706 ( .A(top_core_io_Plain_text_w_37_), .B(
        top_core_io_Plain_text_w_45_), .C(top_core_io_Plain_text_w_53_), .D(
        top_core_io_Plain_text_w_61_), .S0(n_ADDR[0]), .S1(n4133), .Y(
        top_core_io_n1301) );
  MX4X1 top_core_io_U1696 ( .A(top_core_io_CipherKey_w_37_), .B(
        top_core_io_CipherKey_w_45_), .C(top_core_io_CipherKey_w_53_), .D(
        top_core_io_CipherKey_w_61_), .S0(n4118), .S1(n4133), .Y(
        top_core_io_n1291) );
  MX4X1 top_core_io_U1727 ( .A(top_core_io_Plain_text_w_38_), .B(
        top_core_io_Plain_text_w_46_), .C(top_core_io_Plain_text_w_54_), .D(
        top_core_io_Plain_text_w_62_), .S0(n4123), .S1(n4135), .Y(
        top_core_io_n1321) );
  MX4X1 top_core_io_U1717 ( .A(top_core_io_CipherKey_w_38_), .B(
        top_core_io_CipherKey_w_46_), .C(top_core_io_CipherKey_w_54_), .D(
        top_core_io_CipherKey_w_62_), .S0(n4122), .S1(n4134), .Y(
        top_core_io_n1311) );
  MX4X1 top_core_io_U1748 ( .A(top_core_io_Plain_text_w_39_), .B(
        top_core_io_Plain_text_w_47_), .C(top_core_io_Plain_text_w_55_), .D(
        top_core_io_Plain_text_w_63_), .S0(n4124), .S1(n4135), .Y(
        top_core_io_n1341) );
  MX4X1 top_core_io_U1622 ( .A(top_core_io_Plain_text_w_33_), .B(
        top_core_io_Plain_text_w_41_), .C(top_core_io_Plain_text_w_49_), .D(
        top_core_io_Plain_text_w_57_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1221) );
  MX4X1 top_core_io_U1643 ( .A(top_core_io_Plain_text_w_34_), .B(
        top_core_io_Plain_text_w_42_), .C(top_core_io_Plain_text_w_50_), .D(
        top_core_io_Plain_text_w_58_), .S0(n4119), .S1(n4131), .Y(
        top_core_io_n1241) );
  MX4X1 top_core_io_U1603 ( .A(top_core_io_n1202), .B(top_core_io_n1200), .C(
        top_core_io_n1201), .D(top_core_io_n1199), .S0(n4141), .S1(n_ADDR[2]), 
        .Y(top_core_io_n1203) );
  MX4X1 top_core_io_U1604 ( .A(top_core_io_n1203), .B(top_core_io_n1193), .C(
        top_core_io_n1198), .D(top_core_io_n1188), .S0(n_ADDR[5]), .S1(
        n_ADDR[4]), .Y(top_core_io_N81) );
  MX4X1 top_core_io_U1607 ( .A(top_core_io_CipherKey_w_161_), .B(
        top_core_io_CipherKey_w_169_), .C(top_core_io_CipherKey_w_177_), .D(
        top_core_io_CipherKey_w_185_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1206) );
  MX4X1 top_core_io_U1606 ( .A(top_core_io_CipherKey_w_193_), .B(
        top_core_io_CipherKey_w_201_), .C(top_core_io_CipherKey_w_209_), .D(
        top_core_io_CipherKey_w_217_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1205) );
  MX4X1 top_core_io_U1608 ( .A(top_core_io_CipherKey_w_129_), .B(
        top_core_io_CipherKey_w_137_), .C(top_core_io_CipherKey_w_145_), .D(
        top_core_io_CipherKey_w_153_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1207) );
  MX4X1 top_core_io_U1609 ( .A(top_core_io_n1207), .B(top_core_io_n1205), .C(
        top_core_io_n1206), .D(top_core_io_n1204), .S0(n4141), .S1(n4139), .Y(
        top_core_io_n1208) );
  MX4X1 top_core_io_U1628 ( .A(top_core_io_CipherKey_w_162_), .B(
        top_core_io_CipherKey_w_170_), .C(top_core_io_CipherKey_w_178_), .D(
        top_core_io_CipherKey_w_186_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1226) );
  MX4X1 top_core_io_U1627 ( .A(top_core_io_CipherKey_w_194_), .B(
        top_core_io_CipherKey_w_202_), .C(top_core_io_CipherKey_w_210_), .D(
        top_core_io_CipherKey_w_218_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1225) );
  MX4X1 top_core_io_U1629 ( .A(top_core_io_CipherKey_w_130_), .B(
        top_core_io_CipherKey_w_138_), .C(top_core_io_CipherKey_w_146_), .D(
        top_core_io_CipherKey_w_154_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1227) );
  MX4X1 top_core_io_U1630 ( .A(top_core_io_n1227), .B(top_core_io_n1225), .C(
        top_core_io_n1226), .D(top_core_io_n1224), .S0(n4141), .S1(n4139), .Y(
        top_core_io_n1228) );
  MX4X1 top_core_io_U1617 ( .A(top_core_io_Data_reg_20__1_), .B(
        top_core_io_Data_reg_21__1_), .C(top_core_io_Data_reg_22__1_), .D(
        top_core_io_Data_reg_23__1_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1216) );
  MX4X1 top_core_io_U1616 ( .A(top_core_io_Data_reg_24__1_), .B(
        top_core_io_Data_reg_25__1_), .C(top_core_io_Data_reg_26__1_), .D(
        top_core_io_Data_reg_27__1_), .S0(n4118), .S1(n4129), .Y(
        top_core_io_n1215) );
  MX4X1 top_core_io_U1618 ( .A(top_core_io_Data_reg_16__1_), .B(
        top_core_io_Data_reg_17__1_), .C(top_core_io_Data_reg_18__1_), .D(
        top_core_io_Data_reg_19__1_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1217) );
  MX4X1 top_core_io_U1619 ( .A(top_core_io_n1217), .B(top_core_io_n1215), .C(
        top_core_io_n1216), .D(top_core_io_n1214), .S0(n4141), .S1(n4139), .Y(
        top_core_io_n1218) );
  MX4X1 top_core_io_U1638 ( .A(top_core_io_Data_reg_20__2_), .B(
        top_core_io_Data_reg_21__2_), .C(top_core_io_Data_reg_22__2_), .D(
        top_core_io_Data_reg_23__2_), .S0(n4119), .S1(n4131), .Y(
        top_core_io_n1236) );
  MX4X1 top_core_io_U1637 ( .A(top_core_io_Data_reg_24__2_), .B(
        top_core_io_Data_reg_25__2_), .C(top_core_io_Data_reg_26__2_), .D(
        top_core_io_Data_reg_27__2_), .S0(n4119), .S1(n4131), .Y(
        top_core_io_n1235) );
  MX4X1 top_core_io_U1639 ( .A(top_core_io_Data_reg_16__2_), .B(
        top_core_io_Data_reg_17__2_), .C(top_core_io_Data_reg_18__2_), .D(
        top_core_io_Data_reg_19__2_), .S0(n4119), .S1(n4131), .Y(
        top_core_io_n1237) );
  MX4X1 top_core_io_U1640 ( .A(top_core_io_n1237), .B(top_core_io_n1235), .C(
        top_core_io_n1236), .D(top_core_io_n1234), .S0(n4141), .S1(n4139), .Y(
        top_core_io_n1238) );
  MX4X1 top_core_io_U1615 ( .A(top_core_io_Data_reg_28__1_), .B(
        top_core_io_Data_reg_29__1_), .C(top_core_io_Data_reg_30__1_), .D(
        top_core_io_Data_reg_31__1_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1214) );
  MX4X1 top_core_io_U1636 ( .A(top_core_io_Data_reg_28__2_), .B(
        top_core_io_Data_reg_29__2_), .C(top_core_io_Data_reg_30__2_), .D(
        top_core_io_Data_reg_31__2_), .S0(n4119), .S1(n4131), .Y(
        top_core_io_n1234) );
  MX4X1 top_core_io_U1605 ( .A(top_core_io_CipherKey_w_225_), .B(
        top_core_io_CipherKey_w_233_), .C(top_core_io_CipherKey_w_241_), .D(
        top_core_io_CipherKey_w_249_), .S0(n4117), .S1(n4129), .Y(
        top_core_io_n1204) );
  MX4X1 top_core_io_U1626 ( .A(top_core_io_CipherKey_w_226_), .B(
        top_core_io_CipherKey_w_234_), .C(top_core_io_CipherKey_w_242_), .D(
        top_core_io_CipherKey_w_250_), .S0(n4118), .S1(n4130), .Y(
        top_core_io_n1224) );
  DFFSX1 top_core_EC_Addr_reg_0_ ( .D(top_core_EC_n1294), .CK(n3906), .SN(
        n_RSTB), .Q(top_core_Addr[0]), .QN(top_core_EC_n25) );
  DFFRHQX1 top_core_KE_key_mem_ctrl_reg_reg_0_ ( .D(top_core_KE_n4933), .CK(
        n3906), .RN(n_RSTB), .Q(top_core_KE_key_mem_ctrl_reg_0_) );
  MX4X1 top_core_io_U1656 ( .A(top_core_io_n1252), .B(top_core_io_n1250), .C(
        top_core_io_n1251), .D(top_core_io_n1249), .S0(n_ADDR[3]), .S1(n4139), 
        .Y(top_core_io_n1253) );
  MX4X1 top_core_io_U1666 ( .A(top_core_io_n1262), .B(top_core_io_n1260), .C(
        top_core_io_n1261), .D(top_core_io_n1259), .S0(n4142), .S1(n4139), .Y(
        top_core_io_n1263) );
  MX4X1 top_core_io_U1667 ( .A(top_core_io_n1263), .B(top_core_io_n1253), .C(
        top_core_io_n1258), .D(top_core_io_n1248), .S0(n_ADDR[5]), .S1(
        n_ADDR[4]), .Y(top_core_io_N78) );
  MX4X1 top_core_io_U1677 ( .A(top_core_io_n1272), .B(top_core_io_n1270), .C(
        top_core_io_n1271), .D(top_core_io_n1269), .S0(n_ADDR[3]), .S1(n4139), 
        .Y(top_core_io_n1273) );
  MX4X1 top_core_io_U1687 ( .A(top_core_io_n1282), .B(top_core_io_n1280), .C(
        top_core_io_n1281), .D(top_core_io_n1279), .S0(n_ADDR[3]), .S1(n4139), 
        .Y(top_core_io_n1283) );
  MX4X1 top_core_io_U1688 ( .A(top_core_io_n1283), .B(top_core_io_n1273), .C(
        top_core_io_n1278), .D(top_core_io_n1268), .S0(n_ADDR[5]), .S1(
        n_ADDR[4]), .Y(top_core_io_N77) );
  MX4X1 top_core_io_U1698 ( .A(top_core_io_n1292), .B(top_core_io_n1290), .C(
        top_core_io_n1291), .D(top_core_io_n1289), .S0(n_ADDR[3]), .S1(n4138), 
        .Y(top_core_io_n1293) );
  MX4X1 top_core_io_U1708 ( .A(top_core_io_n1302), .B(top_core_io_n1300), .C(
        top_core_io_n1301), .D(top_core_io_n1299), .S0(n_ADDR[3]), .S1(n4138), 
        .Y(top_core_io_n1303) );
  MX4X1 top_core_io_U1709 ( .A(top_core_io_n1303), .B(top_core_io_n1293), .C(
        top_core_io_n1298), .D(top_core_io_n1288), .S0(n_ADDR[5]), .S1(
        n_ADDR[4]), .Y(top_core_io_N76) );
  MX4X1 top_core_io_U1730 ( .A(top_core_io_n1323), .B(top_core_io_n1313), .C(
        top_core_io_n1318), .D(top_core_io_n1308), .S0(n_ADDR[5]), .S1(
        n_ADDR[4]), .Y(top_core_io_N75) );
  MX4X1 top_core_io_U1751 ( .A(top_core_io_n1343), .B(top_core_io_n1333), .C(
        top_core_io_n1338), .D(top_core_io_n1328), .S0(n_ADDR[5]), .S1(
        n_ADDR[4]), .Y(top_core_io_N74) );
  MX4X1 top_core_io_U1624 ( .A(top_core_io_n1222), .B(top_core_io_n1220), .C(
        top_core_io_n1221), .D(top_core_io_n1219), .S0(n4141), .S1(n4139), .Y(
        top_core_io_n1223) );
  MX4X1 top_core_io_U1625 ( .A(top_core_io_n1223), .B(top_core_io_n1213), .C(
        top_core_io_n1218), .D(top_core_io_n1208), .S0(n_ADDR[5]), .S1(
        n_ADDR[4]), .Y(top_core_io_N80) );
  MX4X1 top_core_io_U1645 ( .A(top_core_io_n1242), .B(top_core_io_n1240), .C(
        top_core_io_n1241), .D(top_core_io_n1239), .S0(n4141), .S1(n4139), .Y(
        top_core_io_n1243) );
  MX4X1 top_core_io_U1646 ( .A(top_core_io_n1243), .B(top_core_io_n1233), .C(
        top_core_io_n1238), .D(top_core_io_n1228), .S0(n_ADDR[5]), .S1(
        n_ADDR[4]), .Y(top_core_io_N79) );
  DFFRHQX1 top_core_io_Nk_val_reg_1_ ( .D(top_core_io_n1180), .CK(n3781), .RN(
        n_RSTB), .Q(top_core_Nk[1]) );
  DFFRHQX1 top_core_io_Nk_val_reg_2_ ( .D(top_core_io_n1179), .CK(n3769), .RN(
        n_RSTB), .Q(top_core_Nk[2]) );
  DFFRHQX1 top_core_io_Nk_val_reg_0_ ( .D(n4258), .CK(n3769), .RN(n_RSTB), .Q(
        top_core_Nk[0]) );
  DFFRHQX1 top_core_io_CipherKey_reg_0_ ( .D(top_core_io_N259), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[0]) );
  DFFRHQX1 top_core_io_CipherKey_reg_1_ ( .D(top_core_io_N260), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[1]) );
  DFFRHQX1 top_core_io_CipherKey_reg_2_ ( .D(top_core_io_N261), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[2]) );
  DFFRHQX1 top_core_io_CipherKey_reg_3_ ( .D(top_core_io_N262), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[3]) );
  DFFRHQX1 top_core_io_CipherKey_reg_4_ ( .D(top_core_io_N263), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[4]) );
  DFFRHQX1 top_core_io_CipherKey_reg_5_ ( .D(top_core_io_N264), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[5]) );
  DFFRHQX1 top_core_io_CipherKey_reg_6_ ( .D(top_core_io_N265), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[6]) );
  DFFRHQX1 top_core_io_CipherKey_reg_7_ ( .D(top_core_io_N266), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[7]) );
  DFFRHQX1 top_core_io_CipherKey_reg_8_ ( .D(top_core_io_N267), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[8]) );
  DFFRHQX1 top_core_io_CipherKey_reg_9_ ( .D(top_core_io_N268), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[9]) );
  DFFRHQX1 top_core_io_CipherKey_reg_10_ ( .D(top_core_io_N269), .CK(n3778), 
        .RN(n_RSTB), .Q(top_core_CipherKey[10]) );
  DFFRHQX1 top_core_io_CipherKey_reg_11_ ( .D(top_core_io_N270), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[11]) );
  DFFRHQX1 top_core_io_CipherKey_reg_12_ ( .D(top_core_io_N271), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[12]) );
  DFFRHQX1 top_core_io_CipherKey_reg_13_ ( .D(top_core_io_N272), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[13]) );
  DFFRHQX1 top_core_io_CipherKey_reg_14_ ( .D(top_core_io_N273), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[14]) );
  DFFRHQX1 top_core_io_CipherKey_reg_15_ ( .D(top_core_io_N274), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[15]) );
  DFFRHQX1 top_core_io_CipherKey_reg_16_ ( .D(top_core_io_N275), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[16]) );
  DFFRHQX1 top_core_io_CipherKey_reg_17_ ( .D(top_core_io_N276), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[17]) );
  DFFRHQX1 top_core_io_CipherKey_reg_18_ ( .D(top_core_io_N277), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[18]) );
  DFFRHQX1 top_core_io_CipherKey_reg_19_ ( .D(top_core_io_N278), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[19]) );
  DFFRHQX1 top_core_io_CipherKey_reg_20_ ( .D(top_core_io_N279), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[20]) );
  DFFRHQX1 top_core_io_CipherKey_reg_21_ ( .D(top_core_io_N280), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[21]) );
  DFFRHQX1 top_core_io_CipherKey_reg_22_ ( .D(top_core_io_N281), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[22]) );
  DFFRHQX1 top_core_io_CipherKey_reg_23_ ( .D(top_core_io_N282), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[23]) );
  DFFRHQX1 top_core_io_CipherKey_reg_24_ ( .D(top_core_io_N283), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[24]) );
  DFFRHQX1 top_core_io_CipherKey_reg_25_ ( .D(top_core_io_N284), .CK(n3779), 
        .RN(n_RSTB), .Q(top_core_CipherKey[25]) );
  DFFRHQX1 top_core_io_CipherKey_reg_26_ ( .D(top_core_io_N285), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[26]) );
  DFFRHQX1 top_core_io_CipherKey_reg_27_ ( .D(top_core_io_N286), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[27]) );
  DFFRHQX1 top_core_io_CipherKey_reg_28_ ( .D(top_core_io_N287), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[28]) );
  DFFRHQX1 top_core_io_CipherKey_reg_29_ ( .D(top_core_io_N288), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[29]) );
  DFFRHQX1 top_core_io_CipherKey_reg_30_ ( .D(top_core_io_N289), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[30]) );
  DFFRHQX1 top_core_io_CipherKey_reg_31_ ( .D(top_core_io_N290), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[31]) );
  DFFRHQX1 top_core_io_CipherKey_reg_32_ ( .D(top_core_io_N291), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[32]) );
  DFFRHQX1 top_core_io_CipherKey_reg_33_ ( .D(top_core_io_N292), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[33]) );
  DFFRHQX1 top_core_io_CipherKey_reg_34_ ( .D(top_core_io_N293), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[34]) );
  DFFRHQX1 top_core_io_CipherKey_reg_35_ ( .D(top_core_io_N294), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[35]) );
  DFFRHQX1 top_core_io_CipherKey_reg_36_ ( .D(top_core_io_N295), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[36]) );
  DFFRHQX1 top_core_io_CipherKey_reg_37_ ( .D(top_core_io_N296), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[37]) );
  DFFRHQX1 top_core_io_CipherKey_reg_38_ ( .D(top_core_io_N297), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[38]) );
  DFFRHQX1 top_core_io_CipherKey_reg_39_ ( .D(top_core_io_N298), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[39]) );
  DFFRHQX1 top_core_io_CipherKey_reg_40_ ( .D(top_core_io_N299), .CK(n3780), 
        .RN(n_RSTB), .Q(top_core_CipherKey[40]) );
  DFFRHQX1 top_core_io_CipherKey_reg_41_ ( .D(top_core_io_N300), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[41]) );
  DFFRHQX1 top_core_io_CipherKey_reg_42_ ( .D(top_core_io_N301), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[42]) );
  DFFRHQX1 top_core_io_CipherKey_reg_43_ ( .D(top_core_io_N302), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[43]) );
  DFFRHQX1 top_core_io_CipherKey_reg_44_ ( .D(top_core_io_N303), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[44]) );
  DFFRHQX1 top_core_io_CipherKey_reg_45_ ( .D(top_core_io_N304), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[45]) );
  DFFRHQX1 top_core_io_CipherKey_reg_46_ ( .D(top_core_io_N305), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[46]) );
  DFFRHQX1 top_core_io_CipherKey_reg_47_ ( .D(top_core_io_N306), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[47]) );
  DFFRHQX1 top_core_io_CipherKey_reg_48_ ( .D(top_core_io_N307), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[48]) );
  DFFRHQX1 top_core_io_CipherKey_reg_49_ ( .D(top_core_io_N308), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[49]) );
  DFFRHQX1 top_core_io_CipherKey_reg_50_ ( .D(top_core_io_N309), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[50]) );
  DFFRHQX1 top_core_io_CipherKey_reg_51_ ( .D(top_core_io_N310), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[51]) );
  DFFRHQX1 top_core_io_CipherKey_reg_52_ ( .D(top_core_io_N311), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[52]) );
  DFFRHQX1 top_core_io_CipherKey_reg_53_ ( .D(top_core_io_N312), .CK(n3781), 
        .RN(n_RSTB), .Q(top_core_CipherKey[53]) );
  DFFRHQX1 top_core_io_CipherKey_reg_54_ ( .D(top_core_io_N313), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[54]) );
  DFFRHQX1 top_core_io_CipherKey_reg_55_ ( .D(top_core_io_N314), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[55]) );
  DFFRHQX1 top_core_io_CipherKey_reg_56_ ( .D(top_core_io_N315), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[56]) );
  DFFRHQX1 top_core_io_CipherKey_reg_57_ ( .D(top_core_io_N316), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[57]) );
  DFFRHQX1 top_core_io_CipherKey_reg_58_ ( .D(top_core_io_N317), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[58]) );
  DFFRHQX1 top_core_io_CipherKey_reg_59_ ( .D(top_core_io_N318), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[59]) );
  DFFRHQX1 top_core_io_CipherKey_reg_60_ ( .D(top_core_io_N319), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[60]) );
  DFFRHQX1 top_core_io_CipherKey_reg_61_ ( .D(top_core_io_N320), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[61]) );
  DFFRHQX1 top_core_io_CipherKey_reg_62_ ( .D(top_core_io_N321), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[62]) );
  DFFRHQX1 top_core_io_CipherKey_reg_63_ ( .D(top_core_io_N322), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[63]) );
  DFFRHQX1 top_core_io_CipherKey_reg_64_ ( .D(top_core_io_N323), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[64]) );
  DFFRHQX1 top_core_io_CipherKey_reg_65_ ( .D(top_core_io_N324), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[65]) );
  DFFRHQX1 top_core_io_CipherKey_reg_66_ ( .D(top_core_io_N325), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[66]) );
  DFFRHQX1 top_core_io_CipherKey_reg_67_ ( .D(top_core_io_N326), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[67]) );
  DFFRHQX1 top_core_io_CipherKey_reg_68_ ( .D(top_core_io_N327), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[68]) );
  DFFRHQX1 top_core_io_CipherKey_reg_69_ ( .D(top_core_io_N328), .CK(n3757), 
        .RN(n_RSTB), .Q(top_core_CipherKey[69]) );
  DFFRHQX1 top_core_io_CipherKey_reg_70_ ( .D(top_core_io_N329), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[70]) );
  DFFRHQX1 top_core_io_CipherKey_reg_71_ ( .D(top_core_io_N330), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[71]) );
  DFFRHQX1 top_core_io_CipherKey_reg_72_ ( .D(top_core_io_N331), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[72]) );
  DFFRHQX1 top_core_io_CipherKey_reg_73_ ( .D(top_core_io_N332), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[73]) );
  DFFRHQX1 top_core_io_CipherKey_reg_74_ ( .D(top_core_io_N333), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[74]) );
  DFFRHQX1 top_core_io_CipherKey_reg_75_ ( .D(top_core_io_N334), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[75]) );
  DFFRHQX1 top_core_io_CipherKey_reg_76_ ( .D(top_core_io_N335), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[76]) );
  DFFRHQX1 top_core_io_CipherKey_reg_77_ ( .D(top_core_io_N336), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[77]) );
  DFFRHQX1 top_core_io_CipherKey_reg_78_ ( .D(top_core_io_N337), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[78]) );
  DFFRHQX1 top_core_io_CipherKey_reg_79_ ( .D(top_core_io_N338), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[79]) );
  DFFRHQX1 top_core_io_CipherKey_reg_80_ ( .D(top_core_io_N339), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[80]) );
  DFFRHQX1 top_core_io_CipherKey_reg_81_ ( .D(top_core_io_N340), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[81]) );
  DFFRHQX1 top_core_io_CipherKey_reg_82_ ( .D(top_core_io_N341), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[82]) );
  DFFRHQX1 top_core_io_CipherKey_reg_83_ ( .D(top_core_io_N342), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[83]) );
  DFFRHQX1 top_core_io_CipherKey_reg_84_ ( .D(top_core_io_N343), .CK(n3758), 
        .RN(n_RSTB), .Q(top_core_CipherKey[84]) );
  DFFRHQX1 top_core_io_CipherKey_reg_85_ ( .D(top_core_io_N344), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[85]) );
  DFFRHQX1 top_core_io_CipherKey_reg_86_ ( .D(top_core_io_N345), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[86]) );
  DFFRHQX1 top_core_io_CipherKey_reg_87_ ( .D(top_core_io_N346), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[87]) );
  DFFRHQX1 top_core_io_CipherKey_reg_88_ ( .D(top_core_io_N347), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[88]) );
  DFFRHQX1 top_core_io_CipherKey_reg_89_ ( .D(top_core_io_N348), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[89]) );
  DFFRHQX1 top_core_io_CipherKey_reg_90_ ( .D(top_core_io_N349), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[90]) );
  DFFRHQX1 top_core_io_CipherKey_reg_91_ ( .D(top_core_io_N350), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[91]) );
  DFFRHQX1 top_core_io_CipherKey_reg_92_ ( .D(top_core_io_N351), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[92]) );
  DFFRHQX1 top_core_io_CipherKey_reg_93_ ( .D(top_core_io_N352), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[93]) );
  DFFRHQX1 top_core_io_CipherKey_reg_94_ ( .D(top_core_io_N353), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[94]) );
  DFFRHQX1 top_core_io_CipherKey_reg_95_ ( .D(top_core_io_N354), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[95]) );
  DFFRHQX1 top_core_io_CipherKey_reg_96_ ( .D(top_core_io_N355), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[96]) );
  DFFRHQX1 top_core_io_CipherKey_reg_97_ ( .D(top_core_io_N356), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[97]) );
  DFFRHQX1 top_core_io_CipherKey_reg_98_ ( .D(top_core_io_N357), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[98]) );
  DFFRHQX1 top_core_io_CipherKey_reg_99_ ( .D(top_core_io_N358), .CK(n3759), 
        .RN(n_RSTB), .Q(top_core_CipherKey[99]) );
  DFFRHQX1 top_core_io_CipherKey_reg_100_ ( .D(top_core_io_N359), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[100]) );
  DFFRHQX1 top_core_io_CipherKey_reg_101_ ( .D(top_core_io_N360), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[101]) );
  DFFRHQX1 top_core_io_CipherKey_reg_102_ ( .D(top_core_io_N361), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[102]) );
  DFFRHQX1 top_core_io_CipherKey_reg_103_ ( .D(top_core_io_N362), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[103]) );
  DFFRHQX1 top_core_io_CipherKey_reg_104_ ( .D(top_core_io_N363), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[104]) );
  DFFRHQX1 top_core_io_CipherKey_reg_105_ ( .D(top_core_io_N364), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[105]) );
  DFFRHQX1 top_core_io_CipherKey_reg_106_ ( .D(top_core_io_N365), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[106]) );
  DFFRHQX1 top_core_io_CipherKey_reg_107_ ( .D(top_core_io_N366), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[107]) );
  DFFRHQX1 top_core_io_CipherKey_reg_108_ ( .D(top_core_io_N367), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[108]) );
  DFFRHQX1 top_core_io_CipherKey_reg_109_ ( .D(top_core_io_N368), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[109]) );
  DFFRHQX1 top_core_io_CipherKey_reg_110_ ( .D(top_core_io_N369), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[110]) );
  DFFRHQX1 top_core_io_CipherKey_reg_111_ ( .D(top_core_io_N370), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[111]) );
  DFFRHQX1 top_core_io_CipherKey_reg_112_ ( .D(top_core_io_N371), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[112]) );
  DFFRHQX1 top_core_io_CipherKey_reg_113_ ( .D(top_core_io_N372), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[113]) );
  DFFRHQX1 top_core_io_CipherKey_reg_114_ ( .D(top_core_io_N373), .CK(n3760), 
        .RN(n_RSTB), .Q(top_core_CipherKey[114]) );
  DFFRHQX1 top_core_io_CipherKey_reg_115_ ( .D(top_core_io_N374), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[115]) );
  DFFRHQX1 top_core_io_CipherKey_reg_116_ ( .D(top_core_io_N375), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[116]) );
  DFFRHQX1 top_core_io_CipherKey_reg_117_ ( .D(top_core_io_N376), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[117]) );
  DFFRHQX1 top_core_io_CipherKey_reg_118_ ( .D(top_core_io_N377), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[118]) );
  DFFRHQX1 top_core_io_CipherKey_reg_119_ ( .D(top_core_io_N378), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[119]) );
  DFFRHQX1 top_core_io_CipherKey_reg_120_ ( .D(top_core_io_N379), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[120]) );
  DFFRHQX1 top_core_io_CipherKey_reg_121_ ( .D(top_core_io_N380), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[121]) );
  DFFRHQX1 top_core_io_CipherKey_reg_122_ ( .D(top_core_io_N381), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[122]) );
  DFFRHQX1 top_core_io_CipherKey_reg_123_ ( .D(top_core_io_N382), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[123]) );
  DFFRHQX1 top_core_io_CipherKey_reg_124_ ( .D(top_core_io_N383), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[124]) );
  DFFRHQX1 top_core_io_CipherKey_reg_125_ ( .D(top_core_io_N384), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[125]) );
  DFFRHQX1 top_core_io_CipherKey_reg_126_ ( .D(top_core_io_N385), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[126]) );
  DFFRHQX1 top_core_io_CipherKey_reg_127_ ( .D(top_core_io_N386), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[127]) );
  DFFRHQX1 top_core_io_CipherKey_reg_128_ ( .D(top_core_io_N387), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[128]) );
  DFFRHQX1 top_core_io_CipherKey_reg_129_ ( .D(top_core_io_N388), .CK(n3761), 
        .RN(n_RSTB), .Q(top_core_CipherKey[129]) );
  DFFRHQX1 top_core_io_CipherKey_reg_130_ ( .D(top_core_io_N389), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[130]) );
  DFFRHQX1 top_core_io_CipherKey_reg_131_ ( .D(top_core_io_N390), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[131]) );
  DFFRHQX1 top_core_io_CipherKey_reg_132_ ( .D(top_core_io_N391), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[132]) );
  DFFRHQX1 top_core_io_CipherKey_reg_133_ ( .D(top_core_io_N392), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[133]) );
  DFFRHQX1 top_core_io_CipherKey_reg_134_ ( .D(top_core_io_N393), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[134]) );
  DFFRHQX1 top_core_io_CipherKey_reg_135_ ( .D(top_core_io_N394), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[135]) );
  DFFRHQX1 top_core_io_CipherKey_reg_136_ ( .D(top_core_io_N395), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[136]) );
  DFFRHQX1 top_core_io_CipherKey_reg_137_ ( .D(top_core_io_N396), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[137]) );
  DFFRHQX1 top_core_io_CipherKey_reg_138_ ( .D(top_core_io_N397), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[138]) );
  DFFRHQX1 top_core_io_CipherKey_reg_139_ ( .D(top_core_io_N398), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[139]) );
  DFFRHQX1 top_core_io_CipherKey_reg_140_ ( .D(top_core_io_N399), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[140]) );
  DFFRHQX1 top_core_io_CipherKey_reg_141_ ( .D(top_core_io_N400), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[141]) );
  DFFRHQX1 top_core_io_CipherKey_reg_142_ ( .D(top_core_io_N401), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[142]) );
  DFFRHQX1 top_core_io_CipherKey_reg_143_ ( .D(top_core_io_N402), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[143]) );
  DFFRHQX1 top_core_io_CipherKey_reg_144_ ( .D(top_core_io_N403), .CK(n3762), 
        .RN(n_RSTB), .Q(top_core_CipherKey[144]) );
  DFFRHQX1 top_core_io_CipherKey_reg_145_ ( .D(top_core_io_N404), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[145]) );
  DFFRHQX1 top_core_io_CipherKey_reg_146_ ( .D(top_core_io_N405), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[146]) );
  DFFRHQX1 top_core_io_CipherKey_reg_147_ ( .D(top_core_io_N406), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[147]) );
  DFFRHQX1 top_core_io_CipherKey_reg_148_ ( .D(top_core_io_N407), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[148]) );
  DFFRHQX1 top_core_io_CipherKey_reg_149_ ( .D(top_core_io_N408), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[149]) );
  DFFRHQX1 top_core_io_CipherKey_reg_150_ ( .D(top_core_io_N409), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[150]) );
  DFFRHQX1 top_core_io_CipherKey_reg_151_ ( .D(top_core_io_N410), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[151]) );
  DFFRHQX1 top_core_io_CipherKey_reg_152_ ( .D(top_core_io_N411), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[152]) );
  DFFRHQX1 top_core_io_CipherKey_reg_153_ ( .D(top_core_io_N412), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[153]) );
  DFFRHQX1 top_core_io_CipherKey_reg_154_ ( .D(top_core_io_N413), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[154]) );
  DFFRHQX1 top_core_io_CipherKey_reg_155_ ( .D(top_core_io_N414), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[155]) );
  DFFRHQX1 top_core_io_CipherKey_reg_156_ ( .D(top_core_io_N415), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[156]) );
  DFFRHQX1 top_core_io_CipherKey_reg_157_ ( .D(top_core_io_N416), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[157]) );
  DFFRHQX1 top_core_io_CipherKey_reg_158_ ( .D(top_core_io_N417), .CK(n3763), 
        .RN(n_RSTB), .Q(top_core_CipherKey[158]) );
  DFFRHQX1 top_core_io_CipherKey_reg_159_ ( .D(top_core_io_N418), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[159]) );
  DFFRHQX1 top_core_io_CipherKey_reg_160_ ( .D(top_core_io_N419), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[160]) );
  DFFRHQX1 top_core_io_CipherKey_reg_161_ ( .D(top_core_io_N420), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[161]) );
  DFFRHQX1 top_core_io_CipherKey_reg_162_ ( .D(top_core_io_N421), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[162]) );
  DFFRHQX1 top_core_io_CipherKey_reg_163_ ( .D(top_core_io_N422), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[163]) );
  DFFRHQX1 top_core_io_CipherKey_reg_164_ ( .D(top_core_io_N423), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[164]) );
  DFFRHQX1 top_core_io_CipherKey_reg_165_ ( .D(top_core_io_N424), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[165]) );
  DFFRHQX1 top_core_io_CipherKey_reg_166_ ( .D(top_core_io_N425), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[166]) );
  DFFRHQX1 top_core_io_CipherKey_reg_167_ ( .D(top_core_io_N426), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[167]) );
  DFFRHQX1 top_core_io_CipherKey_reg_168_ ( .D(top_core_io_N427), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[168]) );
  DFFRHQX1 top_core_io_CipherKey_reg_169_ ( .D(top_core_io_N428), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[169]) );
  DFFRHQX1 top_core_io_CipherKey_reg_170_ ( .D(top_core_io_N429), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[170]) );
  DFFRHQX1 top_core_io_CipherKey_reg_171_ ( .D(top_core_io_N430), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[171]) );
  DFFRHQX1 top_core_io_CipherKey_reg_172_ ( .D(top_core_io_N431), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[172]) );
  DFFRHQX1 top_core_io_CipherKey_reg_173_ ( .D(top_core_io_N432), .CK(n3764), 
        .RN(n_RSTB), .Q(top_core_CipherKey[173]) );
  DFFRHQX1 top_core_io_CipherKey_reg_174_ ( .D(top_core_io_N433), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[174]) );
  DFFRHQX1 top_core_io_CipherKey_reg_175_ ( .D(top_core_io_N434), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[175]) );
  DFFRHQX1 top_core_io_CipherKey_reg_176_ ( .D(top_core_io_N435), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[176]) );
  DFFRHQX1 top_core_io_CipherKey_reg_177_ ( .D(top_core_io_N436), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[177]) );
  DFFRHQX1 top_core_io_CipherKey_reg_178_ ( .D(top_core_io_N437), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[178]) );
  DFFRHQX1 top_core_io_CipherKey_reg_179_ ( .D(top_core_io_N438), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[179]) );
  DFFRHQX1 top_core_io_CipherKey_reg_180_ ( .D(top_core_io_N439), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[180]) );
  DFFRHQX1 top_core_io_CipherKey_reg_181_ ( .D(top_core_io_N440), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[181]) );
  DFFRHQX1 top_core_io_CipherKey_reg_182_ ( .D(top_core_io_N441), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[182]) );
  DFFRHQX1 top_core_io_CipherKey_reg_183_ ( .D(top_core_io_N442), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[183]) );
  DFFRHQX1 top_core_io_CipherKey_reg_184_ ( .D(top_core_io_N443), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[184]) );
  DFFRHQX1 top_core_io_CipherKey_reg_185_ ( .D(top_core_io_N444), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[185]) );
  DFFRHQX1 top_core_io_CipherKey_reg_186_ ( .D(top_core_io_N445), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[186]) );
  DFFRHQX1 top_core_io_CipherKey_reg_187_ ( .D(top_core_io_N446), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[187]) );
  DFFRHQX1 top_core_io_CipherKey_reg_188_ ( .D(top_core_io_N447), .CK(n3765), 
        .RN(n_RSTB), .Q(top_core_CipherKey[188]) );
  DFFRHQX1 top_core_io_CipherKey_reg_189_ ( .D(top_core_io_N448), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[189]) );
  DFFRHQX1 top_core_io_CipherKey_reg_190_ ( .D(top_core_io_N449), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[190]) );
  DFFRHQX1 top_core_io_CipherKey_reg_191_ ( .D(top_core_io_N450), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[191]) );
  DFFRHQX1 top_core_io_CipherKey_reg_192_ ( .D(top_core_io_N451), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[192]) );
  DFFRHQX1 top_core_io_CipherKey_reg_193_ ( .D(top_core_io_N452), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[193]) );
  DFFRHQX1 top_core_io_CipherKey_reg_194_ ( .D(top_core_io_N453), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[194]) );
  DFFRHQX1 top_core_io_CipherKey_reg_195_ ( .D(top_core_io_N454), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[195]) );
  DFFRHQX1 top_core_io_CipherKey_reg_196_ ( .D(top_core_io_N455), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[196]) );
  DFFRHQX1 top_core_io_CipherKey_reg_197_ ( .D(top_core_io_N456), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[197]) );
  DFFRHQX1 top_core_io_CipherKey_reg_198_ ( .D(top_core_io_N457), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[198]) );
  DFFRHQX1 top_core_io_CipherKey_reg_199_ ( .D(top_core_io_N458), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[199]) );
  DFFRHQX1 top_core_io_CipherKey_reg_200_ ( .D(top_core_io_N459), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[200]) );
  DFFRHQX1 top_core_io_CipherKey_reg_201_ ( .D(top_core_io_N460), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[201]) );
  DFFRHQX1 top_core_io_CipherKey_reg_202_ ( .D(top_core_io_N461), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[202]) );
  DFFRHQX1 top_core_io_CipherKey_reg_203_ ( .D(top_core_io_N462), .CK(n3766), 
        .RN(n_RSTB), .Q(top_core_CipherKey[203]) );
  DFFRHQX1 top_core_io_CipherKey_reg_204_ ( .D(top_core_io_N463), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[204]) );
  DFFRHQX1 top_core_io_CipherKey_reg_205_ ( .D(top_core_io_N464), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[205]) );
  DFFRHQX1 top_core_io_CipherKey_reg_206_ ( .D(top_core_io_N465), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[206]) );
  DFFRHQX1 top_core_io_CipherKey_reg_207_ ( .D(top_core_io_N466), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[207]) );
  DFFRHQX1 top_core_io_CipherKey_reg_208_ ( .D(top_core_io_N467), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[208]) );
  DFFRHQX1 top_core_io_CipherKey_reg_209_ ( .D(top_core_io_N468), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[209]) );
  DFFRHQX1 top_core_io_CipherKey_reg_210_ ( .D(top_core_io_N469), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[210]) );
  DFFRHQX1 top_core_io_CipherKey_reg_211_ ( .D(top_core_io_N470), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[211]) );
  DFFRHQX1 top_core_io_CipherKey_reg_212_ ( .D(top_core_io_N471), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[212]) );
  DFFRHQX1 top_core_io_CipherKey_reg_213_ ( .D(top_core_io_N472), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[213]) );
  DFFRHQX1 top_core_io_CipherKey_reg_214_ ( .D(top_core_io_N473), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[214]) );
  DFFRHQX1 top_core_io_CipherKey_reg_215_ ( .D(top_core_io_N474), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[215]) );
  DFFRHQX1 top_core_io_CipherKey_reg_216_ ( .D(top_core_io_N475), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[216]) );
  DFFRHQX1 top_core_io_CipherKey_reg_217_ ( .D(top_core_io_N476), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[217]) );
  DFFRHQX1 top_core_io_CipherKey_reg_218_ ( .D(top_core_io_N477), .CK(n3767), 
        .RN(n_RSTB), .Q(top_core_CipherKey[218]) );
  DFFRHQX1 top_core_io_CipherKey_reg_219_ ( .D(top_core_io_N478), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[219]) );
  DFFRHQX1 top_core_io_CipherKey_reg_220_ ( .D(top_core_io_N479), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[220]) );
  DFFRHQX1 top_core_io_CipherKey_reg_221_ ( .D(top_core_io_N480), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[221]) );
  DFFRHQX1 top_core_io_CipherKey_reg_222_ ( .D(top_core_io_N481), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[222]) );
  DFFRHQX1 top_core_io_CipherKey_reg_223_ ( .D(top_core_io_N482), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[223]) );
  DFFRHQX1 top_core_io_CipherKey_reg_224_ ( .D(top_core_io_N483), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[224]) );
  DFFRHQX1 top_core_io_CipherKey_reg_225_ ( .D(top_core_io_N484), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[225]) );
  DFFRHQX1 top_core_io_CipherKey_reg_226_ ( .D(top_core_io_N485), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[226]) );
  DFFRHQX1 top_core_io_CipherKey_reg_227_ ( .D(top_core_io_N486), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[227]) );
  DFFRHQX1 top_core_io_CipherKey_reg_228_ ( .D(top_core_io_N487), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[228]) );
  DFFRHQX1 top_core_io_CipherKey_reg_229_ ( .D(top_core_io_N488), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[229]) );
  DFFRHQX1 top_core_io_CipherKey_reg_230_ ( .D(top_core_io_N489), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[230]) );
  DFFRHQX1 top_core_io_CipherKey_reg_231_ ( .D(top_core_io_N490), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[231]) );
  DFFRHQX1 top_core_io_CipherKey_reg_232_ ( .D(top_core_io_N491), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[232]) );
  DFFRHQX1 top_core_io_CipherKey_reg_233_ ( .D(top_core_io_N492), .CK(n3768), 
        .RN(n_RSTB), .Q(top_core_CipherKey[233]) );
  DFFRHQX1 top_core_io_CipherKey_reg_234_ ( .D(top_core_io_N493), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_CipherKey[234]) );
  DFFRHQX1 top_core_io_CipherKey_reg_235_ ( .D(top_core_io_N494), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_CipherKey[235]) );
  DFFRHQX1 top_core_io_CipherKey_reg_236_ ( .D(top_core_io_N495), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_CipherKey[236]) );
  DFFRHQX1 top_core_io_CipherKey_reg_237_ ( .D(top_core_io_N496), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_CipherKey[237]) );
  DFFRHQX1 top_core_io_CipherKey_reg_238_ ( .D(top_core_io_N497), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_CipherKey[238]) );
  DFFRHQX1 top_core_io_CipherKey_reg_239_ ( .D(top_core_io_N498), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_CipherKey[239]) );
  DFFRHQX1 top_core_io_CipherKey_reg_240_ ( .D(top_core_io_N499), .CK(n3769), 
        .RN(n_RSTB), .Q(top_core_CipherKey[240]) );
  DFFRHQX1 top_core_io_CipherKey_reg_241_ ( .D(top_core_io_N500), .CK(n3800), 
        .RN(n_RSTB), .Q(top_core_CipherKey[241]) );
  DFFRHQX1 top_core_io_CipherKey_reg_242_ ( .D(top_core_io_N501), .CK(n3794), 
        .RN(n_RSTB), .Q(top_core_CipherKey[242]) );
  DFFRHQX1 top_core_io_CipherKey_reg_243_ ( .D(top_core_io_N502), .CK(n3794), 
        .RN(n_RSTB), .Q(top_core_CipherKey[243]) );
  DFFRHQX1 top_core_io_CipherKey_reg_244_ ( .D(top_core_io_N503), .CK(n3794), 
        .RN(n_RSTB), .Q(top_core_CipherKey[244]) );
  DFFRHQX1 top_core_io_CipherKey_reg_245_ ( .D(top_core_io_N504), .CK(n3794), 
        .RN(n_RSTB), .Q(top_core_CipherKey[245]) );
  DFFRHQX1 top_core_io_CipherKey_reg_246_ ( .D(top_core_io_N505), .CK(n3794), 
        .RN(n_RSTB), .Q(top_core_CipherKey[246]) );
  DFFRHQX1 top_core_io_CipherKey_reg_247_ ( .D(top_core_io_N506), .CK(n3794), 
        .RN(n_RSTB), .Q(top_core_CipherKey[247]) );
  DFFRHQX1 top_core_io_CipherKey_reg_248_ ( .D(top_core_io_N507), .CK(n3794), 
        .RN(n_RSTB), .Q(top_core_CipherKey[248]) );
  DFFRHQX1 top_core_io_CipherKey_reg_249_ ( .D(top_core_io_N508), .CK(n3794), 
        .RN(n_RSTB), .Q(top_core_CipherKey[249]) );
  DFFRHQX1 top_core_io_CipherKey_reg_250_ ( .D(top_core_io_N509), .CK(n3794), 
        .RN(n_RSTB), .Q(top_core_CipherKey[250]) );
  DFFRHQX1 top_core_io_CipherKey_reg_251_ ( .D(top_core_io_N510), .CK(n3795), 
        .RN(n_RSTB), .Q(top_core_CipherKey[251]) );
  DFFRHQX1 top_core_io_CipherKey_reg_252_ ( .D(top_core_io_N511), .CK(n3795), 
        .RN(n_RSTB), .Q(top_core_CipherKey[252]) );
  DFFRHQX1 top_core_io_CipherKey_reg_253_ ( .D(top_core_io_N512), .CK(n3795), 
        .RN(n_RSTB), .Q(top_core_CipherKey[253]) );
  DFFRHQX1 top_core_io_CipherKey_reg_254_ ( .D(top_core_io_N513), .CK(n3795), 
        .RN(n_RSTB), .Q(top_core_CipherKey[254]) );
  DFFRHQX1 top_core_io_CipherKey_reg_255_ ( .D(top_core_io_N514), .CK(n3795), 
        .RN(n_RSTB), .Q(top_core_CipherKey[255]) );
  MX4XL top_core_io_U1740 ( .A(top_core_io_n1332), .B(top_core_io_n1330), .C(
        top_core_io_n1331), .D(top_core_io_n1329), .S0(n4142), .S1(n4138), .Y(
        top_core_io_n1333) );
  MX4XL top_core_io_U1724 ( .A(top_core_io_n1317), .B(top_core_io_n1315), .C(
        top_core_io_n1316), .D(top_core_io_n1314), .S0(n4142), .S1(n4138), .Y(
        top_core_io_n1318) );
  MX4XL top_core_io_U1714 ( .A(top_core_io_n1307), .B(top_core_io_n1305), .C(
        top_core_io_n1306), .D(top_core_io_n1304), .S0(n4142), .S1(n4138), .Y(
        top_core_io_n1308) );
  MX4XL top_core_io_U1735 ( .A(top_core_io_n1327), .B(top_core_io_n1325), .C(
        top_core_io_n1326), .D(top_core_io_n1324), .S0(n4142), .S1(n4138), .Y(
        top_core_io_n1328) );
  MX4XL top_core_io_U1719 ( .A(top_core_io_n1312), .B(top_core_io_n1310), .C(
        top_core_io_n1311), .D(top_core_io_n1309), .S0(n4142), .S1(n4138), .Y(
        top_core_io_n1313) );
  MX4XL top_core_io_U1729 ( .A(top_core_io_n1322), .B(top_core_io_n1320), .C(
        top_core_io_n1321), .D(top_core_io_n1319), .S0(n4142), .S1(n4138), .Y(
        top_core_io_n1323) );
  MX4XL top_core_io_U1745 ( .A(top_core_io_n1337), .B(top_core_io_n1335), .C(
        top_core_io_n1336), .D(top_core_io_n1334), .S0(n4142), .S1(n4138), .Y(
        top_core_io_n1338) );
  MX4XL top_core_io_U1750 ( .A(top_core_io_n1342), .B(top_core_io_n1340), .C(
        top_core_io_n1341), .D(top_core_io_n1339), .S0(n4142), .S1(n4138), .Y(
        top_core_io_n1343) );
  MX4XL top_core_io_U1591 ( .A(top_core_io_CipherKey_w_32_), .B(
        top_core_io_CipherKey_w_40_), .C(top_core_io_CipherKey_w_48_), .D(
        top_core_io_CipherKey_w_56_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1191) );
  MX4XL top_core_io_U1590 ( .A(top_core_io_CipherKey_w_64_), .B(
        top_core_io_CipherKey_w_72_), .C(top_core_io_CipherKey_w_80_), .D(
        top_core_io_CipherKey_w_88_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1190) );
  MX4XL top_core_io_U1592 ( .A(top_core_io_CipherKey_w_0_), .B(
        top_core_io_CipherKey_w_8_), .C(top_core_io_CipherKey_w_16_), .D(
        top_core_io_CipherKey_w_24_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1192) );
  MX4XL top_core_io_U1596 ( .A(top_core_io_Data_reg_20__0_), .B(
        top_core_io_Data_reg_21__0_), .C(top_core_io_Data_reg_22__0_), .D(
        top_core_io_Data_reg_23__0_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1196) );
  MX4XL top_core_io_U1595 ( .A(top_core_io_Data_reg_24__0_), .B(
        top_core_io_Data_reg_25__0_), .C(top_core_io_Data_reg_26__0_), .D(
        top_core_io_Data_reg_27__0_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1195) );
  MX4XL top_core_io_U1597 ( .A(top_core_io_Data_reg_16__0_), .B(
        top_core_io_Data_reg_17__0_), .C(top_core_io_Data_reg_18__0_), .D(
        top_core_io_Data_reg_19__0_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1197) );
  MX4XL top_core_io_U1586 ( .A(top_core_io_CipherKey_w_160_), .B(
        top_core_io_CipherKey_w_168_), .C(top_core_io_CipherKey_w_176_), .D(
        top_core_io_CipherKey_w_184_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1186) );
  MX4XL top_core_io_U1585 ( .A(top_core_io_CipherKey_w_192_), .B(
        top_core_io_CipherKey_w_200_), .C(top_core_io_CipherKey_w_208_), .D(
        top_core_io_CipherKey_w_216_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1185) );
  MX4XL top_core_io_U1587 ( .A(top_core_io_CipherKey_w_128_), .B(
        top_core_io_CipherKey_w_136_), .C(top_core_io_CipherKey_w_144_), .D(
        top_core_io_CipherKey_w_152_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1187) );
  MX4XL top_core_io_U1589 ( .A(top_core_io_CipherKey_w_96_), .B(
        top_core_io_CipherKey_w_104_), .C(top_core_io_CipherKey_w_112_), .D(
        top_core_io_CipherKey_w_120_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1189) );
  MX4XL top_core_io_U1594 ( .A(top_core_io_Data_reg_28__0_), .B(
        top_core_io_Data_reg_29__0_), .C(top_core_io_Data_reg_30__0_), .D(
        top_core_io_Data_reg_31__0_), .S0(n4116), .S1(n4128), .Y(
        top_core_io_n1194) );
  DFFRX1 top_core_io_NK_reg_0_ ( .D(top_core_io_n664), .CK(n_CLK), .RN(n_RSTB), 
        .Q(top_core_io_NK_0_) );
  DFFRX1 top_core_io_Data_reg_reg_7__7_ ( .D(top_core_io_n1122), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_63_), .QN(n4718) );
  DFFRX1 top_core_io_Data_reg_reg_7__6_ ( .D(top_core_io_n1121), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_62_), .QN(n4717) );
  DFFRX1 top_core_io_Data_reg_reg_7__5_ ( .D(top_core_io_n1120), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_61_), .QN(n4716) );
  DFFRX1 top_core_io_Data_reg_reg_7__4_ ( .D(top_core_io_n1119), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_60_), .QN(n4715) );
  DFFRX1 top_core_io_Data_reg_reg_7__3_ ( .D(top_core_io_n1118), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_59_), .QN(n4714) );
  DFFRX1 top_core_io_Data_reg_reg_7__2_ ( .D(top_core_io_n1117), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_58_), .QN(n4713) );
  DFFRX1 top_core_io_Data_reg_reg_7__1_ ( .D(top_core_io_n1116), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_57_), .QN(n4712) );
  DFFRX1 top_core_io_Data_reg_reg_7__0_ ( .D(top_core_io_n1115), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_56_), .QN(n4711) );
  DFFRX1 top_core_io_Data_reg_reg_55__7_ ( .D(top_core_io_n738), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_191_), .QN(n4334) );
  DFFRX1 top_core_io_Data_reg_reg_55__6_ ( .D(top_core_io_n737), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_190_), .QN(n4333) );
  DFFRX1 top_core_io_Data_reg_reg_55__5_ ( .D(top_core_io_n736), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_189_), .QN(n4332) );
  DFFRX1 top_core_io_Data_reg_reg_55__4_ ( .D(top_core_io_n735), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_188_), .QN(n4331) );
  DFFRX1 top_core_io_Data_reg_reg_55__3_ ( .D(top_core_io_n734), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_187_), .QN(n4330) );
  DFFRX1 top_core_io_Data_reg_reg_55__2_ ( .D(top_core_io_n733), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_186_), .QN(n4329) );
  DFFRX1 top_core_io_Data_reg_reg_55__1_ ( .D(top_core_io_n732), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_185_), .QN(n4328) );
  DFFRX1 top_core_io_Data_reg_reg_55__0_ ( .D(top_core_io_n731), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_184_), .QN(n4327) );
  DFFRX1 top_core_io_Data_reg_reg_3__7_ ( .D(top_core_io_n1154), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_31_), .QN(n4750) );
  DFFRX1 top_core_io_Data_reg_reg_3__6_ ( .D(top_core_io_n1153), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_30_), .QN(n4749) );
  DFFRX1 top_core_io_Data_reg_reg_3__5_ ( .D(top_core_io_n1152), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_29_), .QN(n4748) );
  DFFRX1 top_core_io_Data_reg_reg_3__4_ ( .D(top_core_io_n1151), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_28_), .QN(n4747) );
  DFFRX1 top_core_io_Data_reg_reg_3__3_ ( .D(top_core_io_n1150), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_27_), .QN(n4746) );
  DFFRX1 top_core_io_Data_reg_reg_3__2_ ( .D(top_core_io_n1149), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_26_), .QN(n4745) );
  DFFRX1 top_core_io_Data_reg_reg_3__1_ ( .D(top_core_io_n1148), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_25_), .QN(n4744) );
  DFFRX1 top_core_io_Data_reg_reg_3__0_ ( .D(top_core_io_n1147), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_24_), .QN(n4743) );
  DFFRX1 top_core_io_Data_reg_reg_51__7_ ( .D(top_core_io_n770), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_159_), .QN(n4366) );
  DFFRX1 top_core_io_Data_reg_reg_51__6_ ( .D(top_core_io_n769), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_158_), .QN(n4365) );
  DFFRX1 top_core_io_Data_reg_reg_51__5_ ( .D(top_core_io_n768), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_157_), .QN(n4364) );
  DFFRX1 top_core_io_Data_reg_reg_51__4_ ( .D(top_core_io_n767), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_156_), .QN(n4363) );
  DFFRX1 top_core_io_Data_reg_reg_51__3_ ( .D(top_core_io_n766), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_155_), .QN(n4362) );
  DFFRX1 top_core_io_Data_reg_reg_51__2_ ( .D(top_core_io_n765), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_154_), .QN(n4361) );
  DFFRX1 top_core_io_Data_reg_reg_51__1_ ( .D(top_core_io_n764), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_153_), .QN(n4360) );
  DFFRX1 top_core_io_Data_reg_reg_51__0_ ( .D(top_core_io_n763), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_152_), .QN(n4359) );
  DFFRX1 top_core_io_Data_reg_reg_35__7_ ( .D(top_core_io_n898), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_31_), .QN(n4494) );
  DFFRX1 top_core_io_Data_reg_reg_35__6_ ( .D(top_core_io_n897), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_30_), .QN(n4493) );
  DFFRX1 top_core_io_Data_reg_reg_35__5_ ( .D(top_core_io_n896), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_29_), .QN(n4492) );
  DFFRX1 top_core_io_Data_reg_reg_35__4_ ( .D(top_core_io_n895), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_28_), .QN(n4491) );
  DFFRX1 top_core_io_Data_reg_reg_35__3_ ( .D(top_core_io_n894), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_27_), .QN(n4490) );
  DFFRX1 top_core_io_Data_reg_reg_35__2_ ( .D(top_core_io_n893), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_26_), .QN(n4489) );
  DFFRX1 top_core_io_Data_reg_reg_35__1_ ( .D(top_core_io_n892), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_25_), .QN(n4488) );
  DFFRX1 top_core_io_Data_reg_reg_35__0_ ( .D(top_core_io_n891), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_24_), .QN(n4487) );
  DFFRX1 top_core_io_Data_reg_reg_39__7_ ( .D(top_core_io_n866), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_63_), .QN(n4462) );
  DFFRX1 top_core_io_Data_reg_reg_39__6_ ( .D(top_core_io_n865), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_62_), .QN(n4461) );
  DFFRX1 top_core_io_Data_reg_reg_39__5_ ( .D(top_core_io_n864), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_61_), .QN(n4460) );
  DFFRX1 top_core_io_Data_reg_reg_39__4_ ( .D(top_core_io_n863), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_60_), .QN(n4459) );
  DFFRX1 top_core_io_Data_reg_reg_39__3_ ( .D(top_core_io_n862), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_59_), .QN(n4458) );
  DFFRX1 top_core_io_Data_reg_reg_39__2_ ( .D(top_core_io_n861), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_58_), .QN(n4457) );
  DFFRX1 top_core_io_Data_reg_reg_39__1_ ( .D(top_core_io_n860), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_57_), .QN(n4456) );
  DFFRX1 top_core_io_Data_reg_reg_39__0_ ( .D(top_core_io_n859), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_56_), .QN(n4455) );
  DFFRX1 top_core_io_Data_reg_reg_33__7_ ( .D(top_core_io_n914), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_15_), .QN(n4510) );
  DFFRX1 top_core_io_Data_reg_reg_33__6_ ( .D(top_core_io_n913), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_14_), .QN(n4509) );
  DFFRX1 top_core_io_Data_reg_reg_33__5_ ( .D(top_core_io_n912), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_13_), .QN(n4508) );
  DFFRX1 top_core_io_Data_reg_reg_33__4_ ( .D(top_core_io_n911), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_12_), .QN(n4507) );
  DFFRX1 top_core_io_Data_reg_reg_33__3_ ( .D(top_core_io_n910), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_11_), .QN(n4506) );
  DFFRX1 top_core_io_Data_reg_reg_33__2_ ( .D(top_core_io_n909), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_10_), .QN(n4505) );
  DFFRX1 top_core_io_Data_reg_reg_33__1_ ( .D(top_core_io_n908), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_9_), .QN(n4504) );
  DFFRX1 top_core_io_Data_reg_reg_33__0_ ( .D(top_core_io_n907), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_8_), .QN(n4503) );
  DFFRX1 top_core_io_Data_reg_reg_1__7_ ( .D(top_core_io_n1170), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_15_), .QN(n4766) );
  DFFRX1 top_core_io_Data_reg_reg_1__6_ ( .D(top_core_io_n1169), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_14_), .QN(n4765) );
  DFFRX1 top_core_io_Data_reg_reg_1__5_ ( .D(top_core_io_n1168), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_13_), .QN(n4764) );
  DFFRX1 top_core_io_Data_reg_reg_1__4_ ( .D(top_core_io_n1167), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_12_), .QN(n4763) );
  DFFRX1 top_core_io_Data_reg_reg_1__3_ ( .D(top_core_io_n1166), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_11_), .QN(n4762) );
  DFFRX1 top_core_io_Data_reg_reg_1__2_ ( .D(top_core_io_n1165), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_10_), .QN(n4761) );
  DFFRX1 top_core_io_Data_reg_reg_1__1_ ( .D(top_core_io_n1164), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_9_), .QN(n4760) );
  DFFRX1 top_core_io_Data_reg_reg_1__0_ ( .D(top_core_io_n1163), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_8_), .QN(n4759) );
  DFFRX1 top_core_io_Data_reg_reg_37__7_ ( .D(top_core_io_n882), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_47_), .QN(n4478) );
  DFFRX1 top_core_io_Data_reg_reg_37__6_ ( .D(top_core_io_n881), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_46_), .QN(n4477) );
  DFFRX1 top_core_io_Data_reg_reg_37__5_ ( .D(top_core_io_n880), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_45_), .QN(n4476) );
  DFFRX1 top_core_io_Data_reg_reg_37__4_ ( .D(top_core_io_n879), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_44_), .QN(n4475) );
  DFFRX1 top_core_io_Data_reg_reg_37__3_ ( .D(top_core_io_n878), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_43_), .QN(n4474) );
  DFFRX1 top_core_io_Data_reg_reg_37__2_ ( .D(top_core_io_n877), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_42_), .QN(n4473) );
  DFFRX1 top_core_io_Data_reg_reg_37__1_ ( .D(top_core_io_n876), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_41_), .QN(n4472) );
  DFFRX1 top_core_io_Data_reg_reg_37__0_ ( .D(top_core_io_n875), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_40_), .QN(n4471) );
  DFFRX1 top_core_io_Data_reg_reg_5__7_ ( .D(top_core_io_n1138), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_47_), .QN(n4734) );
  DFFRX1 top_core_io_Data_reg_reg_5__6_ ( .D(top_core_io_n1137), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_46_), .QN(n4733) );
  DFFRX1 top_core_io_Data_reg_reg_5__5_ ( .D(top_core_io_n1136), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_45_), .QN(n4732) );
  DFFRX1 top_core_io_Data_reg_reg_5__4_ ( .D(top_core_io_n1135), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_44_), .QN(n4731) );
  DFFRX1 top_core_io_Data_reg_reg_5__3_ ( .D(top_core_io_n1134), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_43_), .QN(n4730) );
  DFFRX1 top_core_io_Data_reg_reg_5__2_ ( .D(top_core_io_n1133), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_42_), .QN(n4729) );
  DFFRX1 top_core_io_Data_reg_reg_5__1_ ( .D(top_core_io_n1132), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_41_), .QN(n4728) );
  DFFRX1 top_core_io_Data_reg_reg_5__0_ ( .D(top_core_io_n1131), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_40_), .QN(n4727) );
  DFFRX1 top_core_io_Data_reg_reg_50__7_ ( .D(top_core_io_n778), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_151_), .QN(n4374) );
  DFFRX1 top_core_io_Data_reg_reg_50__6_ ( .D(top_core_io_n777), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_150_), .QN(n4373) );
  DFFRX1 top_core_io_Data_reg_reg_50__5_ ( .D(top_core_io_n776), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_149_), .QN(n4372) );
  DFFRX1 top_core_io_Data_reg_reg_50__4_ ( .D(top_core_io_n775), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_148_), .QN(n4371) );
  DFFRX1 top_core_io_Data_reg_reg_50__3_ ( .D(top_core_io_n774), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_147_), .QN(n4370) );
  DFFRX1 top_core_io_Data_reg_reg_50__2_ ( .D(top_core_io_n773), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_146_), .QN(n4369) );
  DFFRX1 top_core_io_Data_reg_reg_50__1_ ( .D(top_core_io_n772), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_145_), .QN(n4368) );
  DFFRX1 top_core_io_Data_reg_reg_50__0_ ( .D(top_core_io_n771), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_144_), .QN(n4367) );
  DFFRX1 top_core_io_Data_reg_reg_2__7_ ( .D(top_core_io_n1162), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_23_), .QN(n4758) );
  DFFRX1 top_core_io_Data_reg_reg_2__6_ ( .D(top_core_io_n1161), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_22_), .QN(n4757) );
  DFFRX1 top_core_io_Data_reg_reg_2__5_ ( .D(top_core_io_n1160), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_21_), .QN(n4756) );
  DFFRX1 top_core_io_Data_reg_reg_2__4_ ( .D(top_core_io_n1159), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_20_), .QN(n4755) );
  DFFRX1 top_core_io_Data_reg_reg_2__3_ ( .D(top_core_io_n1158), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_19_), .QN(n4754) );
  DFFRX1 top_core_io_Data_reg_reg_2__2_ ( .D(top_core_io_n1157), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_18_), .QN(n4753) );
  DFFRX1 top_core_io_Data_reg_reg_2__1_ ( .D(top_core_io_n1156), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_17_), .QN(n4752) );
  DFFRX1 top_core_io_Data_reg_reg_2__0_ ( .D(top_core_io_n1155), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_16_), .QN(n4751) );
  DFFRX1 top_core_io_Data_reg_reg_34__7_ ( .D(top_core_io_n906), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_23_), .QN(n4502) );
  DFFRX1 top_core_io_Data_reg_reg_34__6_ ( .D(top_core_io_n905), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_22_), .QN(n4501) );
  DFFRX1 top_core_io_Data_reg_reg_34__5_ ( .D(top_core_io_n904), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_21_), .QN(n4500) );
  DFFRX1 top_core_io_Data_reg_reg_34__4_ ( .D(top_core_io_n903), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_20_), .QN(n4499) );
  DFFRX1 top_core_io_Data_reg_reg_34__3_ ( .D(top_core_io_n902), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_19_), .QN(n4498) );
  DFFRX1 top_core_io_Data_reg_reg_34__2_ ( .D(top_core_io_n901), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_18_), .QN(n4497) );
  DFFRX1 top_core_io_Data_reg_reg_34__1_ ( .D(top_core_io_n900), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_17_), .QN(n4496) );
  DFFRX1 top_core_io_Data_reg_reg_34__0_ ( .D(top_core_io_n899), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_16_), .QN(n4495) );
  DFFRX1 top_core_io_Data_reg_reg_54__7_ ( .D(top_core_io_n746), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_183_), .QN(n4342) );
  DFFRX1 top_core_io_Data_reg_reg_54__6_ ( .D(top_core_io_n745), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_182_), .QN(n4341) );
  DFFRX1 top_core_io_Data_reg_reg_54__5_ ( .D(top_core_io_n744), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_181_), .QN(n4340) );
  DFFRX1 top_core_io_Data_reg_reg_54__4_ ( .D(top_core_io_n743), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_180_), .QN(n4339) );
  DFFRX1 top_core_io_Data_reg_reg_54__3_ ( .D(top_core_io_n742), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_179_), .QN(n4338) );
  DFFRX1 top_core_io_Data_reg_reg_54__2_ ( .D(top_core_io_n741), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_178_), .QN(n4337) );
  DFFRX1 top_core_io_Data_reg_reg_54__1_ ( .D(top_core_io_n740), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_177_), .QN(n4336) );
  DFFRX1 top_core_io_Data_reg_reg_54__0_ ( .D(top_core_io_n739), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_176_), .QN(n4335) );
  DFFRX1 top_core_io_Data_reg_reg_6__7_ ( .D(top_core_io_n1130), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_55_), .QN(n4726) );
  DFFRX1 top_core_io_Data_reg_reg_6__6_ ( .D(top_core_io_n1129), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_54_), .QN(n4725) );
  DFFRX1 top_core_io_Data_reg_reg_6__5_ ( .D(top_core_io_n1128), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_53_), .QN(n4724) );
  DFFRX1 top_core_io_Data_reg_reg_6__4_ ( .D(top_core_io_n1127), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_52_), .QN(n4723) );
  DFFRX1 top_core_io_Data_reg_reg_6__3_ ( .D(top_core_io_n1126), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_51_), .QN(n4722) );
  DFFRX1 top_core_io_Data_reg_reg_6__2_ ( .D(top_core_io_n1125), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_50_), .QN(n4721) );
  DFFRX1 top_core_io_Data_reg_reg_6__1_ ( .D(top_core_io_n1124), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_49_), .QN(n4720) );
  DFFRX1 top_core_io_Data_reg_reg_6__0_ ( .D(top_core_io_n1123), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_48_), .QN(n4719) );
  DFFRX1 top_core_io_Data_reg_reg_38__7_ ( .D(top_core_io_n874), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_55_), .QN(n4470) );
  DFFRX1 top_core_io_Data_reg_reg_38__6_ ( .D(top_core_io_n873), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_54_), .QN(n4469) );
  DFFRX1 top_core_io_Data_reg_reg_38__5_ ( .D(top_core_io_n872), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_53_), .QN(n4468) );
  DFFRX1 top_core_io_Data_reg_reg_38__4_ ( .D(top_core_io_n871), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_52_), .QN(n4467) );
  DFFRX1 top_core_io_Data_reg_reg_38__3_ ( .D(top_core_io_n870), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_51_), .QN(n4466) );
  DFFRX1 top_core_io_Data_reg_reg_38__2_ ( .D(top_core_io_n869), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_50_), .QN(n4465) );
  DFFRX1 top_core_io_Data_reg_reg_38__1_ ( .D(top_core_io_n868), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_49_), .QN(n4464) );
  DFFRX1 top_core_io_Data_reg_reg_38__0_ ( .D(top_core_io_n867), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_48_), .QN(n4463) );
  DFFRX1 top_core_io_Data_reg_reg_49__7_ ( .D(top_core_io_n786), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_143_), .QN(n4382) );
  DFFRX1 top_core_io_Data_reg_reg_49__6_ ( .D(top_core_io_n785), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_142_), .QN(n4381) );
  DFFRX1 top_core_io_Data_reg_reg_49__5_ ( .D(top_core_io_n784), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_141_), .QN(n4380) );
  DFFRX1 top_core_io_Data_reg_reg_49__4_ ( .D(top_core_io_n783), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_140_), .QN(n4379) );
  DFFRX1 top_core_io_Data_reg_reg_49__3_ ( .D(top_core_io_n782), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_139_), .QN(n4378) );
  DFFRX1 top_core_io_Data_reg_reg_49__2_ ( .D(top_core_io_n781), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_138_), .QN(n4377) );
  DFFRX1 top_core_io_Data_reg_reg_49__1_ ( .D(top_core_io_n780), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_137_), .QN(n4376) );
  DFFRX1 top_core_io_Data_reg_reg_49__0_ ( .D(top_core_io_n779), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_136_), .QN(n4375) );
  DFFRX1 top_core_io_Data_reg_reg_53__7_ ( .D(top_core_io_n754), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_175_), .QN(n4350) );
  DFFRX1 top_core_io_Data_reg_reg_53__6_ ( .D(top_core_io_n753), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_174_), .QN(n4349) );
  DFFRX1 top_core_io_Data_reg_reg_53__5_ ( .D(top_core_io_n752), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_173_), .QN(n4348) );
  DFFRX1 top_core_io_Data_reg_reg_53__4_ ( .D(top_core_io_n751), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_172_), .QN(n4347) );
  DFFRX1 top_core_io_Data_reg_reg_53__3_ ( .D(top_core_io_n750), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_171_), .QN(n4346) );
  DFFRX1 top_core_io_Data_reg_reg_53__2_ ( .D(top_core_io_n749), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_170_), .QN(n4345) );
  DFFRX1 top_core_io_Data_reg_reg_53__1_ ( .D(top_core_io_n748), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_169_), .QN(n4344) );
  DFFRX1 top_core_io_Data_reg_reg_53__0_ ( .D(top_core_io_n747), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_168_), .QN(n4343) );
  DFFRX1 top_core_io_Data_reg_reg_32__7_ ( .D(top_core_io_n922), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_7_), .QN(n4518) );
  DFFRX1 top_core_io_Data_reg_reg_32__6_ ( .D(top_core_io_n921), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_6_), .QN(n4517) );
  DFFRX1 top_core_io_Data_reg_reg_32__5_ ( .D(top_core_io_n920), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_5_), .QN(n4516) );
  DFFRX1 top_core_io_Data_reg_reg_32__4_ ( .D(top_core_io_n919), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_4_), .QN(n4515) );
  DFFRX1 top_core_io_Data_reg_reg_32__3_ ( .D(top_core_io_n918), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_3_), .QN(n4514) );
  DFFRX1 top_core_io_Data_reg_reg_32__2_ ( .D(top_core_io_n917), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_2_), .QN(n4513) );
  DFFRX1 top_core_io_Data_reg_reg_32__1_ ( .D(top_core_io_n916), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_1_), .QN(n4512) );
  DFFRX1 top_core_io_Data_reg_reg_32__0_ ( .D(top_core_io_n915), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_0_), .QN(n4511) );
  DFFRX1 top_core_io_Data_reg_reg_0__7_ ( .D(top_core_io_n1178), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_7_), .QN(n4774) );
  DFFRX1 top_core_io_Data_reg_reg_0__6_ ( .D(top_core_io_n1177), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_6_), .QN(n4773) );
  DFFRX1 top_core_io_Data_reg_reg_0__5_ ( .D(top_core_io_n1176), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_5_), .QN(n4772) );
  DFFRX1 top_core_io_Data_reg_reg_0__4_ ( .D(top_core_io_n1175), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_4_), .QN(n4771) );
  DFFRX1 top_core_io_Data_reg_reg_0__3_ ( .D(top_core_io_n1174), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_3_), .QN(n4770) );
  DFFRX1 top_core_io_Data_reg_reg_0__2_ ( .D(top_core_io_n1173), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_2_), .QN(n4769) );
  DFFRX1 top_core_io_Data_reg_reg_0__1_ ( .D(top_core_io_n1172), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_1_), .QN(n4768) );
  DFFRX1 top_core_io_Data_reg_reg_0__0_ ( .D(top_core_io_n1171), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_0_), .QN(n4767) );
  DFFRX1 top_core_io_Data_reg_reg_48__7_ ( .D(top_core_io_n794), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_135_), .QN(n4390) );
  DFFRX1 top_core_io_Data_reg_reg_48__6_ ( .D(top_core_io_n793), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_134_), .QN(n4389) );
  DFFRX1 top_core_io_Data_reg_reg_48__5_ ( .D(top_core_io_n792), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_133_), .QN(n4388) );
  DFFRX1 top_core_io_Data_reg_reg_48__4_ ( .D(top_core_io_n791), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_132_), .QN(n4387) );
  DFFRX1 top_core_io_Data_reg_reg_48__3_ ( .D(top_core_io_n790), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_131_), .QN(n4386) );
  DFFRX1 top_core_io_Data_reg_reg_48__2_ ( .D(top_core_io_n789), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_130_), .QN(n4385) );
  DFFRX1 top_core_io_Data_reg_reg_48__1_ ( .D(top_core_io_n788), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_129_), .QN(n4384) );
  DFFRX1 top_core_io_Data_reg_reg_48__0_ ( .D(top_core_io_n787), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_128_), .QN(n4383) );
  DFFRX1 top_core_io_Data_reg_reg_36__7_ ( .D(top_core_io_n890), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_39_), .QN(n4486) );
  DFFRX1 top_core_io_Data_reg_reg_36__6_ ( .D(top_core_io_n889), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_38_), .QN(n4485) );
  DFFRX1 top_core_io_Data_reg_reg_36__5_ ( .D(top_core_io_n888), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_37_), .QN(n4484) );
  DFFRX1 top_core_io_Data_reg_reg_36__4_ ( .D(top_core_io_n887), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_36_), .QN(n4483) );
  DFFRX1 top_core_io_Data_reg_reg_36__3_ ( .D(top_core_io_n886), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_35_), .QN(n4482) );
  DFFRX1 top_core_io_Data_reg_reg_36__2_ ( .D(top_core_io_n885), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_34_), .QN(n4481) );
  DFFRX1 top_core_io_Data_reg_reg_36__1_ ( .D(top_core_io_n884), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_33_), .QN(n4480) );
  DFFRX1 top_core_io_Data_reg_reg_36__0_ ( .D(top_core_io_n883), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_32_), .QN(n4479) );
  DFFRX1 top_core_io_Data_reg_reg_4__7_ ( .D(top_core_io_n1146), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_39_), .QN(n4742) );
  DFFRX1 top_core_io_Data_reg_reg_4__6_ ( .D(top_core_io_n1145), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_38_), .QN(n4741) );
  DFFRX1 top_core_io_Data_reg_reg_4__5_ ( .D(top_core_io_n1144), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_37_), .QN(n4740) );
  DFFRX1 top_core_io_Data_reg_reg_4__4_ ( .D(top_core_io_n1143), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_36_), .QN(n4739) );
  DFFRX1 top_core_io_Data_reg_reg_4__3_ ( .D(top_core_io_n1142), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_35_), .QN(n4738) );
  DFFRX1 top_core_io_Data_reg_reg_4__2_ ( .D(top_core_io_n1141), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_34_), .QN(n4737) );
  DFFRX1 top_core_io_Data_reg_reg_4__1_ ( .D(top_core_io_n1140), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_33_), .QN(n4736) );
  DFFRX1 top_core_io_Data_reg_reg_4__0_ ( .D(top_core_io_n1139), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_32_), .QN(n4735) );
  DFFRX1 top_core_io_Data_reg_reg_40__7_ ( .D(top_core_io_n858), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_71_), .QN(n4454) );
  DFFRX1 top_core_io_Data_reg_reg_40__6_ ( .D(top_core_io_n857), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_70_), .QN(n4453) );
  DFFRX1 top_core_io_Data_reg_reg_40__5_ ( .D(top_core_io_n856), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_69_), .QN(n4452) );
  DFFRX1 top_core_io_Data_reg_reg_40__4_ ( .D(top_core_io_n855), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_68_), .QN(n4451) );
  DFFRX1 top_core_io_Data_reg_reg_40__3_ ( .D(top_core_io_n854), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_67_), .QN(n4450) );
  DFFRX1 top_core_io_Data_reg_reg_40__2_ ( .D(top_core_io_n853), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_66_), .QN(n4449) );
  DFFRX1 top_core_io_Data_reg_reg_40__1_ ( .D(top_core_io_n852), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_65_), .QN(n4448) );
  DFFRX1 top_core_io_Data_reg_reg_40__0_ ( .D(top_core_io_n851), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_64_), .QN(n4447) );
  DFFRX1 top_core_io_Data_reg_reg_8__7_ ( .D(top_core_io_n1114), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_71_), .QN(n4710) );
  DFFRX1 top_core_io_Data_reg_reg_8__6_ ( .D(top_core_io_n1113), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_70_), .QN(n4709) );
  DFFRX1 top_core_io_Data_reg_reg_8__5_ ( .D(top_core_io_n1112), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_69_), .QN(n4708) );
  DFFRX1 top_core_io_Data_reg_reg_8__4_ ( .D(top_core_io_n1111), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_68_), .QN(n4707) );
  DFFRX1 top_core_io_Data_reg_reg_8__3_ ( .D(top_core_io_n1110), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_67_), .QN(n4706) );
  DFFRX1 top_core_io_Data_reg_reg_8__2_ ( .D(top_core_io_n1109), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_66_), .QN(n4705) );
  DFFRX1 top_core_io_Data_reg_reg_8__1_ ( .D(top_core_io_n1108), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_65_), .QN(n4704) );
  DFFRX1 top_core_io_Data_reg_reg_8__0_ ( .D(top_core_io_n1107), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_Plain_text_w_64_), .QN(n4703) );
  DFFRX1 top_core_io_Data_reg_reg_52__7_ ( .D(top_core_io_n762), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_167_), .QN(n4358) );
  DFFRX1 top_core_io_Data_reg_reg_52__6_ ( .D(top_core_io_n761), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_166_), .QN(n4357) );
  DFFRX1 top_core_io_Data_reg_reg_52__5_ ( .D(top_core_io_n760), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_165_), .QN(n4356) );
  DFFRX1 top_core_io_Data_reg_reg_52__4_ ( .D(top_core_io_n759), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_164_), .QN(n4355) );
  DFFRX1 top_core_io_Data_reg_reg_52__3_ ( .D(top_core_io_n758), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_163_), .QN(n4354) );
  DFFRX1 top_core_io_Data_reg_reg_52__2_ ( .D(top_core_io_n757), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_162_), .QN(n4353) );
  DFFRX1 top_core_io_Data_reg_reg_52__1_ ( .D(top_core_io_n756), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_161_), .QN(n4352) );
  DFFRX1 top_core_io_Data_reg_reg_52__0_ ( .D(top_core_io_n755), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_160_), .QN(n4351) );
  DFFRX1 top_core_io_Data_reg_reg_56__7_ ( .D(top_core_io_n730), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_199_), .QN(n4326) );
  DFFRX1 top_core_io_Data_reg_reg_56__6_ ( .D(top_core_io_n729), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_198_), .QN(n4325) );
  DFFRX1 top_core_io_Data_reg_reg_56__5_ ( .D(top_core_io_n728), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_197_), .QN(n4324) );
  DFFRX1 top_core_io_Data_reg_reg_56__4_ ( .D(top_core_io_n727), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_196_), .QN(n4323) );
  DFFRX1 top_core_io_Data_reg_reg_56__3_ ( .D(top_core_io_n726), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_195_), .QN(n4322) );
  DFFRX1 top_core_io_Data_reg_reg_56__2_ ( .D(top_core_io_n725), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_194_), .QN(n4321) );
  DFFRX1 top_core_io_Data_reg_reg_56__1_ ( .D(top_core_io_n724), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_193_), .QN(n4320) );
  DFFRX1 top_core_io_Data_reg_reg_56__0_ ( .D(top_core_io_n723), .CK(n_CLK), 
        .RN(n_RSTB), .Q(top_core_io_CipherKey_w_192_), .QN(n4319) );
  OAI221XL U4 ( .A0(n13985), .A1(n13857), .B0(n3494), .B1(n107), .C0(n13980), 
        .Y(n14148) );
  CLKINVX3 U5 ( .A(n3497), .Y(n3493) );
  AOI221X1 U6 ( .A0(n6137), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .B0(
        n6165), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n328), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n327) );
  OAI221XL U7 ( .A0(n385), .A1(n58), .B0(n13925), .B1(n13867), .C0(n14099), 
        .Y(n14098) );
  OAI221XL U8 ( .A0(n497), .A1(n107), .B0(n13925), .B1(n3501), .C0(n14105), 
        .Y(n14100) );
  OAI221XL U9 ( .A0(n13857), .A1(n13864), .B0(n3483), .B1(n165), .C0(n14070), 
        .Y(n14068) );
  OAI222XL U10 ( .A0(n91), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .B0(
        n3483), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n101), .C0(n1145), .C1(
        n1140), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n291) );
  AOI221X1 U11 ( .A0(n1139), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), 
        .B0(n1145), .B1(n545), .C0(top_core_EC_ss_gen_tbox_0__sboxs_r_n75), 
        .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n284) );
  AOI211X1 U12 ( .A0(n14033), .A1(n3483), .B0(n14042), .C0(n258), .Y(n14041)
         );
  OAI221XL U13 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n71), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .B0(n3491), .B1(n91), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n207), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n219) );
  OAI221XL U14 ( .A0(n15560), .A1(n15432), .B0(n3192), .B1(n110), .C0(n15555), 
        .Y(n15723) );
  CLKINVX3 U15 ( .A(n3195), .Y(n3191) );
  AOI221X1 U16 ( .A0(n5071), .A1(n10776), .B0(n5105), .B1(n10789), .C0(n11018), 
        .Y(n11017) );
  OAI221XL U17 ( .A0(n389), .A1(n61), .B0(n15500), .B1(n15442), .C0(n15674), 
        .Y(n15673) );
  OAI221XL U18 ( .A0(n499), .A1(n110), .B0(n15500), .B1(n3199), .C0(n15680), 
        .Y(n15675) );
  OAI221XL U19 ( .A0(n15432), .A1(n15439), .B0(n3181), .B1(n168), .C0(n15645), 
        .Y(n15643) );
  OAI222XL U20 ( .A0(n94), .A1(n10776), .B0(n2701), .B1(n10793), .C0(n962), 
        .C1(n958), .Y(n10981) );
  AOI221X1 U21 ( .A0(n954), .A1(n10846), .B0(n962), .B1(n549), .C0(n10768), 
        .Y(n10974) );
  AOI211X1 U22 ( .A0(n15608), .A1(n3181), .B0(n15617), .C0(n255), .Y(n15616)
         );
  OAI221XL U23 ( .A0(n10765), .A1(n10776), .B0(n2706), .B1(n94), .C0(n10897), 
        .Y(n10909) );
  OAI221XL U24 ( .A0(n17135), .A1(n17007), .B0(n2893), .B1(n106), .C0(n17130), 
        .Y(n17298) );
  CLKINVX3 U25 ( .A(n2896), .Y(n2892) );
  AOI221X1 U26 ( .A0(n5341), .A1(n9900), .B0(n5375), .B1(n9913), .C0(n10142), 
        .Y(n10141) );
  OAI221XL U27 ( .A0(n386), .A1(n57), .B0(n17075), .B1(n17017), .C0(n17249), 
        .Y(n17248) );
  OAI221XL U28 ( .A0(n498), .A1(n106), .B0(n17075), .B1(n2900), .C0(n17255), 
        .Y(n17250) );
  OAI221XL U29 ( .A0(n17007), .A1(n17014), .B0(n2882), .B1(n164), .C0(n17220), 
        .Y(n17218) );
  OAI222XL U30 ( .A0(n90), .A1(n9900), .B0(n2882), .B1(n9917), .C0(n1004), 
        .C1(n1000), .Y(n10105) );
  AOI221X1 U31 ( .A0(n996), .A1(n9970), .B0(n1004), .B1(n546), .C0(n9892), .Y(
        n10098) );
  AOI211X1 U32 ( .A0(n17183), .A1(n2882), .B0(n17192), .C0(n259), .Y(n17191)
         );
  OAI221XL U33 ( .A0(n9889), .A1(n9900), .B0(n2887), .B1(n90), .C0(n10021), 
        .Y(n10033) );
  OAI221XL U34 ( .A0(n18710), .A1(n18582), .B0(n2590), .B1(n111), .C0(n18705), 
        .Y(n18873) );
  CLKINVX3 U35 ( .A(n2592), .Y(n2589) );
  AOI221X1 U36 ( .A0(n5577), .A1(n9024), .B0(n5611), .B1(n9037), .C0(n9266), 
        .Y(n9265) );
  OAI221XL U37 ( .A0(n390), .A1(n63), .B0(n18650), .B1(n18592), .C0(n18824), 
        .Y(n18823) );
  OAI221XL U38 ( .A0(n502), .A1(n111), .B0(n18650), .B1(n2596), .C0(n18830), 
        .Y(n18825) );
  OAI221XL U39 ( .A0(n18582), .A1(n18589), .B0(n2579), .B1(n169), .C0(n18795), 
        .Y(n18793) );
  OAI222XL U40 ( .A0(n96), .A1(n9024), .B0(n3062), .B1(n9041), .C0(n1046), 
        .C1(n1042), .Y(n9229) );
  AOI221X1 U41 ( .A0(n1038), .A1(n9094), .B0(n1046), .B1(n550), .C0(n9016), 
        .Y(n9222) );
  AOI211X1 U42 ( .A0(n18758), .A1(n2579), .B0(n18767), .C0(n253), .Y(n18766)
         );
  OAI221XL U43 ( .A0(n9013), .A1(n9024), .B0(n3066), .B1(n96), .C0(n9145), .Y(
        n9157) );
  OAI221XL U44 ( .A0(n15245), .A1(n15117), .B0(n3253), .B1(n109), .C0(n15240), 
        .Y(n15408) );
  CLKINVX3 U45 ( .A(n3256), .Y(n3252) );
  AOI221X1 U46 ( .A0(n5813), .A1(n8148), .B0(n5847), .B1(n8161), .C0(n8390), 
        .Y(n8389) );
  OAI221XL U47 ( .A0(n388), .A1(n60), .B0(n15185), .B1(n15127), .C0(n15359), 
        .Y(n15358) );
  OAI221XL U48 ( .A0(n500), .A1(n109), .B0(n15185), .B1(n3260), .C0(n15365), 
        .Y(n15360) );
  OAI221XL U49 ( .A0(n15117), .A1(n15124), .B0(n3242), .B1(n167), .C0(n15330), 
        .Y(n15328) );
  OAI222XL U50 ( .A0(n93), .A1(n8148), .B0(n3242), .B1(n8165), .C0(n1088), 
        .C1(n1084), .Y(n8353) );
  AOI221X1 U51 ( .A0(n1080), .A1(n8218), .B0(n1088), .B1(n548), .C0(n8140), 
        .Y(n8346) );
  AOI211X1 U52 ( .A0(n15293), .A1(n3242), .B0(n15302), .C0(n256), .Y(n15301)
         );
  OAI221XL U53 ( .A0(n8137), .A1(n8148), .B0(n3246), .B1(n93), .C0(n8269), .Y(
        n8281) );
  OAI221XL U54 ( .A0(n16820), .A1(n16692), .B0(n2954), .B1(n112), .C0(n16815), 
        .Y(n16983) );
  CLKINVX3 U55 ( .A(n2957), .Y(n2953) );
  AOI221X1 U56 ( .A0(n6041), .A1(n7272), .B0(n6075), .B1(n7285), .C0(n7514), 
        .Y(n7513) );
  OAI221XL U57 ( .A0(n391), .A1(n62), .B0(n16760), .B1(n16702), .C0(n16934), 
        .Y(n16933) );
  OAI221XL U58 ( .A0(n503), .A1(n112), .B0(n16760), .B1(n2961), .C0(n16940), 
        .Y(n16935) );
  OAI221XL U59 ( .A0(n16692), .A1(n16699), .B0(n2943), .B1(n170), .C0(n16905), 
        .Y(n16903) );
  OAI222XL U60 ( .A0(n95), .A1(n7272), .B0(n3422), .B1(n7289), .C0(n1130), 
        .C1(n1126), .Y(n7477) );
  AOI221X1 U61 ( .A0(n1122), .A1(n7342), .B0(n1130), .B1(n551), .C0(n7264), 
        .Y(n7470) );
  AOI211X1 U62 ( .A0(n16868), .A1(n2943), .B0(n16877), .C0(n254), .Y(n16876)
         );
  OAI221XL U63 ( .A0(n7261), .A1(n7272), .B0(n3426), .B1(n95), .C0(n7393), .Y(
        n7405) );
  OAI221XL U64 ( .A0(n18395), .A1(n18267), .B0(n2650), .B1(n108), .C0(n18390), 
        .Y(n18558) );
  AOI221X1 U65 ( .A0(n4987), .A1(n11068), .B0(n5021), .B1(n11081), .C0(n11310), 
        .Y(n11309) );
  OAI221XL U66 ( .A0(n387), .A1(n59), .B0(n18335), .B1(n18277), .C0(n18509), 
        .Y(n18508) );
  OAI221XL U67 ( .A0(n501), .A1(n108), .B0(n18335), .B1(n2657), .C0(n18515), 
        .Y(n18510) );
  OAI221XL U68 ( .A0(n18267), .A1(n18274), .B0(n2640), .B1(n166), .C0(n18480), 
        .Y(n18478) );
  OAI222XL U69 ( .A0(n92), .A1(n11068), .B0(n2640), .B1(n11085), .C0(n948), 
        .C1(n944), .Y(n11273) );
  AOI221X1 U70 ( .A0(n940), .A1(n11138), .B0(n948), .B1(n547), .C0(n11060), 
        .Y(n11266) );
  AOI211X1 U71 ( .A0(n18443), .A1(n2640), .B0(n18452), .C0(n257), .Y(n18451)
         );
  OAI221XL U72 ( .A0(n11057), .A1(n11068), .B0(n2644), .B1(n92), .C0(n11189), 
        .Y(n11201) );
  OAI221XL U73 ( .A0(n14930), .A1(n14802), .B0(n3314), .B1(n113), .C0(n14925), 
        .Y(n15093) );
  CLKINVX3 U74 ( .A(n3319), .Y(n3313) );
  AOI221X1 U75 ( .A0(n5257), .A1(n10192), .B0(n5291), .B1(n10205), .C0(n10434), 
        .Y(n10433) );
  OAI221XL U76 ( .A0(n392), .A1(n64), .B0(n14870), .B1(n14812), .C0(n15044), 
        .Y(n15043) );
  OAI221XL U77 ( .A0(n504), .A1(n113), .B0(n14870), .B1(n3323), .C0(n15050), 
        .Y(n15045) );
  OAI221XL U78 ( .A0(n14802), .A1(n14809), .B0(n3303), .B1(n171), .C0(n15015), 
        .Y(n15013) );
  OAI222XL U79 ( .A0(n97), .A1(n10192), .B0(n2822), .B1(n10209), .C0(n990), 
        .C1(n986), .Y(n10397) );
  AOI221X1 U80 ( .A0(n982), .A1(n10262), .B0(n990), .B1(n552), .C0(n10184), 
        .Y(n10390) );
  AOI211X1 U81 ( .A0(n14978), .A1(n3303), .B0(n14987), .C0(n252), .Y(n14986)
         );
  OAI221XL U82 ( .A0(n10181), .A1(n10192), .B0(n2826), .B1(n97), .C0(n10313), 
        .Y(n10325) );
  OAI221XL U83 ( .A0(n16505), .A1(n16377), .B0(n3015), .B1(n114), .C0(n16500), 
        .Y(n16668) );
  CLKINVX3 U84 ( .A(n3020), .Y(n3014) );
  AOI221X1 U85 ( .A0(n5501), .A1(n9316), .B0(n5535), .B1(n9329), .C0(n9558), 
        .Y(n9557) );
  OAI221XL U86 ( .A0(n393), .A1(n65), .B0(n16445), .B1(n16387), .C0(n16619), 
        .Y(n16618) );
  OAI221XL U87 ( .A0(n505), .A1(n114), .B0(n16445), .B1(n3024), .C0(n16625), 
        .Y(n16620) );
  OAI221XL U88 ( .A0(n16377), .A1(n16384), .B0(n3004), .B1(n172), .C0(n16590), 
        .Y(n16588) );
  OAI222XL U89 ( .A0(n98), .A1(n9316), .B0(n3004), .B1(n9333), .C0(n1032), 
        .C1(n1028), .Y(n9521) );
  AOI221X1 U90 ( .A0(n1024), .A1(n9386), .B0(n1032), .B1(n553), .C0(n9308), 
        .Y(n9514) );
  AOI211X1 U91 ( .A0(n16553), .A1(n3004), .B0(n16562), .C0(n251), .Y(n16561)
         );
  OAI221XL U92 ( .A0(n9305), .A1(n9316), .B0(n3008), .B1(n98), .C0(n9437), .Y(
        n9449) );
  OAI221XL U93 ( .A0(n18080), .A1(n17952), .B0(n2711), .B1(n115), .C0(n18075), 
        .Y(n18243) );
  CLKINVX3 U94 ( .A(n2714), .Y(n2710) );
  AOI221X1 U95 ( .A0(n5729), .A1(n8440), .B0(n5763), .B1(n8453), .C0(n8682), 
        .Y(n8681) );
  OAI221XL U96 ( .A0(n394), .A1(n66), .B0(n18020), .B1(n17962), .C0(n18194), 
        .Y(n18193) );
  OAI221XL U97 ( .A0(n506), .A1(n115), .B0(n18020), .B1(n2718), .C0(n18200), 
        .Y(n18195) );
  OAI221XL U98 ( .A0(n17952), .A1(n17959), .B0(n2701), .B1(n173), .C0(n18165), 
        .Y(n18163) );
  OAI222XL U99 ( .A0(n99), .A1(n8440), .B0(n3181), .B1(n8457), .C0(n1074), 
        .C1(n1070), .Y(n8645) );
  AOI221X1 U100 ( .A0(n1066), .A1(n8510), .B0(n1074), .B1(n554), .C0(n8432), 
        .Y(n8638) );
  AOI211X1 U101 ( .A0(n18128), .A1(n2701), .B0(n18137), .C0(n250), .Y(n18136)
         );
  OAI221XL U102 ( .A0(n8429), .A1(n8440), .B0(n3186), .B1(n99), .C0(n8561), 
        .Y(n8573) );
  OAI221XL U103 ( .A0(n14615), .A1(n14487), .B0(n3375), .B1(n116), .C0(n14610), 
        .Y(n14778) );
  CLKINVX3 U104 ( .A(n3380), .Y(n3374) );
  AOI221X1 U105 ( .A0(n5965), .A1(n7564), .B0(n5999), .B1(n7577), .C0(n7806), 
        .Y(n7805) );
  OAI221XL U106 ( .A0(n395), .A1(n67), .B0(n14555), .B1(n14497), .C0(n14729), 
        .Y(n14728) );
  OAI221XL U107 ( .A0(n507), .A1(n116), .B0(n14555), .B1(n3384), .C0(n14735), 
        .Y(n14730) );
  OAI221XL U108 ( .A0(n14487), .A1(n14494), .B0(n3364), .B1(n174), .C0(n14700), 
        .Y(n14698) );
  OAI222XL U109 ( .A0(n100), .A1(n7564), .B0(n3364), .B1(n7581), .C0(n1116), 
        .C1(n1112), .Y(n7769) );
  AOI221X1 U110 ( .A0(n1108), .A1(n7634), .B0(n1116), .B1(n555), .C0(n7556), 
        .Y(n7762) );
  AOI211X1 U111 ( .A0(n14663), .A1(n3364), .B0(n14672), .C0(n249), .Y(n14671)
         );
  OAI221XL U112 ( .A0(n7553), .A1(n7564), .B0(n3369), .B1(n100), .C0(n7685), 
        .Y(n7697) );
  OAI221XL U113 ( .A0(n16190), .A1(n16062), .B0(n3072), .B1(n117), .C0(n16185), 
        .Y(n16353) );
  AOI221X1 U114 ( .A0(n4871), .A1(n11360), .B0(n4905), .B1(n11373), .C0(n11602), .Y(n11601) );
  OAI221XL U115 ( .A0(n396), .A1(n68), .B0(n16130), .B1(n16072), .C0(n16304), 
        .Y(n16303) );
  OAI221XL U116 ( .A0(n508), .A1(n117), .B0(n16130), .B1(n3079), .C0(n16310), 
        .Y(n16305) );
  OAI221XL U117 ( .A0(n16062), .A1(n16069), .B0(n3062), .B1(n175), .C0(n16275), 
        .Y(n16273) );
  OAI222XL U118 ( .A0(n101), .A1(n11360), .B0(n2579), .B1(n11377), .C0(n934), 
        .C1(n930), .Y(n11565) );
  AOI221X1 U119 ( .A0(n926), .A1(n11430), .B0(n934), .B1(n556), .C0(n11352), 
        .Y(n11558) );
  AOI211X1 U120 ( .A0(n16238), .A1(n3062), .B0(n16247), .C0(n248), .Y(n16246)
         );
  OAI221XL U121 ( .A0(n11349), .A1(n11360), .B0(n2584), .B1(n101), .C0(n11481), 
        .Y(n11493) );
  OAI221XL U122 ( .A0(n17765), .A1(n17637), .B0(n2772), .B1(n118), .C0(n17760), 
        .Y(n17928) );
  CLKINVX3 U123 ( .A(n2779), .Y(n2771) );
  AOI221X1 U124 ( .A0(n5179), .A1(n10484), .B0(n5213), .B1(n10497), .C0(n10726), .Y(n10725) );
  OAI221XL U125 ( .A0(n397), .A1(n69), .B0(n17705), .B1(n17647), .C0(n17879), 
        .Y(n17878) );
  OAI221XL U126 ( .A0(n509), .A1(n118), .B0(n17705), .B1(n2781), .C0(n17885), 
        .Y(n17880) );
  OAI221XL U127 ( .A0(n17637), .A1(n17644), .B0(n2761), .B1(n176), .C0(n17850), 
        .Y(n17848) );
  OAI222XL U128 ( .A0(n102), .A1(n10484), .B0(n2761), .B1(n10501), .C0(n976), 
        .C1(n972), .Y(n10689) );
  AOI221X1 U129 ( .A0(n968), .A1(n10554), .B0(n976), .B1(n557), .C0(n10476), 
        .Y(n10682) );
  AOI211X1 U130 ( .A0(n17813), .A1(n2761), .B0(n17822), .C0(n247), .Y(n17821)
         );
  OAI221XL U131 ( .A0(n10473), .A1(n10484), .B0(n2766), .B1(n102), .C0(n10605), 
        .Y(n10617) );
  OAI221XL U132 ( .A0(n14300), .A1(n14172), .B0(n3433), .B1(n119), .C0(n14295), 
        .Y(n14463) );
  CLKINVX3 U133 ( .A(n3436), .Y(n3432) );
  AOI221X1 U134 ( .A0(n5425), .A1(n9608), .B0(n5459), .B1(n9621), .C0(n9850), 
        .Y(n9849) );
  OAI221XL U135 ( .A0(n398), .A1(n70), .B0(n14240), .B1(n14182), .C0(n14414), 
        .Y(n14413) );
  OAI221XL U136 ( .A0(n510), .A1(n119), .B0(n14240), .B1(n3440), .C0(n14420), 
        .Y(n14415) );
  OAI221XL U137 ( .A0(n14172), .A1(n14179), .B0(n3422), .B1(n177), .C0(n14385), 
        .Y(n14383) );
  OAI222XL U138 ( .A0(n103), .A1(n9608), .B0(n2943), .B1(n9625), .C0(n1018), 
        .C1(n1014), .Y(n9813) );
  AOI221X1 U139 ( .A0(n1010), .A1(n9678), .B0(n1018), .B1(n558), .C0(n9600), 
        .Y(n9806) );
  AOI211X1 U140 ( .A0(n14348), .A1(n3422), .B0(n14357), .C0(n246), .Y(n14356)
         );
  OAI221XL U141 ( .A0(n9597), .A1(n9608), .B0(n2948), .B1(n103), .C0(n9729), 
        .Y(n9741) );
  OAI221XL U142 ( .A0(n15875), .A1(n15747), .B0(n3134), .B1(n120), .C0(n15870), 
        .Y(n16038) );
  CLKINVX3 U143 ( .A(n3139), .Y(n3133) );
  AOI221X1 U144 ( .A0(n5653), .A1(n8732), .B0(n5687), .B1(n8745), .C0(n8974), 
        .Y(n8973) );
  OAI221XL U145 ( .A0(n399), .A1(n71), .B0(n15815), .B1(n15757), .C0(n15989), 
        .Y(n15988) );
  OAI221XL U146 ( .A0(n511), .A1(n120), .B0(n15815), .B1(n3143), .C0(n15995), 
        .Y(n15990) );
  OAI221XL U147 ( .A0(n15747), .A1(n15754), .B0(n3123), .B1(n178), .C0(n15960), 
        .Y(n15958) );
  OAI222XL U148 ( .A0(n104), .A1(n8732), .B0(n3123), .B1(n8749), .C0(n1060), 
        .C1(n1056), .Y(n8937) );
  AOI221X1 U149 ( .A0(n1052), .A1(n8802), .B0(n1060), .B1(n559), .C0(n8724), 
        .Y(n8930) );
  AOI211X1 U150 ( .A0(n15923), .A1(n3123), .B0(n15932), .C0(n245), .Y(n15931)
         );
  OAI221XL U151 ( .A0(n8721), .A1(n8732), .B0(n3128), .B1(n104), .C0(n8853), 
        .Y(n8865) );
  OAI221XL U152 ( .A0(n17450), .A1(n17322), .B0(n2833), .B1(n121), .C0(n17445), 
        .Y(n17613) );
  CLKINVX3 U153 ( .A(n2839), .Y(n2832) );
  AOI221X1 U154 ( .A0(n5889), .A1(n7856), .B0(n5923), .B1(n7869), .C0(n8098), 
        .Y(n8097) );
  OAI221XL U155 ( .A0(n400), .A1(n72), .B0(n17390), .B1(n17332), .C0(n17564), 
        .Y(n17563) );
  OAI221XL U156 ( .A0(n512), .A1(n121), .B0(n17390), .B1(n2843), .C0(n17570), 
        .Y(n17565) );
  OAI221XL U157 ( .A0(n17322), .A1(n17329), .B0(n2822), .B1(n179), .C0(n17535), 
        .Y(n17533) );
  OAI222XL U158 ( .A0(n105), .A1(n7856), .B0(n3303), .B1(n7873), .C0(n1102), 
        .C1(n1098), .Y(n8061) );
  AOI221X1 U159 ( .A0(n1094), .A1(n7926), .B0(n1102), .B1(n560), .C0(n7848), 
        .Y(n8054) );
  AOI211X1 U160 ( .A0(n17498), .A1(n2822), .B0(n17507), .C0(n244), .Y(n17506)
         );
  OAI221XL U161 ( .A0(n7845), .A1(n7856), .B0(n3307), .B1(n105), .C0(n7977), 
        .Y(n7989) );
  OAI22X2 U162 ( .A0(n2396), .A1(top_core_EC_ss_n146), .B0(n2374), .B1(n125), 
        .Y(top_core_EC_mc_mix_in_8[80]) );
  OAI22X2 U163 ( .A0(n2396), .A1(top_core_EC_ss_n145), .B0(n2374), .B1(n124), 
        .Y(top_core_EC_mc_mix_in_4_80_) );
  OAI22X2 U164 ( .A0(n2401), .A1(top_core_EC_ss_n144), .B0(n2374), .B1(n123), 
        .Y(top_core_EC_mc_mix_in_2_80_) );
  OAI22X2 U165 ( .A0(n2439), .A1(top_core_EC_ss_n164), .B0(n2372), .B1(n127), 
        .Y(top_core_EC_mc_mix_in_8[64]) );
  OAI22X2 U166 ( .A0(n2439), .A1(top_core_EC_ss_n162), .B0(n2372), .B1(n126), 
        .Y(top_core_EC_mc_mix_in_4_64_) );
  OAI22X2 U167 ( .A0(n2428), .A1(top_core_EC_ss_n238), .B0(
        top_core_EC_operation), .B1(n132), .Y(top_core_EC_mc_mix_in_8[112]) );
  OAI22X2 U168 ( .A0(n2531), .A1(top_core_EC_ss_n237), .B0(n2536), .B1(n131), 
        .Y(top_core_EC_mc_mix_in_4_112_) );
  OAI22X2 U169 ( .A0(n2528), .A1(top_core_EC_ss_n236), .B0(n2539), .B1(n130), 
        .Y(top_core_EC_mc_mix_in_2_112_) );
  OAI22X2 U170 ( .A0(n2419), .A1(top_core_EC_ss_n255), .B0(n2367), .B1(n134), 
        .Y(top_core_EC_mc_mix_in_8[96]) );
  OAI22X2 U171 ( .A0(n2437), .A1(top_core_EC_ss_n254), .B0(n2367), .B1(n133), 
        .Y(top_core_EC_mc_mix_in_4_96_) );
  AOI211X1 U172 ( .A0(n12588), .A1(n12638), .B0(n12628), .C0(n6841), .Y(n12784) );
  AOI211X1 U173 ( .A0(n13218), .A1(n13268), .B0(n13258), .C0(n6546), .Y(n13414) );
  AOI211X1 U174 ( .A0(n12903), .A1(n12953), .B0(n12943), .C0(n6887), .Y(n13099) );
  OAI222XL U175 ( .A0(n191), .A1(n12908), .B0(n12978), .B1(n12923), .C0(n12979), .C1(n12980), .Y(n12975) );
  OAI222XL U176 ( .A0(n189), .A1(n12593), .B0(n12663), .B1(n12608), .C0(n12664), .C1(n12665), .Y(n12660) );
  AOI211X1 U177 ( .A0(n13533), .A1(n13583), .B0(n13573), .C0(n6594), .Y(n13729) );
  OAI222XL U178 ( .A0(n190), .A1(n13538), .B0(n13608), .B1(n13553), .C0(n13609), .C1(n13610), .Y(n13605) );
  OAI22X2 U179 ( .A0(n2420), .A1(top_core_EC_ss_n215), .B0(n2369), .B1(n5310), 
        .Y(top_core_EC_mc_mix_in_4_16_) );
  OAI22X2 U180 ( .A0(n2439), .A1(top_core_EC_ss_n163), .B0(n2372), .B1(n6093), 
        .Y(top_core_EC_mc_mix_in_4_0_) );
  OAI22X2 U181 ( .A0(n2493), .A1(top_core_EC_ss_n174), .B0(n2372), .B1(n6097), 
        .Y(top_core_EC_mc_mix_in_8[0]) );
  OAI22X2 U182 ( .A0(n2424), .A1(top_core_EC_ss_n216), .B0(n2369), .B1(n5311), 
        .Y(top_core_EC_mc_mix_in_8[16]) );
  OAI22X2 U183 ( .A0(n2395), .A1(top_core_EC_ss_n152), .B0(n2373), .B1(n6096), 
        .Y(top_core_EC_mc_mix_in_2_0_) );
  OAI22X2 U184 ( .A0(n2436), .A1(top_core_EC_ss_n179), .B0(n2371), .B1(n4950), 
        .Y(top_core_EC_mc_mix_in_2_48_) );
  OAI22X2 U185 ( .A0(n2436), .A1(top_core_EC_ss_n180), .B0(n2371), .B1(n4955), 
        .Y(top_core_EC_mc_mix_in_4_48_) );
  OAI22X2 U186 ( .A0(n2430), .A1(top_core_EC_ss_n198), .B0(n2370), .B1(n5782), 
        .Y(top_core_EC_mc_mix_in_4_32_) );
  OAI22X2 U187 ( .A0(n2436), .A1(top_core_EC_ss_n181), .B0(n2371), .B1(n4957), 
        .Y(top_core_EC_mc_mix_in_8[48]) );
  OAI22X2 U188 ( .A0(n2430), .A1(top_core_EC_ss_n199), .B0(n2370), .B1(n5783), 
        .Y(top_core_EC_mc_mix_in_8[32]) );
  OAI221XL U189 ( .A0(n1182), .A1(n12410), .B0(n12349), .B1(n1263), .C0(n12524), .Y(n12523) );
  OAI221XL U190 ( .A0(n11779), .A1(n11691), .B0(n11929), .B1(n185), .C0(n11673), .Y(n11933) );
  OAI221XL U191 ( .A0(top_core_KE_sb1_n207), .A1(top_core_KE_sb1_n116), .B0(
        top_core_KE_sb1_n358), .B1(n186), .C0(top_core_KE_sb1_n98), .Y(
        top_core_KE_sb1_n362) );
  OAI221XL U192 ( .A0(n1223), .A1(n11779), .B0(n11718), .B1(n11661), .C0(
        n11893), .Y(n11892) );
  OAI221XL U193 ( .A0(n1217), .A1(top_core_KE_sb1_n207), .B0(
        top_core_KE_sb1_n145), .B1(top_core_KE_sb1_n86), .C0(
        top_core_KE_sb1_n322), .Y(top_core_KE_sb1_n321) );
  OAI221XL U194 ( .A0(n12410), .A1(n12322), .B0(n12560), .B1(n46), .C0(n12304), 
        .Y(n12564) );
  OAI221XL U195 ( .A0(n12095), .A1(n12007), .B0(n12245), .B1(n188), .C0(n11989), .Y(n12249) );
  OAI221XL U196 ( .A0(n1177), .A1(n12095), .B0(n12034), .B1(n11977), .C0(
        n12209), .Y(n12208) );
  OAI222XL U197 ( .A0(top_core_KE_sb1_n145), .A1(top_core_KE_sb1_n130), .B0(
        n1824), .B1(top_core_KE_sb1_n143), .C0(n1352), .C1(
        top_core_KE_sb1_n162), .Y(top_core_KE_sb1_n158) );
  AOI222X1 U198 ( .A0(n6915), .A1(n11705), .B0(n6919), .B1(n1808), .C0(n6904), 
        .C1(n1257), .Y(n11871) );
  OAI221XL U199 ( .A0(n11651), .A1(n11658), .B0(n1803), .B1(n77), .C0(n11864), 
        .Y(n11862) );
  AOI222X1 U200 ( .A0(n6869), .A1(top_core_KE_sb1_n130), .B0(n6873), .B1(n1829), .C0(n6858), .C1(n1329), .Y(top_core_KE_sb1_n300) );
  OAI221XL U201 ( .A0(top_core_KE_sb1_n76), .A1(top_core_KE_sb1_n83), .B0(
        n1824), .B1(n78), .C0(top_core_KE_sb1_n293), .Y(top_core_KE_sb1_n291)
         );
  AOI211X1 U202 ( .A0(n11827), .A1(n1803), .B0(n11836), .C0(n243), .Y(n11835)
         );
  AOI211X1 U203 ( .A0(top_core_KE_sb1_n256), .A1(n1824), .B0(
        top_core_KE_sb1_n265), .C0(n242), .Y(top_core_KE_sb1_n264) );
  OAI222XL U204 ( .A0(n11718), .A1(n11705), .B0(n1803), .B1(n11716), .C0(n1350), .C1(n11735), .Y(n11731) );
  OAI222XL U205 ( .A0(n12034), .A1(n12021), .B0(n1782), .B1(n12032), .C0(n1366), .C1(n12051), .Y(n12047) );
  AOI222X1 U206 ( .A0(n6622), .A1(n12336), .B0(n6626), .B1(n1764), .C0(n6611), 
        .C1(n1264), .Y(n12502) );
  OAI221XL U207 ( .A0(n12283), .A1(n12290), .B0(n1761), .B1(n184), .C0(n12495), 
        .Y(n12493) );
  AOI222X1 U208 ( .A0(n6575), .A1(n12021), .B0(n6579), .B1(n1787), .C0(n6564), 
        .C1(n1260), .Y(n12187) );
  OAI221XL U209 ( .A0(n11967), .A1(n11974), .B0(n1782), .B1(n79), .C0(n12180), 
        .Y(n12178) );
  AOI211X1 U210 ( .A0(n12458), .A1(n1761), .B0(n12467), .C0(n241), .Y(n12466)
         );
  AOI211X1 U211 ( .A0(n12143), .A1(n1782), .B0(n12152), .C0(n240), .Y(n12151)
         );
  OAI222XL U212 ( .A0(n12349), .A1(n12336), .B0(n1761), .B1(n12347), .C0(n1364), .C1(n12366), .Y(n12362) );
  OAI221XL U213 ( .A0(n58), .A1(n13897), .B0(n14135), .B1(n13922), .C0(n13879), 
        .Y(n14139) );
  AOI222X1 U214 ( .A0(n1625), .A1(n585), .B0(n6156), .B1(n1327), .C0(n1139), 
        .C1(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n301) );
  AOI222X1 U215 ( .A0(n545), .A1(n3488), .B0(n6146), .B1(n1327), .C0(n1625), 
        .C1(n561), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n304) );
  NAND4BXL U216 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n106), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n108), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n234), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n228) );
  OAI221XL U217 ( .A0(n61), .A1(n15472), .B0(n15710), .B1(n15497), .C0(n15454), 
        .Y(n15714) );
  AOI222X1 U218 ( .A0(n1612), .A1(n589), .B0(n5096), .B1(n1251), .C0(n954), 
        .C1(n10846), .Y(n10991) );
  AOI222X1 U219 ( .A0(n549), .A1(n2705), .B0(n5080), .B1(n1251), .C0(n1612), 
        .C1(n565), .Y(n10994) );
  NAND4BXL U220 ( .AN(n10797), .B(n10799), .C(n10772), .D(n10924), .Y(n10918)
         );
  OAI221XL U221 ( .A0(n57), .A1(n17047), .B0(n17285), .B1(n17072), .C0(n17029), 
        .Y(n17289) );
  AOI222X1 U222 ( .A0(n1615), .A1(n586), .B0(n5366), .B1(n1245), .C0(n996), 
        .C1(n9970), .Y(n10115) );
  AOI222X1 U223 ( .A0(n546), .A1(n2888), .B0(n5350), .B1(n1245), .C0(n1615), 
        .C1(n562), .Y(n10118) );
  NAND4BXL U224 ( .AN(n9921), .B(n9923), .C(n9896), .D(n10048), .Y(n10042) );
  OAI221XL U225 ( .A0(n63), .A1(n18622), .B0(n18860), .B1(n18647), .C0(n18604), 
        .Y(n18864) );
  AOI222X1 U226 ( .A0(n1618), .A1(n590), .B0(n5602), .B1(n1239), .C0(n1038), 
        .C1(n9094), .Y(n9239) );
  AOI222X1 U227 ( .A0(n550), .A1(n3070), .B0(n5586), .B1(n1239), .C0(n1618), 
        .C1(n566), .Y(n9242) );
  NAND4BXL U228 ( .AN(n9045), .B(n9047), .C(n9020), .D(n9172), .Y(n9166) );
  OAI221XL U229 ( .A0(n60), .A1(n15157), .B0(n15395), .B1(n15182), .C0(n15139), 
        .Y(n15399) );
  AOI222X1 U230 ( .A0(n1621), .A1(n588), .B0(n5838), .B1(n1233), .C0(n1080), 
        .C1(n8218), .Y(n8363) );
  AOI222X1 U231 ( .A0(n548), .A1(n3245), .B0(n5822), .B1(n1233), .C0(n1621), 
        .C1(n564), .Y(n8366) );
  NAND4BXL U232 ( .AN(n8169), .B(n8171), .C(n8144), .D(n8296), .Y(n8290) );
  OAI221XL U233 ( .A0(n62), .A1(n16732), .B0(n16970), .B1(n16757), .C0(n16714), 
        .Y(n16974) );
  AOI222X1 U234 ( .A0(n1624), .A1(n591), .B0(n6066), .B1(n1227), .C0(n1122), 
        .C1(n7342), .Y(n7487) );
  AOI222X1 U235 ( .A0(n551), .A1(n3425), .B0(n6050), .B1(n1227), .C0(n1624), 
        .C1(n567), .Y(n7490) );
  NAND4BXL U236 ( .AN(n7293), .B(n7295), .C(n7268), .D(n7420), .Y(n7414) );
  OAI221XL U237 ( .A0(n59), .A1(n18307), .B0(n18545), .B1(n18332), .C0(n18289), 
        .Y(n18549) );
  AOI222X1 U238 ( .A0(n1611), .A1(n587), .B0(n5012), .B1(n1253), .C0(n940), 
        .C1(n11138), .Y(n11283) );
  AOI222X1 U239 ( .A0(n547), .A1(n2643), .B0(n4996), .B1(n1253), .C0(n1611), 
        .C1(n563), .Y(n11286) );
  NAND4BXL U240 ( .AN(n11089), .B(n11091), .C(n11064), .D(n11216), .Y(n11210)
         );
  OAI221XL U241 ( .A0(n64), .A1(n14842), .B0(n15080), .B1(n14867), .C0(n14824), 
        .Y(n15084) );
  AOI222X1 U242 ( .A0(n1614), .A1(n592), .B0(n5282), .B1(n1247), .C0(n982), 
        .C1(n10262), .Y(n10407) );
  AOI222X1 U243 ( .A0(n552), .A1(n2830), .B0(n5266), .B1(n1247), .C0(n1614), 
        .C1(n568), .Y(n10410) );
  NAND4BXL U244 ( .AN(n10213), .B(n10215), .C(n10188), .D(n10340), .Y(n10334)
         );
  OAI221XL U245 ( .A0(n65), .A1(n16417), .B0(n16655), .B1(n16442), .C0(n16399), 
        .Y(n16659) );
  AOI222X1 U246 ( .A0(n1617), .A1(n593), .B0(n5526), .B1(n1241), .C0(n1024), 
        .C1(n9386), .Y(n9531) );
  AOI222X1 U247 ( .A0(n553), .A1(n3007), .B0(n5510), .B1(n1241), .C0(n1617), 
        .C1(n569), .Y(n9534) );
  NAND4BXL U248 ( .AN(n9337), .B(n9339), .C(n9312), .D(n9464), .Y(n9458) );
  OAI221XL U249 ( .A0(n66), .A1(n17992), .B0(n18230), .B1(n18017), .C0(n17974), 
        .Y(n18234) );
  AOI222X1 U250 ( .A0(n1620), .A1(n594), .B0(n5754), .B1(n1235), .C0(n1066), 
        .C1(n8510), .Y(n8655) );
  AOI222X1 U251 ( .A0(n554), .A1(n3185), .B0(n5738), .B1(n1235), .C0(n1620), 
        .C1(n570), .Y(n8658) );
  NAND4BXL U252 ( .AN(n8461), .B(n8463), .C(n8436), .D(n8588), .Y(n8582) );
  OAI221XL U253 ( .A0(n67), .A1(n14527), .B0(n14765), .B1(n14552), .C0(n14509), 
        .Y(n14769) );
  AOI222X1 U254 ( .A0(n1623), .A1(n595), .B0(n5990), .B1(n1229), .C0(n1108), 
        .C1(n7634), .Y(n7779) );
  AOI222X1 U255 ( .A0(n555), .A1(n3368), .B0(n5974), .B1(n1229), .C0(n1623), 
        .C1(n571), .Y(n7782) );
  NAND4BXL U256 ( .AN(n7585), .B(n7587), .C(n7560), .D(n7712), .Y(n7706) );
  OAI221XL U257 ( .A0(n68), .A1(n16102), .B0(n16340), .B1(n16127), .C0(n16084), 
        .Y(n16344) );
  AOI222X1 U258 ( .A0(n1610), .A1(n596), .B0(n4896), .B1(n1255), .C0(n926), 
        .C1(n11430), .Y(n11575) );
  AOI222X1 U259 ( .A0(n556), .A1(n2583), .B0(n4880), .B1(n1255), .C0(n1610), 
        .C1(n572), .Y(n11578) );
  NAND4BXL U260 ( .AN(n11381), .B(n11383), .C(n11356), .D(n11508), .Y(n11502)
         );
  OAI221XL U261 ( .A0(n69), .A1(n17677), .B0(n17915), .B1(n17702), .C0(n17659), 
        .Y(n17919) );
  AOI222X1 U262 ( .A0(n1613), .A1(n597), .B0(n5204), .B1(n1249), .C0(n968), 
        .C1(n10554), .Y(n10699) );
  AOI222X1 U263 ( .A0(n557), .A1(n2765), .B0(n5188), .B1(n1249), .C0(n1613), 
        .C1(n573), .Y(n10702) );
  NAND4BXL U264 ( .AN(n10505), .B(n10507), .C(n10480), .D(n10632), .Y(n10626)
         );
  OAI221XL U265 ( .A0(n70), .A1(n14212), .B0(n14450), .B1(n14237), .C0(n14194), 
        .Y(n14454) );
  AOI222X1 U266 ( .A0(n1616), .A1(n598), .B0(n5450), .B1(n1243), .C0(n1010), 
        .C1(n9678), .Y(n9823) );
  AOI222X1 U267 ( .A0(n558), .A1(n2947), .B0(n5434), .B1(n1243), .C0(n1616), 
        .C1(n574), .Y(n9826) );
  NAND4BXL U268 ( .AN(n9629), .B(n9631), .C(n9604), .D(n9756), .Y(n9750) );
  OAI221XL U269 ( .A0(n71), .A1(n15787), .B0(n16025), .B1(n15812), .C0(n15769), 
        .Y(n16029) );
  AOI222X1 U270 ( .A0(n1619), .A1(n599), .B0(n5678), .B1(n1237), .C0(n1052), 
        .C1(n8802), .Y(n8947) );
  AOI222X1 U271 ( .A0(n559), .A1(n3127), .B0(n5662), .B1(n1237), .C0(n1619), 
        .C1(n575), .Y(n8950) );
  NAND4BXL U272 ( .AN(n8753), .B(n8755), .C(n8728), .D(n8880), .Y(n8874) );
  OAI221XL U273 ( .A0(n72), .A1(n17362), .B0(n17600), .B1(n17387), .C0(n17344), 
        .Y(n17604) );
  AOI222X1 U274 ( .A0(n1622), .A1(n600), .B0(n5914), .B1(n1231), .C0(n1094), 
        .C1(n7926), .Y(n8071) );
  AOI222X1 U275 ( .A0(n560), .A1(n3306), .B0(n5898), .B1(n1231), .C0(n1622), 
        .C1(n576), .Y(n8074) );
  NAND4BXL U276 ( .AN(n7877), .B(n7879), .C(n7852), .D(n8004), .Y(n7998) );
  OAI22X2 U277 ( .A0(n2533), .A1(top_core_EC_ss_n138), .B0(n2374), .B1(n122), 
        .Y(top_core_EC_mc_mix_in_8[95]) );
  OAI22X2 U278 ( .A0(n2532), .A1(top_core_EC_ss_n230), .B0(n2368), .B1(n129), 
        .Y(top_core_EC_mc_mix_in_8[127]) );
  AOI221X1 U279 ( .A0(n6597), .A1(n1278), .B0(n1157), .B1(n13538), .C0(n13708), 
        .Y(n13831) );
  OAI221XL U280 ( .A0(n13670), .A1(n13543), .B0(n1659), .B1(n55), .C0(n13665), 
        .Y(n13833) );
  OAI221XL U281 ( .A0(n6), .A1(n13583), .B0(n13820), .B1(n190), .C0(n13565), 
        .Y(n13824) );
  OAI221XL U282 ( .A0(n616), .A1(n6), .B0(n13610), .B1(n13553), .C0(n13784), 
        .Y(n13783) );
  OAI221XL U283 ( .A0(n695), .A1(n55), .B0(n13610), .B1(n1664), .C0(n13790), 
        .Y(n13785) );
  OAI221XL U284 ( .A0(n12598), .A1(n12605), .B0(n1739), .B1(n181), .C0(n12810), 
        .Y(n12808) );
  OAI221XL U285 ( .A0(n13543), .A1(n13550), .B0(n1652), .B1(n183), .C0(n13755), 
        .Y(n13753) );
  AOI211X1 U286 ( .A0(n12773), .A1(n1739), .B0(n12782), .C0(n262), .Y(n12781)
         );
  OAI221XL U287 ( .A0(n3), .A1(n13268), .B0(n13505), .B1(n187), .C0(n13250), 
        .Y(n13509) );
  AOI221X1 U288 ( .A0(n6890), .A1(n1272), .B0(n1197), .B1(n12908), .C0(n13078), 
        .Y(n13201) );
  OAI221XL U289 ( .A0(n13040), .A1(n12913), .B0(n1717), .B1(n56), .C0(n13035), 
        .Y(n13203) );
  OAI221XL U290 ( .A0(n5), .A1(n12953), .B0(n13190), .B1(n191), .C0(n12935), 
        .Y(n13194) );
  OAI221XL U291 ( .A0(n612), .A1(n5), .B0(n12980), .B1(n12923), .C0(n13154), 
        .Y(n13153) );
  OAI221XL U292 ( .A0(n696), .A1(n56), .B0(n12980), .B1(n1721), .C0(n13160), 
        .Y(n13155) );
  OAI221XL U293 ( .A0(n13228), .A1(n13235), .B0(n1681), .B1(n180), .C0(n13440), 
        .Y(n13438) );
  OAI221XL U294 ( .A0(n12913), .A1(n12920), .B0(n1710), .B1(n182), .C0(n13125), 
        .Y(n13123) );
  AOI211X1 U295 ( .A0(n13403), .A1(n1681), .B0(n13412), .C0(n263), .Y(n13411)
         );
  AOI211X1 U296 ( .A0(n13088), .A1(n1710), .B0(n13097), .C0(n260), .Y(n13096)
         );
  OAI222XL U297 ( .A0(n12980), .A1(n12967), .B0(n1710), .B1(n12978), .C0(n1351), .C1(n12997), .Y(n12993) );
  OAI222XL U298 ( .A0(n12665), .A1(n12652), .B0(n1739), .B1(n12663), .C0(n1353), .C1(n12682), .Y(n12678) );
  OAI221XL U299 ( .A0(n610), .A1(n3), .B0(n13295), .B1(n13238), .C0(n13469), 
        .Y(n13468) );
  AOI221X1 U300 ( .A0(n6844), .A1(n1269), .B0(n1188), .B1(n12593), .C0(n12763), 
        .Y(n12886) );
  OAI221XL U301 ( .A0(n12725), .A1(n12598), .B0(n1746), .B1(n54), .C0(n12720), 
        .Y(n12888) );
  OAI221XL U302 ( .A0(n4), .A1(n12638), .B0(n12875), .B1(n189), .C0(n12620), 
        .Y(n12879) );
  OAI221XL U303 ( .A0(n611), .A1(n4), .B0(n12665), .B1(n12608), .C0(n12839), 
        .Y(n12838) );
  OAI221XL U304 ( .A0(n694), .A1(n54), .B0(n12665), .B1(n1750), .C0(n12845), 
        .Y(n12840) );
  AOI211X1 U305 ( .A0(n13718), .A1(n1652), .B0(n13727), .C0(n261), .Y(n13726)
         );
  OAI222XL U306 ( .A0(n13610), .A1(n13597), .B0(n1652), .B1(n13608), .C0(n1365), .C1(n13627), .Y(n13623) );
  OAI22X2 U307 ( .A0(n2480), .A1(top_core_EC_ss_n209), .B0(n2369), .B1(n4836), 
        .Y(top_core_EC_mc_mix_in_8[31]) );
  OAI22X2 U308 ( .A0(n2460), .A1(top_core_EC_ss_n173), .B0(n2372), .B1(n128), 
        .Y(top_core_EC_mc_mix_in_8[63]) );
  CLKINVX3 U309 ( .A(n1713), .Y(n1710) );
  CLKINVX3 U310 ( .A(n1742), .Y(n1739) );
  CLKINVX3 U311 ( .A(n1684), .Y(n1681) );
  NOR2X2 U312 ( .A(top_core_KE_key_mem_ctrl_reg_0_), .B(n7017), .Y(
        top_core_KE_n2705) );
  OR2X2 U313 ( .A(n7020), .B(top_core_KE_n1865), .Y(n739) );
  AND2X2 U314 ( .A(top_core_KE_n896), .B(top_core_KE_n1865), .Y(n740) );
  INVX1 U315 ( .A(n_ADDR[1]), .Y(n4136) );
  NAND2X2 U316 ( .A(n2), .B(top_core_EC_n946), .Y(n1) );
  AND2X2 U317 ( .A(n1), .B(top_core_EC_n868), .Y(n742) );
  NAND2X2 U318 ( .A(top_core_t_ready), .B(n6308), .Y(n2) );
  NAND2X2 U319 ( .A(n1673), .B(n748), .Y(n3) );
  NAND2X2 U320 ( .A(n1731), .B(n749), .Y(n4) );
  NAND2X2 U321 ( .A(n1702), .B(n750), .Y(n5) );
  NAND2X2 U322 ( .A(n1648), .B(n751), .Y(n6) );
  INVX1 U323 ( .A(top_core_KE_n1873), .Y(n2253) );
  INVX1 U324 ( .A(top_core_KE_n1873), .Y(n2252) );
  NAND2X2 U325 ( .A(top_core_io_n233), .B(n85), .Y(n7) );
  NAND2X2 U326 ( .A(top_core_io_n60), .B(n85), .Y(n8) );
  NAND2X2 U327 ( .A(top_core_io_n222), .B(n85), .Y(n9) );
  NAND2X2 U328 ( .A(top_core_io_n211), .B(n85), .Y(n10) );
  NAND2X2 U329 ( .A(top_core_io_n200), .B(n85), .Y(n11) );
  NAND2X2 U330 ( .A(top_core_io_n38), .B(n85), .Y(n12) );
  AND2X2 U331 ( .A(top_core_io_n49), .B(n85), .Y(n13) );
  INVX1 U332 ( .A(n_ADDR[2]), .Y(n4140) );
  NAND2X4 U333 ( .A(n6165), .B(n3479), .Y(n14) );
  NAND2X4 U334 ( .A(n5375), .B(n2877), .Y(n15) );
  NAND2X4 U335 ( .A(n5021), .B(n2635), .Y(n16) );
  NAND2X4 U336 ( .A(n5847), .B(n3237), .Y(n17) );
  NAND2X4 U337 ( .A(n5105), .B(n2693), .Y(n18) );
  NAND2X4 U338 ( .A(n5611), .B(n3057), .Y(n19) );
  NAND2X4 U339 ( .A(n6075), .B(n3414), .Y(n20) );
  NAND2X4 U340 ( .A(n5291), .B(n2816), .Y(n21) );
  NAND2X4 U341 ( .A(n5535), .B(n2996), .Y(n22) );
  NAND2X4 U342 ( .A(n5763), .B(n3176), .Y(n23) );
  NAND2X4 U343 ( .A(n5999), .B(n3359), .Y(n24) );
  NAND2X4 U344 ( .A(n4905), .B(n2574), .Y(n25) );
  NAND2X4 U345 ( .A(n5213), .B(n2756), .Y(n26) );
  NAND2X4 U346 ( .A(n5459), .B(n2935), .Y(n27) );
  NAND2X4 U347 ( .A(n5687), .B(n3118), .Y(n28) );
  NAND2X4 U348 ( .A(n5923), .B(n3297), .Y(n29) );
  AND2X2 U349 ( .A(n17017), .B(n1310), .Y(n337) );
  CLKBUFX3 U350 ( .A(n337), .Y(n1003) );
  AND2X2 U351 ( .A(n13867), .B(n1280), .Y(n338) );
  CLKBUFX3 U352 ( .A(n338), .Y(n1142) );
  AND2X2 U353 ( .A(n15127), .B(n1292), .Y(n340) );
  CLKBUFX3 U354 ( .A(n340), .Y(n1087) );
  AND2X2 U355 ( .A(n18277), .B(n1322), .Y(n339) );
  CLKBUFX3 U356 ( .A(n339), .Y(n947) );
  AND2X2 U357 ( .A(n15442), .B(n1295), .Y(n341) );
  CLKBUFX3 U358 ( .A(n341), .Y(n1073) );
  AND2X2 U359 ( .A(n16702), .B(n1307), .Y(n342) );
  CLKBUFX3 U360 ( .A(n342), .Y(n1017) );
  AND2X2 U361 ( .A(n18592), .B(n1325), .Y(n343) );
  CLKBUFX3 U362 ( .A(n343), .Y(n933) );
  AND2X2 U363 ( .A(n14812), .B(n1289), .Y(n344) );
  CLKBUFX3 U364 ( .A(n344), .Y(n1101) );
  AND2X2 U365 ( .A(n16387), .B(n1304), .Y(n345) );
  CLKBUFX3 U366 ( .A(n345), .Y(n1031) );
  AND2X2 U367 ( .A(n17962), .B(n1319), .Y(n346) );
  CLKBUFX3 U368 ( .A(n346), .Y(n961) );
  AND2X2 U369 ( .A(n14497), .B(n1286), .Y(n347) );
  CLKBUFX3 U370 ( .A(n347), .Y(n1115) );
  AND2X2 U371 ( .A(n16072), .B(n1301), .Y(n348) );
  CLKBUFX3 U372 ( .A(n348), .Y(n1045) );
  AND2X2 U373 ( .A(n17647), .B(n1316), .Y(n349) );
  CLKBUFX3 U374 ( .A(n349), .Y(n975) );
  AND2X2 U375 ( .A(n14182), .B(n1283), .Y(n350) );
  CLKBUFX3 U376 ( .A(n350), .Y(n1129) );
  AND2X2 U377 ( .A(n15757), .B(n1298), .Y(n351) );
  CLKBUFX3 U378 ( .A(n351), .Y(n1059) );
  AND2X2 U379 ( .A(n17332), .B(n1313), .Y(n352) );
  CLKBUFX3 U380 ( .A(n352), .Y(n989) );
  NAND2X2 U381 ( .A(top_core_EC_ss_in[82]), .B(n995), .Y(n30) );
  NAND2X2 U382 ( .A(n3477), .B(n1134), .Y(n31) );
  NAND2X2 U383 ( .A(top_core_EC_ss_in[114]), .B(n939), .Y(n32) );
  NAND2X2 U384 ( .A(top_core_EC_ss_in[34]), .B(n1079), .Y(n33) );
  NAND2X2 U385 ( .A(top_core_EC_ss_in[42]), .B(n1065), .Y(n34) );
  NAND2X2 U386 ( .A(top_core_EC_ss_in[122]), .B(n925), .Y(n35) );
  NAND2X2 U387 ( .A(top_core_EC_ss_in[74]), .B(n1009), .Y(n36) );
  NAND2X2 U388 ( .A(top_core_EC_ss_in[26]), .B(n1093), .Y(n37) );
  NAND2X2 U389 ( .A(top_core_EC_ss_in[66]), .B(n1023), .Y(n38) );
  NAND2X2 U390 ( .A(top_core_EC_ss_in[106]), .B(n953), .Y(n39) );
  NAND2X2 U391 ( .A(top_core_EC_ss_in[18]), .B(n1107), .Y(n40) );
  NAND2X2 U392 ( .A(top_core_EC_ss_in[58]), .B(n1037), .Y(n41) );
  NAND2X2 U393 ( .A(top_core_EC_ss_in[98]), .B(n967), .Y(n42) );
  NAND2X2 U394 ( .A(top_core_EC_ss_in[10]), .B(n1121), .Y(n43) );
  NAND2X2 U395 ( .A(top_core_EC_ss_in[50]), .B(n1051), .Y(n44) );
  NAND2X2 U396 ( .A(top_core_EC_ss_in[90]), .B(n981), .Y(n45) );
  NAND2X2 U397 ( .A(n1360), .B(n1164), .Y(n46) );
  NAND2X2 U398 ( .A(top_core_io_n528), .B(n85), .Y(n47) );
  NAND2X2 U399 ( .A(top_core_io_n517), .B(n85), .Y(n48) );
  NAND2X2 U400 ( .A(top_core_io_n506), .B(n85), .Y(n49) );
  NAND2X4 U401 ( .A(n1209), .B(n1204), .Y(n50) );
  NAND2X4 U402 ( .A(n1207), .B(n1195), .Y(n51) );
  NAND2X4 U403 ( .A(n1166), .B(n1150), .Y(n52) );
  NAND2X4 U404 ( .A(n1167), .B(n1155), .Y(n53) );
  NAND2X4 U405 ( .A(n1206), .B(n1190), .Y(n54) );
  NAND2X4 U406 ( .A(n1168), .B(n1159), .Y(n55) );
  NAND2X4 U407 ( .A(n1208), .B(n1199), .Y(n56) );
  NAND2X2 U408 ( .A(n2875), .B(n5375), .Y(n57) );
  NAND2X2 U409 ( .A(n3475), .B(n6165), .Y(n58) );
  NAND2X2 U410 ( .A(n2633), .B(n5021), .Y(n59) );
  NAND2X2 U411 ( .A(n3236), .B(n5847), .Y(n60) );
  NAND2X2 U412 ( .A(n3175), .B(n5763), .Y(n61) );
  NAND2X2 U413 ( .A(n2936), .B(n5459), .Y(n62) );
  NAND2X2 U414 ( .A(n2572), .B(n4905), .Y(n63) );
  NAND2X2 U415 ( .A(n3297), .B(n5923), .Y(n64) );
  NAND2X2 U416 ( .A(n2997), .B(n5535), .Y(n65) );
  NAND2X2 U417 ( .A(n2694), .B(n5105), .Y(n66) );
  NAND2X2 U418 ( .A(n3358), .B(n5999), .Y(n67) );
  NAND2X2 U419 ( .A(n3055), .B(n5611), .Y(n68) );
  NAND2X2 U420 ( .A(n2755), .B(n5213), .Y(n69) );
  NAND2X2 U421 ( .A(n3415), .B(n6075), .Y(n70) );
  NAND2X2 U422 ( .A(n3116), .B(n5687), .Y(n71) );
  NAND2X2 U423 ( .A(n2816), .B(n5291), .Y(n72) );
  AND2X2 U424 ( .A(n1273), .B(n1274), .Y(n580) );
  CLKBUFX3 U425 ( .A(n580), .Y(n1173) );
  AND2X2 U426 ( .A(n1267), .B(n1268), .Y(n584) );
  CLKBUFX3 U427 ( .A(n584), .Y(n1213) );
  AND2X2 U428 ( .A(n1276), .B(n1277), .Y(n583) );
  CLKBUFX3 U429 ( .A(n583), .Y(n1178) );
  AND2X2 U430 ( .A(n1270), .B(n1271), .Y(n582) );
  CLKBUFX3 U431 ( .A(n582), .Y(n1219) );
  AND2X2 U432 ( .A(n1257), .B(n1258), .Y(n577) );
  CLKBUFX3 U433 ( .A(n577), .Y(n1222) );
  AND2X2 U434 ( .A(n1329), .B(n1330), .Y(n578) );
  CLKBUFX3 U435 ( .A(n578), .Y(n1216) );
  AND2X2 U436 ( .A(n1263), .B(n1265), .Y(n579) );
  CLKBUFX3 U437 ( .A(n579), .Y(n1181) );
  AND2X2 U438 ( .A(n1260), .B(n1261), .Y(n581) );
  CLKBUFX3 U439 ( .A(n581), .Y(n1176) );
  NAND2X2 U440 ( .A(n1673), .B(n1149), .Y(n73) );
  NAND2X2 U441 ( .A(n1731), .B(n1189), .Y(n74) );
  NAND2X2 U442 ( .A(n1702), .B(n1198), .Y(n75) );
  NAND2X2 U443 ( .A(n1646), .B(n1158), .Y(n76) );
  NAND2X2 U444 ( .A(n1344), .B(n761), .Y(n77) );
  NAND2X2 U445 ( .A(n1345), .B(n762), .Y(n78) );
  NAND2X2 U446 ( .A(n1359), .B(n763), .Y(n79) );
  NAND2X2 U447 ( .A(n1344), .B(n1203), .Y(n80) );
  NAND2X2 U448 ( .A(n1345), .B(n1194), .Y(n81) );
  NAND2X2 U449 ( .A(n1358), .B(n1163), .Y(n82) );
  NAND2X2 U450 ( .A(n1359), .B(n1154), .Y(n83) );
  NAND2X2 U451 ( .A(top_core_io_n222), .B(n303), .Y(n84) );
  NOR2X4 U452 ( .A(n4143), .B(n4140), .Y(n85) );
  NOR2X4 U453 ( .A(n4138), .B(n4142), .Y(n86) );
  NAND2X2 U454 ( .A(top_core_io_n495), .B(n85), .Y(n87) );
  NAND2X2 U455 ( .A(n85), .B(top_core_io_n27), .Y(n88) );
  NAND2X4 U456 ( .A(n1169), .B(n1164), .Y(n89) );
  NAND2X4 U457 ( .A(n5348), .B(n2876), .Y(n90) );
  NAND2X4 U458 ( .A(n6144), .B(n3479), .Y(n91) );
  NAND2X4 U459 ( .A(n4994), .B(n2634), .Y(n92) );
  NAND2X4 U460 ( .A(n5820), .B(n3236), .Y(n93) );
  NAND2X4 U461 ( .A(n5078), .B(n2695), .Y(n94) );
  NAND2X4 U462 ( .A(n6048), .B(n3416), .Y(n95) );
  NAND2X4 U463 ( .A(n5584), .B(n3056), .Y(n96) );
  NAND2X4 U464 ( .A(n5264), .B(n2815), .Y(n97) );
  NAND2X4 U465 ( .A(n5508), .B(n2998), .Y(n98) );
  NAND2X4 U466 ( .A(n5736), .B(n3175), .Y(n99) );
  NAND2X4 U467 ( .A(n5972), .B(n3358), .Y(n100) );
  NAND2X4 U468 ( .A(n4878), .B(n2573), .Y(n101) );
  NAND2X4 U469 ( .A(n5186), .B(n2755), .Y(n102) );
  NAND2X4 U470 ( .A(n5432), .B(n2937), .Y(n103) );
  NAND2X4 U471 ( .A(n5660), .B(n3117), .Y(n104) );
  NAND2X4 U472 ( .A(n5896), .B(n3296), .Y(n105) );
  NAND2X4 U473 ( .A(n1000), .B(n2868), .Y(n106) );
  NAND2X4 U474 ( .A(n1140), .B(n3470), .Y(n107) );
  NAND2X4 U475 ( .A(n944), .B(n2626), .Y(n108) );
  NAND2X4 U476 ( .A(n1084), .B(n3228), .Y(n109) );
  NAND2X4 U477 ( .A(n1070), .B(n3167), .Y(n110) );
  NAND2X4 U478 ( .A(n930), .B(n2565), .Y(n111) );
  NAND2X4 U479 ( .A(n1014), .B(n2929), .Y(n112) );
  NAND2X4 U480 ( .A(n1098), .B(n3289), .Y(n113) );
  NAND2X4 U481 ( .A(n1028), .B(n2990), .Y(n114) );
  NAND2X4 U482 ( .A(n958), .B(n2689), .Y(n115) );
  NAND2X4 U483 ( .A(n1112), .B(n3350), .Y(n116) );
  NAND2X4 U484 ( .A(n1042), .B(n3048), .Y(n117) );
  NAND2X4 U485 ( .A(n972), .B(n2747), .Y(n118) );
  NAND2X4 U486 ( .A(n1126), .B(n3408), .Y(n119) );
  NAND2X4 U487 ( .A(n1056), .B(n3109), .Y(n120) );
  NAND2X4 U488 ( .A(n986), .B(n2808), .Y(n121) );
  XNOR2X1 U489 ( .A(top_core_Key[36]), .B(top_core_EC_add_in_r[92]), .Y(n122)
         );
  XNOR2X1 U490 ( .A(top_core_Key[47]), .B(top_core_EC_add_in_r[87]), .Y(n123)
         );
  XNOR2X1 U491 ( .A(top_core_Key[46]), .B(top_core_EC_add_in_r[86]), .Y(n124)
         );
  XNOR2X1 U492 ( .A(top_core_Key[45]), .B(top_core_EC_add_in_r[85]), .Y(n125)
         );
  XNOR2X1 U493 ( .A(top_core_Key[62]), .B(top_core_EC_add_in_r[70]), .Y(n126)
         );
  XNOR2X1 U494 ( .A(top_core_Key[61]), .B(top_core_EC_add_in_r[69]), .Y(n127)
         );
  XNOR2X1 U495 ( .A(top_core_Key[68]), .B(top_core_EC_add_in_r[60]), .Y(n128)
         );
  XNOR2X1 U496 ( .A(top_core_Key[4]), .B(top_core_EC_add_in_r[124]), .Y(n129)
         );
  XNOR2X1 U497 ( .A(top_core_Key[15]), .B(top_core_EC_add_in_r[119]), .Y(n130)
         );
  XNOR2X1 U498 ( .A(top_core_Key[14]), .B(top_core_EC_add_in_r[118]), .Y(n131)
         );
  XNOR2X1 U499 ( .A(top_core_Key[13]), .B(top_core_EC_add_in_r[117]), .Y(n132)
         );
  XNOR2X1 U500 ( .A(top_core_Key[30]), .B(top_core_EC_add_in_r[102]), .Y(n133)
         );
  XNOR2X1 U501 ( .A(top_core_Key[29]), .B(top_core_EC_add_in_r[101]), .Y(n134)
         );
  NOR2X2 U502 ( .A(n2874), .B(n2866), .Y(n135) );
  NOR2X2 U503 ( .A(n3476), .B(n3467), .Y(n136) );
  NOR2X2 U504 ( .A(n2632), .B(n2624), .Y(n137) );
  NOR2X2 U505 ( .A(n3235), .B(n3226), .Y(n138) );
  NOR2X2 U506 ( .A(n2693), .B(n2685), .Y(n139) );
  NOR2X2 U507 ( .A(n3054), .B(n3046), .Y(n140) );
  NOR2X2 U508 ( .A(n3414), .B(n3406), .Y(n141) );
  NOR2X2 U509 ( .A(n2814), .B(n2806), .Y(n142) );
  NOR2X2 U510 ( .A(n2996), .B(n2988), .Y(n143) );
  NOR2X2 U511 ( .A(n3174), .B(n3165), .Y(n144) );
  NOR2X2 U512 ( .A(n3357), .B(n3348), .Y(n145) );
  NOR2X2 U513 ( .A(n2571), .B(n2563), .Y(n146) );
  NOR2X2 U514 ( .A(n2754), .B(n2745), .Y(n147) );
  NOR2X2 U515 ( .A(n2935), .B(n2927), .Y(n148) );
  NOR2X2 U516 ( .A(n3115), .B(n3107), .Y(n149) );
  NOR2X2 U517 ( .A(n3295), .B(n3287), .Y(n150) );
  NAND2X2 U518 ( .A(top_core_KE_n2705), .B(n1500), .Y(n151) );
  XNOR2X1 U519 ( .A(top_core_Key[60]), .B(top_core_EC_add_in_r[68]), .Y(n152)
         );
  XNOR2X1 U520 ( .A(top_core_Key[63]), .B(top_core_EC_add_in_r[71]), .Y(n153)
         );
  XNOR2X1 U521 ( .A(top_core_Key[49]), .B(top_core_EC_add_in_r[73]), .Y(n154)
         );
  XNOR2X1 U522 ( .A(top_core_Key[52]), .B(top_core_EC_add_in_r[76]), .Y(n155)
         );
  XNOR2X1 U523 ( .A(top_core_Key[44]), .B(top_core_EC_add_in_r[84]), .Y(n156)
         );
  XNOR2X1 U524 ( .A(top_core_Key[33]), .B(top_core_EC_add_in_r[89]), .Y(n157)
         );
  XNOR2X1 U525 ( .A(top_core_Key[28]), .B(top_core_EC_add_in_r[100]), .Y(n158)
         );
  XNOR2X1 U526 ( .A(top_core_Key[31]), .B(top_core_EC_add_in_r[103]), .Y(n159)
         );
  XNOR2X1 U527 ( .A(top_core_Key[17]), .B(top_core_EC_add_in_r[105]), .Y(n160)
         );
  XNOR2X1 U528 ( .A(top_core_Key[20]), .B(top_core_EC_add_in_r[108]), .Y(n161)
         );
  XNOR2X1 U529 ( .A(top_core_Key[12]), .B(top_core_EC_add_in_r[116]), .Y(n162)
         );
  XNOR2X1 U530 ( .A(top_core_Key[1]), .B(top_core_EC_add_in_r[121]), .Y(n163)
         );
  NAND2X2 U531 ( .A(n2878), .B(n999), .Y(n164) );
  NAND2X2 U532 ( .A(n3477), .B(n1138), .Y(n165) );
  NAND2X2 U533 ( .A(n2636), .B(n943), .Y(n166) );
  NAND2X2 U534 ( .A(n3238), .B(n1083), .Y(n167) );
  NAND2X2 U535 ( .A(n3177), .B(n1069), .Y(n168) );
  NAND2X2 U536 ( .A(n2575), .B(n929), .Y(n169) );
  NAND2X2 U537 ( .A(n2939), .B(n1013), .Y(n170) );
  NAND2X2 U538 ( .A(n3299), .B(n1097), .Y(n171) );
  NAND2X2 U539 ( .A(n3000), .B(n1027), .Y(n172) );
  NAND2X2 U540 ( .A(n2697), .B(n957), .Y(n173) );
  NAND2X2 U541 ( .A(n3360), .B(n1111), .Y(n174) );
  NAND2X2 U542 ( .A(n3058), .B(n1041), .Y(n175) );
  NAND2X2 U543 ( .A(n2757), .B(n971), .Y(n176) );
  NAND2X2 U544 ( .A(n3418), .B(n1125), .Y(n177) );
  NAND2X2 U545 ( .A(n3119), .B(n1055), .Y(n178) );
  NAND2X2 U546 ( .A(n2818), .B(n985), .Y(n179) );
  NAND2X2 U547 ( .A(n1673), .B(n756), .Y(n180) );
  NAND2X2 U548 ( .A(n1731), .B(n757), .Y(n181) );
  NAND2X2 U549 ( .A(n1702), .B(n758), .Y(n182) );
  NAND2X2 U550 ( .A(n1645), .B(n759), .Y(n183) );
  NAND2X2 U551 ( .A(n1358), .B(n760), .Y(n184) );
  NAND2X2 U552 ( .A(n1346), .B(n1204), .Y(n185) );
  NAND2X2 U553 ( .A(n1348), .B(n1195), .Y(n186) );
  NAND2X2 U554 ( .A(n1363), .B(n1150), .Y(n187) );
  NAND2X2 U555 ( .A(n1362), .B(n1155), .Y(n188) );
  NAND2X2 U556 ( .A(n1349), .B(n1190), .Y(n189) );
  NAND2X2 U557 ( .A(n1361), .B(n1159), .Y(n190) );
  NAND2X2 U558 ( .A(n1347), .B(n1199), .Y(n191) );
  XNOR2X1 U559 ( .A(top_core_Key[66]), .B(top_core_EC_add_in_r[58]), .Y(n192)
         );
  XNOR2X1 U560 ( .A(top_core_Key[67]), .B(top_core_EC_add_in_r[59]), .Y(n193)
         );
  XNOR2X1 U561 ( .A(top_core_Key[69]), .B(top_core_EC_add_in_r[61]), .Y(n194)
         );
  XNOR2X1 U562 ( .A(top_core_Key[70]), .B(top_core_EC_add_in_r[62]), .Y(n195)
         );
  XNOR2X1 U563 ( .A(top_core_Key[71]), .B(top_core_EC_add_in_r[63]), .Y(n196)
         );
  XNOR2X1 U564 ( .A(top_core_Key[56]), .B(top_core_EC_add_in_r[64]), .Y(n197)
         );
  XNOR2X1 U565 ( .A(top_core_Key[57]), .B(top_core_EC_add_in_r[65]), .Y(n198)
         );
  XNOR2X1 U566 ( .A(top_core_Key[58]), .B(top_core_EC_add_in_r[66]), .Y(n199)
         );
  XNOR2X1 U567 ( .A(top_core_Key[59]), .B(top_core_EC_add_in_r[67]), .Y(n200)
         );
  XNOR2X1 U568 ( .A(top_core_Key[48]), .B(top_core_EC_add_in_r[72]), .Y(n201)
         );
  XNOR2X1 U569 ( .A(top_core_Key[50]), .B(top_core_EC_add_in_r[74]), .Y(n202)
         );
  XNOR2X1 U570 ( .A(top_core_Key[51]), .B(top_core_EC_add_in_r[75]), .Y(n203)
         );
  XNOR2X1 U571 ( .A(top_core_Key[53]), .B(top_core_EC_add_in_r[77]), .Y(n204)
         );
  XNOR2X1 U572 ( .A(top_core_Key[54]), .B(top_core_EC_add_in_r[78]), .Y(n205)
         );
  XNOR2X1 U573 ( .A(top_core_Key[55]), .B(top_core_EC_add_in_r[79]), .Y(n206)
         );
  XNOR2X1 U574 ( .A(top_core_Key[40]), .B(top_core_EC_add_in_r[80]), .Y(n207)
         );
  XNOR2X1 U575 ( .A(top_core_Key[41]), .B(top_core_EC_add_in_r[81]), .Y(n208)
         );
  XNOR2X1 U576 ( .A(top_core_Key[42]), .B(top_core_EC_add_in_r[82]), .Y(n209)
         );
  XNOR2X1 U577 ( .A(top_core_Key[43]), .B(top_core_EC_add_in_r[83]), .Y(n210)
         );
  XNOR2X1 U578 ( .A(top_core_Key[32]), .B(top_core_EC_add_in_r[88]), .Y(n211)
         );
  XNOR2X1 U579 ( .A(top_core_Key[34]), .B(top_core_EC_add_in_r[90]), .Y(n212)
         );
  XNOR2X1 U580 ( .A(top_core_Key[35]), .B(top_core_EC_add_in_r[91]), .Y(n213)
         );
  XNOR2X1 U581 ( .A(top_core_Key[37]), .B(top_core_EC_add_in_r[93]), .Y(n214)
         );
  XNOR2X1 U582 ( .A(top_core_Key[38]), .B(top_core_EC_add_in_r[94]), .Y(n215)
         );
  XNOR2X1 U583 ( .A(top_core_Key[39]), .B(top_core_EC_add_in_r[95]), .Y(n216)
         );
  XNOR2X1 U584 ( .A(top_core_Key[24]), .B(top_core_EC_add_in_r[96]), .Y(n217)
         );
  XNOR2X1 U585 ( .A(top_core_Key[25]), .B(top_core_EC_add_in_r[97]), .Y(n218)
         );
  XNOR2X1 U586 ( .A(top_core_Key[26]), .B(top_core_EC_add_in_r[98]), .Y(n219)
         );
  XNOR2X1 U587 ( .A(top_core_Key[27]), .B(top_core_EC_add_in_r[99]), .Y(n220)
         );
  XNOR2X1 U588 ( .A(top_core_Key[16]), .B(top_core_EC_add_in_r[104]), .Y(n221)
         );
  XNOR2X1 U589 ( .A(top_core_Key[18]), .B(top_core_EC_add_in_r[106]), .Y(n222)
         );
  XNOR2X1 U590 ( .A(top_core_Key[19]), .B(top_core_EC_add_in_r[107]), .Y(n223)
         );
  XNOR2X1 U591 ( .A(top_core_Key[21]), .B(top_core_EC_add_in_r[109]), .Y(n224)
         );
  XNOR2X1 U592 ( .A(top_core_Key[22]), .B(top_core_EC_add_in_r[110]), .Y(n225)
         );
  XNOR2X1 U593 ( .A(top_core_Key[23]), .B(top_core_EC_add_in_r[111]), .Y(n226)
         );
  XNOR2X1 U594 ( .A(top_core_Key[8]), .B(top_core_EC_add_in_r[112]), .Y(n227)
         );
  XNOR2X1 U595 ( .A(top_core_Key[9]), .B(top_core_EC_add_in_r[113]), .Y(n228)
         );
  XNOR2X1 U596 ( .A(top_core_Key[10]), .B(top_core_EC_add_in_r[114]), .Y(n229)
         );
  XNOR2X1 U597 ( .A(top_core_Key[11]), .B(top_core_EC_add_in_r[115]), .Y(n230)
         );
  XNOR2X1 U598 ( .A(top_core_Key[0]), .B(top_core_EC_add_in_r[120]), .Y(n231)
         );
  XNOR2X1 U599 ( .A(top_core_Key[2]), .B(top_core_EC_add_in_r[122]), .Y(n232)
         );
  XNOR2X1 U600 ( .A(top_core_Key[3]), .B(top_core_EC_add_in_r[123]), .Y(n233)
         );
  XNOR2X1 U601 ( .A(top_core_Key[5]), .B(top_core_EC_add_in_r[125]), .Y(n234)
         );
  XNOR2X1 U602 ( .A(top_core_Key[6]), .B(top_core_EC_add_in_r[126]), .Y(n235)
         );
  XNOR2X1 U603 ( .A(top_core_Key[7]), .B(top_core_EC_add_in_r[127]), .Y(n236)
         );
  NOR2X1 U604 ( .A(n2385), .B(n6306), .Y(n237) );
  AND2X2 U605 ( .A(n2389), .B(n6305), .Y(n238) );
  CLKINVX3 U606 ( .A(n681), .Y(n11705) );
  CLKINVX3 U607 ( .A(n682), .Y(top_core_KE_sb1_n130) );
  CLKINVX3 U608 ( .A(n683), .Y(n12336) );
  CLKINVX3 U609 ( .A(n684), .Y(n12021) );
  CLKINVX3 U610 ( .A(n757), .Y(n12665) );
  CLKINVX3 U611 ( .A(n758), .Y(n12980) );
  CLKINVX3 U612 ( .A(n759), .Y(n13610) );
  NAND2X2 U613 ( .A(top_core_io_n506), .B(n86), .Y(n276) );
  NAND2X2 U614 ( .A(top_core_io_n495), .B(n86), .Y(n277) );
  NAND2X2 U615 ( .A(n302), .B(top_core_io_n49), .Y(n299) );
  NAND2X2 U616 ( .A(n302), .B(top_core_io_n38), .Y(n300) );
  NAND2X2 U617 ( .A(n302), .B(top_core_io_n27), .Y(n301) );
  AOI211X1 U618 ( .A0(n1099), .A1(n7952), .B0(n8057), .C0(n8011), .Y(n8056) );
  NOR2X1 U619 ( .A(n7852), .B(n3313), .Y(n8057) );
  AOI211X1 U620 ( .A0(n1015), .A1(n9704), .B0(n9809), .C0(n9763), .Y(n9808) );
  NOR2X1 U621 ( .A(n9604), .B(n2953), .Y(n9809) );
  AOI211X1 U622 ( .A0(n931), .A1(n11456), .B0(n11561), .C0(n11515), .Y(n11560)
         );
  NOR2X1 U623 ( .A(n11356), .B(n2589), .Y(n11561) );
  AOI211X1 U624 ( .A0(n1071), .A1(n8536), .B0(n8641), .C0(n8595), .Y(n8640) );
  NOR2X1 U625 ( .A(n8436), .B(n3191), .Y(n8641) );
  AOI211X1 U626 ( .A0(n987), .A1(n10288), .B0(n10393), .C0(n10347), .Y(n10392)
         );
  NOR2X1 U627 ( .A(n10188), .B(n2832), .Y(n10393) );
  AOI211X1 U628 ( .A0(n1127), .A1(n7368), .B0(n7473), .C0(n7427), .Y(n7472) );
  NOR2X1 U629 ( .A(n7268), .B(n3432), .Y(n7473) );
  AOI211X1 U630 ( .A0(n1043), .A1(n9120), .B0(n9225), .C0(n9179), .Y(n9224) );
  NOR2X1 U631 ( .A(n9020), .B(n3082), .Y(n9225) );
  AOI211X1 U632 ( .A0(n959), .A1(n10872), .B0(n10977), .C0(n10931), .Y(n10976)
         );
  NOR2X1 U633 ( .A(n10772), .B(n2710), .Y(n10977) );
  AOI211X1 U634 ( .A0(n1085), .A1(n8244), .B0(n8349), .C0(n8303), .Y(n8348) );
  NOR2X1 U635 ( .A(n8144), .B(n3252), .Y(n8349) );
  AOI211X1 U636 ( .A0(n945), .A1(n11164), .B0(n11269), .C0(n11223), .Y(n11268)
         );
  NOR2X1 U637 ( .A(n11064), .B(n2660), .Y(n11269) );
  AOI211X1 U638 ( .A0(n1001), .A1(n9996), .B0(n10101), .C0(n10055), .Y(n10100)
         );
  NOR2X1 U639 ( .A(n9896), .B(n2892), .Y(n10101) );
  AOI211X1 U640 ( .A0(n1143), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n182), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n287), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n241), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n286) );
  NOR2X1 U641 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .B(n3493), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n287) );
  AOI211X1 U642 ( .A0(n1057), .A1(n8828), .B0(n8933), .C0(n8887), .Y(n8932) );
  NOR2X1 U643 ( .A(n8728), .B(n3133), .Y(n8933) );
  AOI211X1 U644 ( .A0(n1113), .A1(n7660), .B0(n7765), .C0(n7719), .Y(n7764) );
  NOR2X1 U645 ( .A(n7560), .B(n3374), .Y(n7765) );
  AOI211X1 U646 ( .A0(n1029), .A1(n9412), .B0(n9517), .C0(n9471), .Y(n9516) );
  NOR2X1 U647 ( .A(n9312), .B(n3014), .Y(n9517) );
  AOI211X1 U648 ( .A0(n973), .A1(n10580), .B0(n10685), .C0(n10639), .Y(n10684)
         );
  NOR2X1 U649 ( .A(n10480), .B(n2771), .Y(n10685) );
  AOI222X1 U650 ( .A0(n1180), .A1(n6604), .B0(n13553), .B1(n13555), .C0(n13583), .C1(n6587), .Y(n13580) );
  OAI222XL U651 ( .A0(n13543), .A1(n76), .B0(n1178), .B1(n13743), .C0(n13670), 
        .C1(n13553), .Y(n13756) );
  AOI222X1 U652 ( .A0(n1161), .A1(n1278), .B0(n6592), .B1(n13553), .C0(n1157), 
        .C1(n13583), .Y(n13815) );
  CLKINVX3 U653 ( .A(n616), .Y(n13553) );
  NAND2X2 U654 ( .A(n302), .B(top_core_io_n60), .Y(n298) );
  NAND2X2 U655 ( .A(top_core_io_n517), .B(n86), .Y(n275) );
  AOI32X1 U656 ( .A0(n16811), .A1(n1306), .A2(n16693), .B0(n5411), .B1(n2964), 
        .Y(n16810) );
  OAI222XL U657 ( .A0(n414), .A1(n62), .B0(n2954), .B1(n36), .C0(n16757), .C1(
        n1306), .Y(n16941) );
  AOI221X1 U658 ( .A0(n5464), .A1(n16702), .B0(n1012), .B1(n1307), .C0(n16703), 
        .Y(n16701) );
  AOI32X1 U659 ( .A0(n13661), .A1(n1276), .A2(n13544), .B0(n6516), .B1(n1659), 
        .Y(n13660) );
  OAI222XL U660 ( .A0(n695), .A1(n6), .B0(n1659), .B1(n76), .C0(n190), .C1(
        n1276), .Y(n13791) );
  AOI221X1 U661 ( .A0(n6604), .A1(n1276), .B0(n1161), .B1(n13538), .C0(n13554), 
        .Y(n13552) );
  CLKINVX3 U662 ( .A(n609), .Y(n1276) );
  AOI32X1 U663 ( .A0(n13976), .A1(n1279), .A2(n13858), .B0(n6111), .B1(n3505), 
        .Y(n13975) );
  OAI222XL U664 ( .A0(n402), .A1(n58), .B0(n3494), .B1(n31), .C0(n13922), .C1(
        n1279), .Y(n14106) );
  AOI221X1 U665 ( .A0(n6151), .A1(n13867), .B0(n1137), .B1(n1280), .C0(n13868), 
        .Y(n13866) );
  AOI32X1 U666 ( .A0(n15236), .A1(n1291), .A2(n15118), .B0(n5799), .B1(n3263), 
        .Y(n15235) );
  OAI222XL U667 ( .A0(n404), .A1(n60), .B0(n3253), .B1(n33), .C0(n15182), .C1(
        n1291), .Y(n15366) );
  AOI221X1 U668 ( .A0(n5852), .A1(n15127), .B0(n1082), .B1(n1292), .C0(n15128), 
        .Y(n15126) );
  AOI32X1 U669 ( .A0(n18386), .A1(n1321), .A2(n18268), .B0(n4973), .B1(n2651), 
        .Y(n18385) );
  OAI222XL U670 ( .A0(n403), .A1(n59), .B0(n2650), .B1(n32), .C0(n18332), .C1(
        n1321), .Y(n18516) );
  AOI221X1 U671 ( .A0(n5026), .A1(n18277), .B0(n942), .B1(n1322), .C0(n18278), 
        .Y(n18276) );
  AOI32X1 U672 ( .A0(n17126), .A1(n1309), .A2(n17008), .B0(n5327), .B1(n2903), 
        .Y(n17125) );
  OAI222XL U673 ( .A0(n401), .A1(n57), .B0(n2893), .B1(n30), .C0(n17072), .C1(
        n1309), .Y(n17256) );
  AOI221X1 U674 ( .A0(n5380), .A1(n17017), .B0(n998), .B1(n1310), .C0(n17018), 
        .Y(n17016) );
  AOI32X1 U675 ( .A0(n15866), .A1(n1297), .A2(n15748), .B0(n5639), .B1(n3135), 
        .Y(n15865) );
  OAI222XL U676 ( .A0(n415), .A1(n71), .B0(n3134), .B1(n44), .C0(n15812), .C1(
        n1297), .Y(n15996) );
  AOI221X1 U677 ( .A0(n5692), .A1(n15757), .B0(n1054), .B1(n1298), .C0(n15758), 
        .Y(n15756) );
  AOI32X1 U678 ( .A0(n14606), .A1(n1285), .A2(n14488), .B0(n5951), .B1(n3376), 
        .Y(n14605) );
  OAI222XL U679 ( .A0(n411), .A1(n67), .B0(n3375), .B1(n40), .C0(n14552), .C1(
        n1285), .Y(n14736) );
  AOI221X1 U680 ( .A0(n6004), .A1(n14497), .B0(n1110), .B1(n1286), .C0(n14498), 
        .Y(n14496) );
  AOI32X1 U681 ( .A0(n16496), .A1(n1303), .A2(n16378), .B0(n5487), .B1(n3016), 
        .Y(n16495) );
  OAI222XL U682 ( .A0(n409), .A1(n65), .B0(n3015), .B1(n38), .C0(n16442), .C1(
        n1303), .Y(n16626) );
  AOI221X1 U683 ( .A0(n5540), .A1(n16387), .B0(n1026), .B1(n1304), .C0(n16388), 
        .Y(n16386) );
  AOI32X1 U684 ( .A0(n17756), .A1(n1315), .A2(n17638), .B0(n5165), .B1(n2773), 
        .Y(n17755) );
  OAI222XL U685 ( .A0(n413), .A1(n69), .B0(n2772), .B1(n42), .C0(n17702), .C1(
        n1315), .Y(n17886) );
  AOI221X1 U686 ( .A0(n5218), .A1(n17647), .B0(n970), .B1(n1316), .C0(n17648), 
        .Y(n17646) );
  AOI32X1 U687 ( .A0(n14921), .A1(n1288), .A2(n14803), .B0(n5875), .B1(n3326), 
        .Y(n14920) );
  OAI222XL U688 ( .A0(n416), .A1(n64), .B0(n3314), .B1(n37), .C0(n14867), .C1(
        n1288), .Y(n15051) );
  AOI221X1 U689 ( .A0(n5928), .A1(n14812), .B0(n1096), .B1(n1289), .C0(n14813), 
        .Y(n14811) );
  AOI32X1 U690 ( .A0(n17441), .A1(n1312), .A2(n17323), .B0(n5243), .B1(n2834), 
        .Y(n17440) );
  OAI222XL U691 ( .A0(n408), .A1(n72), .B0(n2833), .B1(n45), .C0(n17387), .C1(
        n1312), .Y(n17571) );
  AOI221X1 U692 ( .A0(n5296), .A1(n17332), .B0(n984), .B1(n1313), .C0(n17333), 
        .Y(n17331) );
  AOI32X1 U693 ( .A0(n16181), .A1(n1300), .A2(n16063), .B0(n5563), .B1(n3073), 
        .Y(n16180) );
  OAI222XL U694 ( .A0(n406), .A1(n68), .B0(n3072), .B1(n41), .C0(n16127), .C1(
        n1300), .Y(n16311) );
  AOI221X1 U695 ( .A0(n5616), .A1(n16072), .B0(n1040), .B1(n1301), .C0(n16073), 
        .Y(n16071) );
  AOI32X1 U696 ( .A0(n14291), .A1(n1282), .A2(n14173), .B0(n6027), .B1(n3442), 
        .Y(n14290) );
  OAI222XL U697 ( .A0(n407), .A1(n70), .B0(n3433), .B1(n43), .C0(n14237), .C1(
        n1282), .Y(n14421) );
  AOI221X1 U698 ( .A0(n6080), .A1(n14182), .B0(n1124), .B1(n1283), .C0(n14183), 
        .Y(n14181) );
  AOI32X1 U699 ( .A0(n18071), .A1(n1318), .A2(n17953), .B0(n5057), .B1(n2720), 
        .Y(n18070) );
  OAI222XL U700 ( .A0(n405), .A1(n66), .B0(n2711), .B1(n39), .C0(n18017), .C1(
        n1318), .Y(n18201) );
  AOI221X1 U701 ( .A0(n5110), .A1(n17962), .B0(n956), .B1(n1319), .C0(n17963), 
        .Y(n17961) );
  AOI32X1 U702 ( .A0(n15551), .A1(n1294), .A2(n15433), .B0(n5715), .B1(n3202), 
        .Y(n15550) );
  OAI222XL U703 ( .A0(n410), .A1(n61), .B0(n3192), .B1(n34), .C0(n15497), .C1(
        n1294), .Y(n15681) );
  AOI221X1 U704 ( .A0(n5768), .A1(n15442), .B0(n1068), .B1(n1295), .C0(n15443), 
        .Y(n15441) );
  AOI32X1 U705 ( .A0(n18701), .A1(n1324), .A2(n18583), .B0(n4857), .B1(n2590), 
        .Y(n18700) );
  OAI222XL U706 ( .A0(n412), .A1(n63), .B0(n2598), .B1(n35), .C0(n18647), .C1(
        n1324), .Y(n18831) );
  AOI221X1 U707 ( .A0(n4910), .A1(n18592), .B0(n928), .B1(n1325), .C0(n18593), 
        .Y(n18591) );
  AOI222X1 U708 ( .A0(n1197), .A1(n12908), .B0(n13072), .B1(n1710), .C0(n6885), 
        .C1(n672), .Y(n13071) );
  AOI211X1 U709 ( .A0(n1200), .A1(n12908), .B0(n12943), .C0(n6888), .Y(n13053)
         );
  CLKINVX3 U710 ( .A(n696), .Y(n12908) );
  AOI222X1 U711 ( .A0(n1188), .A1(n12593), .B0(n12757), .B1(n1739), .C0(n6839), 
        .C1(n671), .Y(n12756) );
  AOI211X1 U712 ( .A0(n1191), .A1(n12593), .B0(n12628), .C0(n6842), .Y(n12738)
         );
  CLKINVX3 U713 ( .A(n694), .Y(n12593) );
  AOI222X1 U714 ( .A0(n1157), .A1(n13538), .B0(n13702), .B1(n1651), .C0(n6592), 
        .C1(n669), .Y(n13701) );
  AOI211X1 U715 ( .A0(n1160), .A1(n13538), .B0(n13573), .C0(n6595), .Y(n13683)
         );
  CLKINVX3 U716 ( .A(n695), .Y(n13538) );
  NAND2X2 U717 ( .A(top_core_io_n495), .B(n302), .Y(n285) );
  NAND2X2 U718 ( .A(top_core_io_n528), .B(n86), .Y(n274) );
  AOI222X1 U719 ( .A0(n591), .A1(n1228), .B0(n1127), .B1(n1119), .C0(n1122), 
        .C1(n1130), .Y(n7505) );
  OAI222XL U720 ( .A0(n3425), .A1(n7268), .B0(n1228), .B1(n20), .C0(n1130), 
        .C1(n7260), .Y(n7366) );
  AOI222X1 U721 ( .A0(n589), .A1(n1252), .B0(n959), .B1(n951), .C0(n954), .C1(
        n962), .Y(n11009) );
  OAI222XL U722 ( .A0(n2705), .A1(n10772), .B0(n1252), .B1(n18), .C0(n962), 
        .C1(n10764), .Y(n10870) );
  AOI222X1 U723 ( .A0(n592), .A1(n1248), .B0(n987), .B1(n979), .C0(n982), .C1(
        n990), .Y(n10425) );
  OAI222XL U724 ( .A0(n2828), .A1(n10188), .B0(n1248), .B1(n21), .C0(n990), 
        .C1(n10180), .Y(n10286) );
  AOI222X1 U725 ( .A0(n588), .A1(n1234), .B0(n1085), .B1(n1077), .C0(n1080), 
        .C1(n1088), .Y(n8381) );
  OAI222XL U726 ( .A0(n3245), .A1(n8144), .B0(n1234), .B1(n17), .C0(n1088), 
        .C1(n8136), .Y(n8242) );
  AOI222X1 U727 ( .A0(n587), .A1(n1254), .B0(n945), .B1(n937), .C0(n940), .C1(
        n948), .Y(n11301) );
  OAI222XL U728 ( .A0(n2643), .A1(n11064), .B0(n1254), .B1(n16), .C0(n948), 
        .C1(n11056), .Y(n11162) );
  AOI222X1 U729 ( .A0(n585), .A1(n1328), .B0(n1143), .B1(n1135), .C0(n1139), 
        .C1(n1145), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n319) );
  OAI222XL U730 ( .A0(n3492), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n79), 
        .B0(n1328), .B1(n14), .C0(n1145), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n70), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n180) );
  AOI222X1 U731 ( .A0(n586), .A1(n1246), .B0(n1001), .B1(n993), .C0(n996), 
        .C1(n1004), .Y(n10133) );
  OAI222XL U732 ( .A0(n2885), .A1(n9896), .B0(n1246), .B1(n15), .C0(n1004), 
        .C1(n9888), .Y(n9994) );
  AOI222X1 U733 ( .A0(n599), .A1(n1238), .B0(n1057), .B1(n1049), .C0(n1052), 
        .C1(n1060), .Y(n8965) );
  OAI222XL U734 ( .A0(n3127), .A1(n8728), .B0(n1238), .B1(n28), .C0(n1060), 
        .C1(n8720), .Y(n8826) );
  AOI222X1 U735 ( .A0(n595), .A1(n1230), .B0(n1113), .B1(n1105), .C0(n1108), 
        .C1(n1116), .Y(n7797) );
  OAI222XL U736 ( .A0(n3368), .A1(n7560), .B0(n1230), .B1(n24), .C0(n1116), 
        .C1(n7552), .Y(n7658) );
  AOI222X1 U737 ( .A0(n593), .A1(n1242), .B0(n1029), .B1(n1021), .C0(n1024), 
        .C1(n1032), .Y(n9549) );
  OAI222XL U738 ( .A0(n3007), .A1(n9312), .B0(n1242), .B1(n22), .C0(n1032), 
        .C1(n9304), .Y(n9410) );
  AOI222X1 U739 ( .A0(n597), .A1(n1250), .B0(n973), .B1(n965), .C0(n968), .C1(
        n976), .Y(n10717) );
  OAI222XL U740 ( .A0(n2765), .A1(n10480), .B0(n1250), .B1(n26), .C0(n976), 
        .C1(n10472), .Y(n10578) );
  AOI222X1 U741 ( .A0(n598), .A1(n1244), .B0(n1015), .B1(n1007), .C0(n1010), 
        .C1(n1018), .Y(n9841) );
  OAI222XL U742 ( .A0(n2947), .A1(n9604), .B0(n1244), .B1(n27), .C0(n1018), 
        .C1(n9596), .Y(n9702) );
  AOI222X1 U743 ( .A0(n594), .A1(n1236), .B0(n1071), .B1(n1063), .C0(n1066), 
        .C1(n1074), .Y(n8673) );
  OAI222XL U744 ( .A0(n3185), .A1(n8436), .B0(n1236), .B1(n23), .C0(n1074), 
        .C1(n8428), .Y(n8534) );
  AOI222X1 U745 ( .A0(n600), .A1(n1232), .B0(n1099), .B1(n1091), .C0(n1094), 
        .C1(n1102), .Y(n8089) );
  OAI222XL U746 ( .A0(n3306), .A1(n7852), .B0(n1232), .B1(n29), .C0(n1102), 
        .C1(n7844), .Y(n7950) );
  AOI222X1 U747 ( .A0(n596), .A1(n1256), .B0(n931), .B1(n923), .C0(n926), .C1(
        n934), .Y(n11593) );
  OAI222XL U748 ( .A0(n2583), .A1(n11356), .B0(n1256), .B1(n25), .C0(n934), 
        .C1(n11348), .Y(n11454) );
  AOI222X1 U749 ( .A0(n590), .A1(n1240), .B0(n1043), .B1(n1035), .C0(n1038), 
        .C1(n1046), .Y(n9257) );
  OAI222XL U750 ( .A0(n3068), .A1(n9020), .B0(n1240), .B1(n19), .C0(n1046), 
        .C1(n9012), .Y(n9118) );
  OAI222XL U751 ( .A0(n11967), .A1(n83), .B0(n1176), .B1(n12168), .C0(n12094), 
        .C1(n11977), .Y(n12181) );
  AOI222X1 U752 ( .A0(n1156), .A1(n1262), .B0(n6569), .B1(n11977), .C0(n1153), 
        .C1(n12007), .Y(n12240) );
  OAI222XL U753 ( .A0(n188), .A1(n11962), .B0(n12032), .B1(n11977), .C0(n12033), .C1(n12034), .Y(n12029) );
  CLKINVX3 U754 ( .A(n615), .Y(n11977) );
  OAI222XL U755 ( .A0(n12283), .A1(n82), .B0(n1181), .B1(n12483), .C0(n12409), 
        .C1(n1264), .Y(n12496) );
  AOI222X1 U756 ( .A0(n1165), .A1(n1266), .B0(n6616), .B1(n1264), .C0(n1162), 
        .C1(n12322), .Y(n12555) );
  OAI222XL U757 ( .A0(n46), .A1(n12278), .B0(n12347), .B1(n1263), .C0(n12348), 
        .C1(n12349), .Y(n12344) );
  OAI222XL U758 ( .A0(top_core_KE_sb1_n76), .A1(n81), .B0(n1216), .B1(
        top_core_KE_sb1_n281), .C0(top_core_KE_sb1_n206), .C1(
        top_core_KE_sb1_n86), .Y(top_core_KE_sb1_n294) );
  AOI222X1 U759 ( .A0(n1196), .A1(n1331), .B0(n6863), .B1(top_core_KE_sb1_n86), 
        .C0(n1193), .C1(top_core_KE_sb1_n116), .Y(top_core_KE_sb1_n353) );
  OAI222XL U760 ( .A0(n186), .A1(top_core_KE_sb1_n71), .B0(
        top_core_KE_sb1_n143), .B1(top_core_KE_sb1_n86), .C0(
        top_core_KE_sb1_n144), .C1(top_core_KE_sb1_n145), .Y(
        top_core_KE_sb1_n139) );
  CLKINVX3 U761 ( .A(n614), .Y(top_core_KE_sb1_n86) );
  OAI222XL U762 ( .A0(n11651), .A1(n80), .B0(n1222), .B1(n11852), .C0(n11778), 
        .C1(n11661), .Y(n11865) );
  AOI222X1 U763 ( .A0(n1205), .A1(n1259), .B0(n6909), .B1(n11661), .C0(n1202), 
        .C1(n11691), .Y(n11924) );
  OAI222XL U764 ( .A0(n185), .A1(n11646), .B0(n11716), .B1(n11661), .C0(n11717), .C1(n11718), .Y(n11713) );
  CLKINVX3 U765 ( .A(n613), .Y(n11661) );
  AOI221X1 U766 ( .A0(n6556), .A1(n1273), .B0(n1152), .B1(n13223), .C0(n13239), 
        .Y(n13237) );
  AOI221X1 U767 ( .A0(n6851), .A1(n1267), .B0(n1192), .B1(n12593), .C0(n12609), 
        .Y(n12607) );
  AOI221X1 U768 ( .A0(n6897), .A1(n1270), .B0(n1201), .B1(n12908), .C0(n12924), 
        .Y(n12922) );
  AOI222X1 U769 ( .A0(n6598), .A1(n13597), .B0(n6602), .B1(n1655), .C0(n6587), 
        .C1(n1276), .Y(n13762) );
  CLKINVX3 U770 ( .A(n685), .Y(n13597) );
  NAND2X2 U771 ( .A(top_core_io_n506), .B(n302), .Y(n284) );
  NAND2X2 U772 ( .A(top_core_io_n200), .B(n86), .Y(n281) );
  AOI221X1 U773 ( .A0(n1091), .A1(n3303), .B0(n7862), .B1(n1232), .C0(n8011), 
        .Y(n8010) );
  NOR2X1 U774 ( .A(n7845), .B(n3318), .Y(n8011) );
  AOI221X1 U775 ( .A0(n1049), .A1(n3123), .B0(n8738), .B1(n1238), .C0(n8887), 
        .Y(n8886) );
  NOR2X1 U776 ( .A(n8721), .B(n3136), .Y(n8887) );
  AOI221X1 U777 ( .A0(n1007), .A1(n2943), .B0(n9614), .B1(n1244), .C0(n9763), 
        .Y(n9762) );
  NOR2X1 U778 ( .A(n9597), .B(n2966), .Y(n9763) );
  AOI221X1 U779 ( .A0(n965), .A1(n2761), .B0(n10490), .B1(n1250), .C0(n10639), 
        .Y(n10638) );
  NOR2X1 U780 ( .A(n10473), .B(n2777), .Y(n10639) );
  AOI221X1 U781 ( .A0(n923), .A1(n2579), .B0(n11366), .B1(n1256), .C0(n11515), 
        .Y(n11514) );
  NOR2X1 U782 ( .A(n11349), .B(n2597), .Y(n11515) );
  AOI221X1 U783 ( .A0(n1105), .A1(n3364), .B0(n7570), .B1(n1230), .C0(n7719), 
        .Y(n7718) );
  NOR2X1 U784 ( .A(n7553), .B(n3377), .Y(n7719) );
  AOI221X1 U785 ( .A0(n1063), .A1(n3181), .B0(n8446), .B1(n1236), .C0(n8595), 
        .Y(n8594) );
  NOR2X1 U786 ( .A(n8429), .B(n3204), .Y(n8595) );
  AOI221X1 U787 ( .A0(n1021), .A1(n3004), .B0(n9322), .B1(n1242), .C0(n9471), 
        .Y(n9470) );
  NOR2X1 U788 ( .A(n9305), .B(n3017), .Y(n9471) );
  AOI221X1 U789 ( .A0(n979), .A1(n2822), .B0(n10198), .B1(n1248), .C0(n10347), 
        .Y(n10346) );
  NOR2X1 U790 ( .A(n10181), .B(n2842), .Y(n10347) );
  AOI221X1 U791 ( .A0(n1035), .A1(n3062), .B0(n9030), .B1(n1240), .C0(n9179), 
        .Y(n9178) );
  NOR2X1 U792 ( .A(n9013), .B(n3080), .Y(n9179) );
  AOI221X1 U793 ( .A0(n1119), .A1(n3422), .B0(n7278), .B1(n1228), .C0(n7427), 
        .Y(n7426) );
  NOR2X1 U794 ( .A(n7261), .B(n3435), .Y(n7427) );
  AOI221X1 U795 ( .A0(n951), .A1(n2701), .B0(n10782), .B1(n1252), .C0(n10931), 
        .Y(n10930) );
  NOR2X1 U796 ( .A(n10765), .B(n2713), .Y(n10931) );
  AOI221X1 U797 ( .A0(n1077), .A1(n3242), .B0(n8154), .B1(n1234), .C0(n8303), 
        .Y(n8302) );
  NOR2X1 U798 ( .A(n8137), .B(n3265), .Y(n8303) );
  AOI221X1 U799 ( .A0(n937), .A1(n2640), .B0(n11074), .B1(n1254), .C0(n11223), 
        .Y(n11222) );
  NOR2X1 U800 ( .A(n11057), .B(n2658), .Y(n11223) );
  AOI221X1 U801 ( .A0(n993), .A1(n2882), .B0(n9906), .B1(n1246), .C0(n10055), 
        .Y(n10054) );
  NOR2X1 U802 ( .A(n9889), .B(n2905), .Y(n10055) );
  AOI32X1 U803 ( .A0(n13346), .A1(n1273), .A2(n13229), .B0(n6467), .B1(n1688), 
        .Y(n13345) );
  OAI222XL U804 ( .A0(n692), .A1(n3), .B0(n1688), .B1(n73), .C0(n187), .C1(
        n1273), .Y(n13476) );
  CLKINVX3 U805 ( .A(n602), .Y(n1273) );
  AOI32X1 U806 ( .A0(n13031), .A1(n1270), .A2(n12914), .B0(n6812), .B1(n1717), 
        .Y(n13030) );
  OAI222XL U807 ( .A0(n696), .A1(n5), .B0(n1717), .B1(n75), .C0(n191), .C1(
        n1270), .Y(n13161) );
  CLKINVX3 U808 ( .A(n604), .Y(n1270) );
  AOI32X1 U809 ( .A0(n12716), .A1(n1267), .A2(n12599), .B0(n6770), .B1(n1746), 
        .Y(n12715) );
  OAI222XL U810 ( .A0(n694), .A1(n4), .B0(n1746), .B1(n74), .C0(n189), .C1(
        n1267), .Y(n12846) );
  CLKINVX3 U811 ( .A(n603), .Y(n1267) );
  OAI222XL U812 ( .A0(n13857), .A1(n31), .B0(n1142), .B1(n14058), .C0(n13985), 
        .C1(n13867), .Y(n14071) );
  AOI222X1 U813 ( .A0(n1137), .A1(n13911), .B0(n6125), .B1(n13867), .C0(n1133), 
        .C1(n13897), .Y(n14130) );
  OAI222XL U814 ( .A0(n13922), .A1(n1280), .B0(n13923), .B1(n13867), .C0(
        n13924), .C1(n13925), .Y(n13919) );
  CLKINVX3 U815 ( .A(n385), .Y(n13867) );
  OAI222XL U816 ( .A0(n15747), .A1(n44), .B0(n1059), .B1(n15948), .C0(n15875), 
        .C1(n15757), .Y(n15961) );
  AOI222X1 U817 ( .A0(n1054), .A1(n15801), .B0(n5669), .B1(n15757), .C0(n1050), 
        .C1(n15787), .Y(n16020) );
  OAI222XL U818 ( .A0(n15812), .A1(n1298), .B0(n15813), .B1(n15757), .C0(
        n15814), .C1(n15815), .Y(n15809) );
  CLKINVX3 U819 ( .A(n399), .Y(n15757) );
  OAI222XL U820 ( .A0(n17637), .A1(n42), .B0(n975), .B1(n17838), .C0(n17765), 
        .C1(n17647), .Y(n17851) );
  AOI222X1 U821 ( .A0(n970), .A1(n17691), .B0(n5195), .B1(n17647), .C0(n966), 
        .C1(n17677), .Y(n17910) );
  OAI222XL U822 ( .A0(n17702), .A1(n1316), .B0(n17703), .B1(n17647), .C0(
        n17704), .C1(n17705), .Y(n17699) );
  CLKINVX3 U823 ( .A(n397), .Y(n17647) );
  OAI222XL U824 ( .A0(n14487), .A1(n40), .B0(n1115), .B1(n14688), .C0(n14615), 
        .C1(n14497), .Y(n14701) );
  AOI222X1 U825 ( .A0(n1110), .A1(n14541), .B0(n5981), .B1(n14497), .C0(n1106), 
        .C1(n14527), .Y(n14760) );
  OAI222XL U826 ( .A0(n14552), .A1(n1286), .B0(n14553), .B1(n14497), .C0(
        n14554), .C1(n14555), .Y(n14549) );
  CLKINVX3 U827 ( .A(n395), .Y(n14497) );
  OAI222XL U828 ( .A0(n16377), .A1(n38), .B0(n1031), .B1(n16578), .C0(n16505), 
        .C1(n16387), .Y(n16591) );
  AOI222X1 U829 ( .A0(n1026), .A1(n16431), .B0(n5517), .B1(n16387), .C0(n1022), 
        .C1(n16417), .Y(n16650) );
  OAI222XL U830 ( .A0(n16442), .A1(n1304), .B0(n16443), .B1(n16387), .C0(
        n16444), .C1(n16445), .Y(n16439) );
  CLKINVX3 U831 ( .A(n393), .Y(n16387) );
  OAI222XL U832 ( .A0(n16692), .A1(n36), .B0(n1017), .B1(n16893), .C0(n16820), 
        .C1(n16702), .Y(n16906) );
  AOI222X1 U833 ( .A0(n1012), .A1(n16746), .B0(n5441), .B1(n16702), .C0(n1008), 
        .C1(n16732), .Y(n16965) );
  OAI222XL U834 ( .A0(n16757), .A1(n1307), .B0(n16758), .B1(n16702), .C0(
        n16759), .C1(n16760), .Y(n16754) );
  CLKINVX3 U835 ( .A(n391), .Y(n16702) );
  OAI222XL U836 ( .A0(n15117), .A1(n33), .B0(n1087), .B1(n15318), .C0(n15245), 
        .C1(n15127), .Y(n15331) );
  AOI222X1 U837 ( .A0(n1082), .A1(n15171), .B0(n5829), .B1(n15127), .C0(n1078), 
        .C1(n15157), .Y(n15390) );
  OAI222XL U838 ( .A0(n15182), .A1(n1292), .B0(n15183), .B1(n15127), .C0(
        n15184), .C1(n15185), .Y(n15179) );
  CLKINVX3 U839 ( .A(n388), .Y(n15127) );
  OAI222XL U840 ( .A0(n18267), .A1(n32), .B0(n947), .B1(n18468), .C0(n18395), 
        .C1(n18277), .Y(n18481) );
  AOI222X1 U841 ( .A0(n942), .A1(n18321), .B0(n5003), .B1(n18277), .C0(n938), 
        .C1(n18307), .Y(n18540) );
  OAI222XL U842 ( .A0(n18332), .A1(n1322), .B0(n18333), .B1(n18277), .C0(
        n18334), .C1(n18335), .Y(n18329) );
  CLKINVX3 U843 ( .A(n387), .Y(n18277) );
  OAI222XL U844 ( .A0(n17007), .A1(n30), .B0(n1003), .B1(n17208), .C0(n17135), 
        .C1(n17017), .Y(n17221) );
  AOI222X1 U845 ( .A0(n998), .A1(n17061), .B0(n5357), .B1(n17017), .C0(n994), 
        .C1(n17047), .Y(n17280) );
  OAI222XL U846 ( .A0(n17072), .A1(n1310), .B0(n17073), .B1(n17017), .C0(
        n17074), .C1(n17075), .Y(n17069) );
  CLKINVX3 U847 ( .A(n386), .Y(n17017) );
  OAI222XL U848 ( .A0(n14172), .A1(n43), .B0(n1129), .B1(n14373), .C0(n14300), 
        .C1(n14182), .Y(n14386) );
  AOI222X1 U849 ( .A0(n1124), .A1(n14226), .B0(n6057), .B1(n14182), .C0(n1120), 
        .C1(n14212), .Y(n14445) );
  OAI222XL U850 ( .A0(n14237), .A1(n1283), .B0(n14238), .B1(n14182), .C0(
        n14239), .C1(n14240), .Y(n14234) );
  CLKINVX3 U851 ( .A(n398), .Y(n14182) );
  OAI222XL U852 ( .A0(n17952), .A1(n39), .B0(n961), .B1(n18153), .C0(n18080), 
        .C1(n17962), .Y(n18166) );
  AOI222X1 U853 ( .A0(n956), .A1(n18006), .B0(n5087), .B1(n17962), .C0(n952), 
        .C1(n17992), .Y(n18225) );
  OAI222XL U854 ( .A0(n18017), .A1(n1319), .B0(n18018), .B1(n17962), .C0(
        n18019), .C1(n18020), .Y(n18014) );
  CLKINVX3 U855 ( .A(n394), .Y(n17962) );
  OAI222XL U856 ( .A0(n15432), .A1(n34), .B0(n1073), .B1(n15633), .C0(n15560), 
        .C1(n15442), .Y(n15646) );
  AOI222X1 U857 ( .A0(n1068), .A1(n15486), .B0(n5745), .B1(n15442), .C0(n1064), 
        .C1(n15472), .Y(n15705) );
  OAI222XL U858 ( .A0(n15497), .A1(n1295), .B0(n15498), .B1(n15442), .C0(
        n15499), .C1(n15500), .Y(n15494) );
  CLKINVX3 U859 ( .A(n389), .Y(n15442) );
  OAI222XL U860 ( .A0(n17322), .A1(n45), .B0(n989), .B1(n17523), .C0(n17450), 
        .C1(n17332), .Y(n17536) );
  AOI222X1 U861 ( .A0(n984), .A1(n17376), .B0(n5273), .B1(n17332), .C0(n980), 
        .C1(n17362), .Y(n17595) );
  OAI222XL U862 ( .A0(n17387), .A1(n1313), .B0(n17388), .B1(n17332), .C0(
        n17389), .C1(n17390), .Y(n17384) );
  CLKINVX3 U863 ( .A(n400), .Y(n17332) );
  OAI222XL U864 ( .A0(n16062), .A1(n41), .B0(n1045), .B1(n16263), .C0(n16190), 
        .C1(n16072), .Y(n16276) );
  AOI222X1 U865 ( .A0(n1040), .A1(n16116), .B0(n5593), .B1(n16072), .C0(n1036), 
        .C1(n16102), .Y(n16335) );
  OAI222XL U866 ( .A0(n16127), .A1(n1301), .B0(n16128), .B1(n16072), .C0(
        n16129), .C1(n16130), .Y(n16124) );
  CLKINVX3 U867 ( .A(n396), .Y(n16072) );
  OAI222XL U868 ( .A0(n18582), .A1(n35), .B0(n933), .B1(n18783), .C0(n18710), 
        .C1(n18592), .Y(n18796) );
  AOI222X1 U869 ( .A0(n928), .A1(n18636), .B0(n4887), .B1(n18592), .C0(n924), 
        .C1(n18622), .Y(n18855) );
  OAI222XL U870 ( .A0(n18647), .A1(n1325), .B0(n18648), .B1(n18592), .C0(
        n18649), .C1(n18650), .Y(n18644) );
  CLKINVX3 U871 ( .A(n390), .Y(n18592) );
  OAI222XL U872 ( .A0(n14802), .A1(n37), .B0(n1101), .B1(n15003), .C0(n14930), 
        .C1(n14812), .Y(n15016) );
  AOI222X1 U873 ( .A0(n1096), .A1(n14856), .B0(n5905), .B1(n14812), .C0(n1092), 
        .C1(n14842), .Y(n15075) );
  OAI222XL U874 ( .A0(n14867), .A1(n1289), .B0(n14868), .B1(n14812), .C0(
        n14869), .C1(n14870), .Y(n14864) );
  CLKINVX3 U875 ( .A(n392), .Y(n14812) );
  CLKINVX3 U876 ( .A(n601), .Y(n1264) );
  AOI222X1 U877 ( .A0(n6550), .A1(n13282), .B0(n6554), .B1(n1686), .C0(n6539), 
        .C1(n1273), .Y(n13447) );
  OAI222XL U878 ( .A0(n13295), .A1(n13282), .B0(n1681), .B1(n13293), .C0(n1367), .C1(n13312), .Y(n13308) );
  CLKINVX3 U879 ( .A(n686), .Y(n13282) );
  AOI222X1 U880 ( .A0(n5675), .A1(n15801), .B0(n5690), .B1(n3132), .C0(n5665), 
        .C1(n1297), .Y(n15967) );
  OAI222XL U881 ( .A0(n15815), .A1(n15801), .B0(n3123), .B1(n15813), .C0(n3108), .C1(n15832), .Y(n15828) );
  CLKINVX3 U882 ( .A(n527), .Y(n15801) );
  AOI222X1 U883 ( .A0(n5201), .A1(n17691), .B0(n5216), .B1(n2770), .C0(n5191), 
        .C1(n1315), .Y(n17857) );
  OAI222XL U884 ( .A0(n17705), .A1(n17691), .B0(n2761), .B1(n17703), .C0(n2746), .C1(n17722), .Y(n17718) );
  CLKINVX3 U885 ( .A(n525), .Y(n17691) );
  AOI222X1 U886 ( .A0(n5987), .A1(n14541), .B0(n6002), .B1(n3373), .C0(n5977), 
        .C1(n1285), .Y(n14707) );
  OAI222XL U887 ( .A0(n14555), .A1(n14541), .B0(n3364), .B1(n14553), .C0(n3349), .C1(n14572), .Y(n14568) );
  CLKINVX3 U888 ( .A(n523), .Y(n14541) );
  AOI222X1 U889 ( .A0(n5523), .A1(n16431), .B0(n5538), .B1(n3012), .C0(n5513), 
        .C1(n1303), .Y(n16597) );
  OAI222XL U890 ( .A0(n16445), .A1(n16431), .B0(n3004), .B1(n16443), .C0(n2989), .C1(n16462), .Y(n16458) );
  CLKINVX3 U891 ( .A(n521), .Y(n16431) );
  AOI222X1 U892 ( .A0(n5447), .A1(n16746), .B0(n5462), .B1(n2951), .C0(n5437), 
        .C1(n1306), .Y(n16912) );
  OAI222XL U893 ( .A0(n16760), .A1(n16746), .B0(n2943), .B1(n16758), .C0(n2928), .C1(n16777), .Y(n16773) );
  CLKINVX3 U894 ( .A(n519), .Y(n16746) );
  AOI222X1 U895 ( .A0(n5835), .A1(n15171), .B0(n5850), .B1(n3250), .C0(n5825), 
        .C1(n1291), .Y(n15337) );
  OAI222XL U896 ( .A0(n15185), .A1(n15171), .B0(n3242), .B1(n15183), .C0(n3227), .C1(n15202), .Y(n15198) );
  CLKINVX3 U897 ( .A(n516), .Y(n15171) );
  AOI222X1 U898 ( .A0(n5009), .A1(n18321), .B0(n5024), .B1(n2648), .C0(n4999), 
        .C1(n1321), .Y(n18487) );
  OAI222XL U899 ( .A0(n18335), .A1(n18321), .B0(n2640), .B1(n18333), .C0(n2625), .C1(n18352), .Y(n18348) );
  CLKINVX3 U900 ( .A(n515), .Y(n18321) );
  AOI222X1 U901 ( .A0(n6131), .A1(n13911), .B0(n6149), .B1(n3489), .C0(n6121), 
        .C1(n1279), .Y(n14077) );
  OAI222XL U902 ( .A0(n13925), .A1(n13911), .B0(n3483), .B1(n13923), .C0(n3468), .C1(n13942), .Y(n13938) );
  CLKINVX3 U903 ( .A(n514), .Y(n13911) );
  AOI222X1 U904 ( .A0(n5363), .A1(n17061), .B0(n5378), .B1(n2890), .C0(n5353), 
        .C1(n1309), .Y(n17227) );
  OAI222XL U905 ( .A0(n17075), .A1(n17061), .B0(n2882), .B1(n17073), .C0(n2867), .C1(n17092), .Y(n17088) );
  CLKINVX3 U906 ( .A(n513), .Y(n17061) );
  AOI222X1 U907 ( .A0(n6063), .A1(n14226), .B0(n6078), .B1(n3430), .C0(n6053), 
        .C1(n1282), .Y(n14392) );
  OAI222XL U908 ( .A0(n14240), .A1(n14226), .B0(n3422), .B1(n14238), .C0(n3407), .C1(n14257), .Y(n14253) );
  CLKINVX3 U909 ( .A(n526), .Y(n14226) );
  AOI222X1 U910 ( .A0(n5093), .A1(n18006), .B0(n5108), .B1(n2709), .C0(n5083), 
        .C1(n1318), .Y(n18172) );
  OAI222XL U911 ( .A0(n18020), .A1(n18006), .B0(n2701), .B1(n18018), .C0(n2686), .C1(n18037), .Y(n18033) );
  CLKINVX3 U912 ( .A(n522), .Y(n18006) );
  AOI222X1 U913 ( .A0(n5751), .A1(n15486), .B0(n5766), .B1(n3190), .C0(n5741), 
        .C1(n1294), .Y(n15652) );
  OAI222XL U914 ( .A0(n15500), .A1(n15486), .B0(n3181), .B1(n15498), .C0(n3166), .C1(n15517), .Y(n15513) );
  CLKINVX3 U915 ( .A(n517), .Y(n15486) );
  AOI222X1 U916 ( .A0(n5279), .A1(n17376), .B0(n5294), .B1(n2830), .C0(n5269), 
        .C1(n1312), .Y(n17542) );
  OAI222XL U917 ( .A0(n17390), .A1(n17376), .B0(n2822), .B1(n17388), .C0(n2807), .C1(n17407), .Y(n17403) );
  CLKINVX3 U918 ( .A(n528), .Y(n17376) );
  AOI222X1 U919 ( .A0(n5599), .A1(n16116), .B0(n5614), .B1(n3070), .C0(n5589), 
        .C1(n1300), .Y(n16282) );
  OAI222XL U920 ( .A0(n16130), .A1(n16116), .B0(n3062), .B1(n16128), .C0(n3047), .C1(n16147), .Y(n16143) );
  CLKINVX3 U921 ( .A(n524), .Y(n16116) );
  AOI222X1 U922 ( .A0(n5911), .A1(n14856), .B0(n5926), .B1(n3311), .C0(n5901), 
        .C1(n1288), .Y(n15022) );
  OAI222XL U923 ( .A0(n14870), .A1(n14856), .B0(n3303), .B1(n14868), .C0(n3288), .C1(n14887), .Y(n14883) );
  CLKINVX3 U924 ( .A(n520), .Y(n14856) );
  AOI222X1 U925 ( .A0(n4893), .A1(n18636), .B0(n4908), .B1(n2588), .C0(n4883), 
        .C1(n1324), .Y(n18802) );
  OAI222XL U926 ( .A0(n18650), .A1(n18636), .B0(n2579), .B1(n18648), .C0(n2564), .C1(n18667), .Y(n18663) );
  CLKINVX3 U927 ( .A(n518), .Y(n18636) );
  AOI222X1 U928 ( .A0(n6845), .A1(n12652), .B0(n6849), .B1(n1744), .C0(n6834), 
        .C1(n1267), .Y(n12817) );
  CLKINVX3 U929 ( .A(n688), .Y(n12652) );
  AOI222X1 U930 ( .A0(n6891), .A1(n12967), .B0(n6895), .B1(n1715), .C0(n6880), 
        .C1(n1270), .Y(n13132) );
  CLKINVX3 U931 ( .A(n687), .Y(n12967) );
  NAND2X2 U932 ( .A(top_core_io_n517), .B(n302), .Y(n283) );
  NAND2X2 U933 ( .A(top_core_io_n211), .B(n86), .Y(n280) );
  NAND2X2 U934 ( .A(n304), .B(top_core_io_n60), .Y(n290) );
  NOR2X1 U935 ( .A(n7844), .B(n7926), .Y(n7968) );
  NOR2X1 U936 ( .A(n8720), .B(n8802), .Y(n8844) );
  NOR2X1 U937 ( .A(n9596), .B(n9678), .Y(n9720) );
  NOR2X1 U938 ( .A(n10472), .B(n10554), .Y(n10596) );
  NOR2X1 U939 ( .A(n11348), .B(n11430), .Y(n11472) );
  NOR2X1 U940 ( .A(n7552), .B(n7634), .Y(n7676) );
  NOR2X1 U941 ( .A(n8428), .B(n8510), .Y(n8552) );
  NOR2X1 U942 ( .A(n9304), .B(n9386), .Y(n9428) );
  NOR2X1 U943 ( .A(n10180), .B(n10262), .Y(n10304) );
  NOR2X1 U944 ( .A(n9012), .B(n9094), .Y(n9136) );
  NOR2X1 U945 ( .A(n7260), .B(n7342), .Y(n7384) );
  NOR2X1 U946 ( .A(n10764), .B(n10846), .Y(n10888) );
  NOR2X1 U947 ( .A(n8136), .B(n8218), .Y(n8260) );
  NOR2X1 U948 ( .A(n11056), .B(n11138), .Y(n11180) );
  NOR2X1 U949 ( .A(n9888), .B(n9970), .Y(n10012) );
  NOR2X1 U950 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n70), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n198) );
  AOI222X1 U951 ( .A0(n1172), .A1(n6556), .B0(n13238), .B1(n13240), .C0(n13268), .C1(n6539), .Y(n13265) );
  OAI222XL U952 ( .A0(n13228), .A1(n73), .B0(n1173), .B1(n13428), .C0(n13355), 
        .C1(n13238), .Y(n13441) );
  AOI222X1 U953 ( .A0(n1152), .A1(n1275), .B0(n6544), .B1(n13238), .C0(n1148), 
        .C1(n13268), .Y(n13500) );
  OAI222XL U954 ( .A0(n187), .A1(n13223), .B0(n13293), .B1(n13238), .C0(n13294), .C1(n13295), .Y(n13290) );
  CLKINVX3 U955 ( .A(n610), .Y(n13238) );
  OAI221XL U956 ( .A0(n7284), .A1(n1228), .B0(n7285), .B1(n7286), .C0(n7287), 
        .Y(n7283) );
  AOI221X1 U957 ( .A0(n7278), .A1(n3440), .B0(n1119), .B1(n1228), .C0(n6037), 
        .Y(n7269) );
  OAI221XL U958 ( .A0(n7291), .A1(n7285), .B0(n7404), .B1(n1228), .C0(n7460), 
        .Y(n7458) );
  CLKINVX3 U959 ( .A(n535), .Y(n1228) );
  OAI221XL U960 ( .A0(n7868), .A1(n1232), .B0(n7869), .B1(n7870), .C0(n7871), 
        .Y(n7867) );
  AOI221X1 U961 ( .A0(n7862), .A1(n3322), .B0(n1091), .B1(n1232), .C0(n5885), 
        .Y(n7853) );
  OAI221XL U962 ( .A0(n7875), .A1(n7869), .B0(n7988), .B1(n1232), .C0(n8044), 
        .Y(n8042) );
  CLKINVX3 U963 ( .A(n544), .Y(n1232) );
  OAI221XL U964 ( .A0(n11372), .A1(n1256), .B0(n11373), .B1(n11374), .C0(
        n11375), .Y(n11371) );
  AOI221X1 U965 ( .A0(n11366), .A1(n2591), .B0(n923), .B1(n1256), .C0(n4867), 
        .Y(n11357) );
  OAI221XL U966 ( .A0(n11379), .A1(n11373), .B0(n11492), .B1(n1256), .C0(
        n11548), .Y(n11546) );
  CLKINVX3 U967 ( .A(n540), .Y(n1256) );
  OAI221XL U968 ( .A0(n10204), .A1(n1248), .B0(n10205), .B1(n10206), .C0(
        n10207), .Y(n10203) );
  AOI221X1 U969 ( .A0(n10198), .A1(n2839), .B0(n979), .B1(n1248), .C0(n5253), 
        .Y(n10189) );
  OAI221XL U970 ( .A0(n10211), .A1(n10205), .B0(n10324), .B1(n1248), .C0(
        n10380), .Y(n10378) );
  CLKINVX3 U971 ( .A(n536), .Y(n1248) );
  OAI221XL U972 ( .A0(n9620), .A1(n1244), .B0(n9621), .B1(n9622), .C0(n9623), 
        .Y(n9619) );
  AOI221X1 U973 ( .A0(n9614), .A1(n2956), .B0(n1007), .B1(n1244), .C0(n5421), 
        .Y(n9605) );
  OAI221XL U974 ( .A0(n9627), .A1(n9621), .B0(n9740), .B1(n1244), .C0(n9796), 
        .Y(n9794) );
  CLKINVX3 U975 ( .A(n542), .Y(n1244) );
  OAI221XL U976 ( .A0(n8452), .A1(n1236), .B0(n8453), .B1(n8454), .C0(n8455), 
        .Y(n8451) );
  AOI221X1 U977 ( .A0(n8446), .A1(n3194), .B0(n1063), .B1(n1236), .C0(n5725), 
        .Y(n8437) );
  OAI221XL U978 ( .A0(n8459), .A1(n8453), .B0(n8572), .B1(n1236), .C0(n8628), 
        .Y(n8626) );
  CLKINVX3 U979 ( .A(n538), .Y(n1236) );
  OAI221XL U980 ( .A0(n9036), .A1(n1240), .B0(n9037), .B1(n9038), .C0(n9039), 
        .Y(n9035) );
  AOI221X1 U981 ( .A0(n9030), .A1(n3074), .B0(n1035), .B1(n1240), .C0(n5573), 
        .Y(n9021) );
  OAI221XL U982 ( .A0(n9043), .A1(n9037), .B0(n9156), .B1(n1240), .C0(n9212), 
        .Y(n9210) );
  CLKINVX3 U983 ( .A(n534), .Y(n1240) );
  OAI221XL U984 ( .A0(n10788), .A1(n1252), .B0(n10789), .B1(n10790), .C0(
        n10791), .Y(n10787) );
  AOI221X1 U985 ( .A0(n10782), .A1(n2718), .B0(n951), .B1(n1252), .C0(n5067), 
        .Y(n10773) );
  OAI221XL U986 ( .A0(n10795), .A1(n10789), .B0(n10908), .B1(n1252), .C0(
        n10964), .Y(n10962) );
  CLKINVX3 U987 ( .A(n533), .Y(n1252) );
  OAI221XL U988 ( .A0(n8160), .A1(n1234), .B0(n8161), .B1(n8162), .C0(n8163), 
        .Y(n8159) );
  AOI221X1 U989 ( .A0(n8154), .A1(n3255), .B0(n1077), .B1(n1234), .C0(n5809), 
        .Y(n8145) );
  OAI221XL U990 ( .A0(n8167), .A1(n8161), .B0(n8280), .B1(n1234), .C0(n8336), 
        .Y(n8334) );
  CLKINVX3 U991 ( .A(n532), .Y(n1234) );
  OAI221XL U992 ( .A0(n11080), .A1(n1254), .B0(n11081), .B1(n11082), .C0(
        n11083), .Y(n11079) );
  AOI221X1 U993 ( .A0(n11074), .A1(n2652), .B0(n937), .B1(n1254), .C0(n4983), 
        .Y(n11065) );
  OAI221XL U994 ( .A0(n11087), .A1(n11081), .B0(n11200), .B1(n1254), .C0(
        n11256), .Y(n11254) );
  CLKINVX3 U995 ( .A(n531), .Y(n1254) );
  OAI221XL U996 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n96), .A1(n1328), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n98), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n99), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n95) );
  AOI221X1 U997 ( .A0(n1135), .A1(n3483), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n89), .B1(n1328), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n241), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n240) );
  AOI221X1 U998 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n89), .A1(n3502), 
        .B0(n1135), .B1(n1328), .C0(n6133), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n80) );
  OAI221XL U999 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n104), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n218), .B1(n1328), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n274), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n272) );
  CLKINVX3 U1000 ( .A(n530), .Y(n1328) );
  OAI221XL U1001 ( .A0(n9912), .A1(n1246), .B0(n9913), .B1(n9914), .C0(n9915), 
        .Y(n9911) );
  AOI221X1 U1002 ( .A0(n9906), .A1(n2895), .B0(n993), .B1(n1246), .C0(n5337), 
        .Y(n9897) );
  OAI221XL U1003 ( .A0(n9919), .A1(n9913), .B0(n10032), .B1(n1246), .C0(n10088), .Y(n10086) );
  CLKINVX3 U1004 ( .A(n529), .Y(n1246) );
  OAI221XL U1005 ( .A0(n8744), .A1(n1238), .B0(n8745), .B1(n8746), .C0(n8747), 
        .Y(n8743) );
  AOI221X1 U1006 ( .A0(n8738), .A1(n3142), .B0(n1049), .B1(n1238), .C0(n5649), 
        .Y(n8729) );
  OAI221XL U1007 ( .A0(n8751), .A1(n8745), .B0(n8864), .B1(n1238), .C0(n8920), 
        .Y(n8918) );
  CLKINVX3 U1008 ( .A(n543), .Y(n1238) );
  OAI221XL U1009 ( .A0(n7576), .A1(n1230), .B0(n7577), .B1(n7578), .C0(n7579), 
        .Y(n7575) );
  AOI221X1 U1010 ( .A0(n7570), .A1(n3383), .B0(n1105), .B1(n1230), .C0(n5961), 
        .Y(n7561) );
  OAI221XL U1011 ( .A0(n7583), .A1(n7577), .B0(n7696), .B1(n1230), .C0(n7752), 
        .Y(n7750) );
  CLKINVX3 U1012 ( .A(n539), .Y(n1230) );
  OAI221XL U1013 ( .A0(n9328), .A1(n1242), .B0(n9329), .B1(n9330), .C0(n9331), 
        .Y(n9327) );
  AOI221X1 U1014 ( .A0(n9322), .A1(n3023), .B0(n1021), .B1(n1242), .C0(n5497), 
        .Y(n9313) );
  OAI221XL U1015 ( .A0(n9335), .A1(n9329), .B0(n9448), .B1(n1242), .C0(n9504), 
        .Y(n9502) );
  CLKINVX3 U1016 ( .A(n537), .Y(n1242) );
  OAI221XL U1017 ( .A0(n10496), .A1(n1250), .B0(n10497), .B1(n10498), .C0(
        n10499), .Y(n10495) );
  AOI221X1 U1018 ( .A0(n10490), .A1(n2778), .B0(n965), .B1(n1250), .C0(n5175), 
        .Y(n10481) );
  OAI221XL U1019 ( .A0(n10503), .A1(n10497), .B0(n10616), .B1(n1250), .C0(
        n10672), .Y(n10670) );
  CLKINVX3 U1020 ( .A(n541), .Y(n1250) );
  AOI222X1 U1021 ( .A0(n13294), .A1(n748), .B0(n1148), .B1(n610), .C0(n1152), 
        .C1(n1274), .Y(n13406) );
  AOI222X1 U1022 ( .A0(n1667), .A1(n13498), .B0(n6467), .B1(n1274), .C0(n6470), 
        .C1(n13268), .Y(n13497) );
  AOI222X1 U1023 ( .A0(n6539), .A1(n1275), .B0(n6556), .B1(n1274), .C0(n6544), 
        .C1(n1173), .Y(n13413) );
  OAI221XL U1024 ( .A0(n1691), .A1(n13293), .B0(n180), .B1(n1274), .C0(n13429), 
        .Y(n13416) );
  CLKINVX3 U1025 ( .A(n677), .Y(n1274) );
  AOI222X1 U1026 ( .A0(n12979), .A1(n750), .B0(n1197), .B1(n612), .C0(n1201), 
        .C1(n1271), .Y(n13091) );
  AOI222X1 U1027 ( .A0(n1696), .A1(n13183), .B0(n6812), .B1(n1271), .C0(n6813), 
        .C1(n12953), .Y(n13182) );
  AOI222X1 U1028 ( .A0(n6880), .A1(n1272), .B0(n6897), .B1(n1271), .C0(n6885), 
        .C1(n1219), .Y(n13098) );
  OAI221XL U1029 ( .A0(n1720), .A1(n12978), .B0(n182), .B1(n1271), .C0(n13114), 
        .Y(n13101) );
  CLKINVX3 U1030 ( .A(n680), .Y(n1271) );
  AOI222X1 U1031 ( .A0(n12664), .A1(n749), .B0(n1188), .B1(n611), .C0(n1192), 
        .C1(n1268), .Y(n12776) );
  AOI222X1 U1032 ( .A0(n1725), .A1(n12868), .B0(n6770), .B1(n1268), .C0(n6773), 
        .C1(n12638), .Y(n12867) );
  AOI222X1 U1033 ( .A0(n6834), .A1(n1269), .B0(n6851), .B1(n1268), .C0(n6839), 
        .C1(n1213), .Y(n12783) );
  OAI221XL U1034 ( .A0(n1749), .A1(n12663), .B0(n181), .B1(n1268), .C0(n12799), 
        .Y(n12786) );
  CLKINVX3 U1035 ( .A(n678), .Y(n1268) );
  AOI222X1 U1036 ( .A0(n13609), .A1(n751), .B0(n1157), .B1(n616), .C0(n1161), 
        .C1(n1277), .Y(n13721) );
  AOI222X1 U1037 ( .A0(n6587), .A1(n1278), .B0(n6604), .B1(n1277), .C0(n6592), 
        .C1(n1178), .Y(n13728) );
  OAI221XL U1038 ( .A0(n1663), .A1(n13608), .B0(n183), .B1(n1277), .C0(n13744), 
        .Y(n13731) );
  CLKINVX3 U1039 ( .A(n679), .Y(n1277) );
  AOI222X1 U1040 ( .A0(n6564), .A1(n1262), .B0(n6580), .B1(n1261), .C0(n6569), 
        .C1(n1176), .Y(n12153) );
  OAI221XL U1041 ( .A0(n1791), .A1(n12032), .B0(n79), .B1(n1261), .C0(n12169), 
        .Y(n12156) );
  CLKINVX3 U1042 ( .A(n676), .Y(n1261) );
  AOI222X1 U1043 ( .A0(n6904), .A1(n1259), .B0(n6920), .B1(n1258), .C0(n6909), 
        .C1(n1222), .Y(n11837) );
  OAI221XL U1044 ( .A0(n1812), .A1(n11716), .B0(n77), .B1(n1258), .C0(n11853), 
        .Y(n11840) );
  CLKINVX3 U1045 ( .A(n673), .Y(n1258) );
  AOI222X1 U1046 ( .A0(n6858), .A1(n1331), .B0(n6874), .B1(n1330), .C0(n6863), 
        .C1(n1216), .Y(top_core_KE_sb1_n266) );
  OAI221XL U1047 ( .A0(n1833), .A1(top_core_KE_sb1_n143), .B0(n78), .B1(n1330), 
        .C0(top_core_KE_sb1_n282), .Y(top_core_KE_sb1_n269) );
  CLKINVX3 U1048 ( .A(n674), .Y(n1330) );
  AOI222X1 U1049 ( .A0(n6611), .A1(n1266), .B0(n6627), .B1(n1265), .C0(n6616), 
        .C1(n1181), .Y(n12468) );
  OAI221XL U1050 ( .A0(n1770), .A1(n12347), .B0(n184), .B1(n1265), .C0(n12484), 
        .Y(n12471) );
  CLKINVX3 U1051 ( .A(n675), .Y(n1265) );
  OAI32X1 U1052 ( .A0(n15866), .A1(n3119), .A2(n15747), .B0(n1299), .B1(n15902), .Y(n15901) );
  AOI221X1 U1053 ( .A0(n5674), .A1(n1299), .B0(n1050), .B1(n1298), .C0(n15913), 
        .Y(n16036) );
  CLKINVX3 U1054 ( .A(n463), .Y(n1299) );
  OAI32X1 U1055 ( .A0(n17756), .A1(n2757), .A2(n17637), .B0(n1317), .B1(n17792), .Y(n17791) );
  AOI221X1 U1056 ( .A0(n5200), .A1(n1317), .B0(n966), .B1(n1316), .C0(n17803), 
        .Y(n17926) );
  CLKINVX3 U1057 ( .A(n461), .Y(n1317) );
  OAI32X1 U1058 ( .A0(n14606), .A1(n3360), .A2(n14487), .B0(n1287), .B1(n14642), .Y(n14641) );
  AOI221X1 U1059 ( .A0(n5986), .A1(n1287), .B0(n1106), .B1(n1286), .C0(n14653), 
        .Y(n14776) );
  CLKINVX3 U1060 ( .A(n459), .Y(n1287) );
  OAI32X1 U1061 ( .A0(n16496), .A1(n3000), .A2(n16377), .B0(n1305), .B1(n16532), .Y(n16531) );
  AOI221X1 U1062 ( .A0(n5522), .A1(n1305), .B0(n1022), .B1(n1304), .C0(n16543), 
        .Y(n16666) );
  CLKINVX3 U1063 ( .A(n457), .Y(n1305) );
  OAI32X1 U1064 ( .A0(n16811), .A1(n2939), .A2(n16692), .B0(n1308), .B1(n16847), .Y(n16846) );
  AOI221X1 U1065 ( .A0(n5446), .A1(n1308), .B0(n1008), .B1(n1307), .C0(n16858), 
        .Y(n16981) );
  CLKINVX3 U1066 ( .A(n455), .Y(n1308) );
  OAI32X1 U1067 ( .A0(n15236), .A1(n3238), .A2(n15117), .B0(n1293), .B1(n15272), .Y(n15271) );
  AOI221X1 U1068 ( .A0(n5834), .A1(n1293), .B0(n1078), .B1(n1292), .C0(n15283), 
        .Y(n15406) );
  CLKINVX3 U1069 ( .A(n452), .Y(n1293) );
  OAI32X1 U1070 ( .A0(n18386), .A1(n2636), .A2(n18267), .B0(n1323), .B1(n18422), .Y(n18421) );
  AOI221X1 U1071 ( .A0(n5008), .A1(n1323), .B0(n938), .B1(n1322), .C0(n18433), 
        .Y(n18556) );
  CLKINVX3 U1072 ( .A(n451), .Y(n1323) );
  OAI32X1 U1073 ( .A0(n17126), .A1(n2878), .A2(n17007), .B0(n1311), .B1(n17162), .Y(n17161) );
  AOI221X1 U1074 ( .A0(n5362), .A1(n1311), .B0(n994), .B1(n1310), .C0(n17173), 
        .Y(n17296) );
  CLKINVX3 U1075 ( .A(n450), .Y(n1311) );
  OAI32X1 U1076 ( .A0(n13976), .A1(n3478), .A2(n13857), .B0(n1281), .B1(n14012), .Y(n14011) );
  AOI221X1 U1077 ( .A0(n6130), .A1(n1281), .B0(n1133), .B1(n1280), .C0(n14023), 
        .Y(n14146) );
  CLKINVX3 U1078 ( .A(n449), .Y(n1281) );
  OAI32X1 U1079 ( .A0(n14921), .A1(n3299), .A2(n14802), .B0(n1290), .B1(n14957), .Y(n14956) );
  AOI221X1 U1080 ( .A0(n5910), .A1(n1290), .B0(n1092), .B1(n1289), .C0(n14968), 
        .Y(n15091) );
  CLKINVX3 U1081 ( .A(n456), .Y(n1290) );
  OAI32X1 U1082 ( .A0(n18701), .A1(n2575), .A2(n18582), .B0(n1326), .B1(n18737), .Y(n18736) );
  AOI221X1 U1083 ( .A0(n4892), .A1(n1326), .B0(n924), .B1(n1325), .C0(n18748), 
        .Y(n18871) );
  CLKINVX3 U1084 ( .A(n454), .Y(n1326) );
  OAI32X1 U1085 ( .A0(n17441), .A1(n2818), .A2(n17322), .B0(n1314), .B1(n17477), .Y(n17476) );
  AOI221X1 U1086 ( .A0(n5278), .A1(n1314), .B0(n980), .B1(n1313), .C0(n17488), 
        .Y(n17611) );
  CLKINVX3 U1087 ( .A(n464), .Y(n1314) );
  OAI32X1 U1088 ( .A0(n16181), .A1(n3058), .A2(n16062), .B0(n1302), .B1(n16217), .Y(n16216) );
  AOI221X1 U1089 ( .A0(n5598), .A1(n1302), .B0(n1036), .B1(n1301), .C0(n16228), 
        .Y(n16351) );
  CLKINVX3 U1090 ( .A(n460), .Y(n1302) );
  OAI32X1 U1091 ( .A0(n15551), .A1(n3177), .A2(n15432), .B0(n1296), .B1(n15587), .Y(n15586) );
  AOI221X1 U1092 ( .A0(n5750), .A1(n1296), .B0(n1064), .B1(n1295), .C0(n15598), 
        .Y(n15721) );
  CLKINVX3 U1093 ( .A(n453), .Y(n1296) );
  OAI32X1 U1094 ( .A0(n14291), .A1(n3418), .A2(n14172), .B0(n1284), .B1(n14327), .Y(n14326) );
  AOI221X1 U1095 ( .A0(n6062), .A1(n1284), .B0(n1120), .B1(n1283), .C0(n14338), 
        .Y(n14461) );
  CLKINVX3 U1096 ( .A(n462), .Y(n1284) );
  OAI32X1 U1097 ( .A0(n18071), .A1(n2697), .A2(n17952), .B0(n1320), .B1(n18107), .Y(n18106) );
  AOI221X1 U1098 ( .A0(n5092), .A1(n1320), .B0(n952), .B1(n1319), .C0(n18118), 
        .Y(n18241) );
  CLKINVX3 U1099 ( .A(n458), .Y(n1320) );
  OAI222XL U1100 ( .A0(n691), .A1(n12410), .B0(n1768), .B1(n82), .C0(n46), 
        .C1(n1263), .Y(n12531) );
  OAI222XL U1101 ( .A0(n689), .A1(n11779), .B0(n1810), .B1(n80), .C0(n185), 
        .C1(n1257), .Y(n11900) );
  OAI222XL U1102 ( .A0(n690), .A1(top_core_KE_sb1_n207), .B0(n1831), .B1(n81), 
        .C0(n186), .C1(n1329), .Y(top_core_KE_sb1_n329) );
  OAI222XL U1103 ( .A0(n693), .A1(n12095), .B0(n1789), .B1(n83), .C0(n188), 
        .C1(n1260), .Y(n12216) );
  CLKINVX3 U1104 ( .A(n727), .Y(n16757) );
  CLKINVX3 U1105 ( .A(n725), .Y(n15182) );
  CLKINVX3 U1106 ( .A(n724), .Y(n18332) );
  CLKINVX3 U1107 ( .A(n723), .Y(n13922) );
  CLKINVX3 U1108 ( .A(n722), .Y(n17072) );
  CLKINVX3 U1109 ( .A(n736), .Y(n15812) );
  CLKINVX3 U1110 ( .A(n732), .Y(n14552) );
  CLKINVX3 U1111 ( .A(n730), .Y(n16442) );
  CLKINVX3 U1112 ( .A(n734), .Y(n17702) );
  CLKINVX3 U1113 ( .A(n735), .Y(n14237) );
  CLKINVX3 U1114 ( .A(n731), .Y(n18017) );
  CLKINVX3 U1115 ( .A(n726), .Y(n15497) );
  CLKINVX3 U1116 ( .A(n737), .Y(n17387) );
  CLKINVX3 U1117 ( .A(n733), .Y(n16127) );
  CLKINVX3 U1118 ( .A(n729), .Y(n14867) );
  CLKINVX3 U1119 ( .A(n728), .Y(n18647) );
  NAND2X2 U1120 ( .A(top_core_io_n528), .B(n302), .Y(n282) );
  NAND2X2 U1121 ( .A(top_core_io_n222), .B(n86), .Y(n279) );
  NAND2X2 U1122 ( .A(top_core_io_n233), .B(n303), .Y(n271) );
  NAND2X2 U1123 ( .A(n304), .B(top_core_io_n27), .Y(n293) );
  AOI211X1 U1124 ( .A0(n150), .A1(n1102), .B0(n5891), .C0(n7951), .Y(n8072) );
  NOR2X1 U1125 ( .A(n7845), .B(n440), .Y(n7951) );
  AOI211X1 U1126 ( .A0(n149), .A1(n1060), .B0(n5655), .C0(n8827), .Y(n8948) );
  NOR2X1 U1127 ( .A(n8721), .B(n447), .Y(n8827) );
  AOI211X1 U1128 ( .A0(n148), .A1(n1018), .B0(n5427), .C0(n9703), .Y(n9824) );
  NOR2X1 U1129 ( .A(n9597), .B(n438), .Y(n9703) );
  AOI211X1 U1130 ( .A0(n147), .A1(n976), .B0(n5181), .C0(n10579), .Y(n10700)
         );
  NOR2X1 U1131 ( .A(n10473), .B(n445), .Y(n10579) );
  AOI211X1 U1132 ( .A0(n146), .A1(n934), .B0(n4873), .C0(n11455), .Y(n11576)
         );
  NOR2X1 U1133 ( .A(n11349), .B(n439), .Y(n11455) );
  AOI211X1 U1134 ( .A0(n145), .A1(n1116), .B0(n5967), .C0(n7659), .Y(n7780) );
  NOR2X1 U1135 ( .A(n7553), .B(n443), .Y(n7659) );
  AOI211X1 U1136 ( .A0(n144), .A1(n1074), .B0(n5731), .C0(n8535), .Y(n8656) );
  NOR2X1 U1137 ( .A(n8429), .B(n437), .Y(n8535) );
  AOI211X1 U1138 ( .A0(n143), .A1(n1032), .B0(n5503), .C0(n9411), .Y(n9532) );
  NOR2X1 U1139 ( .A(n9305), .B(n441), .Y(n9411) );
  AOI211X1 U1140 ( .A0(n142), .A1(n990), .B0(n5259), .C0(n10287), .Y(n10408)
         );
  NOR2X1 U1141 ( .A(n10181), .B(n448), .Y(n10287) );
  AOI211X1 U1142 ( .A0(n140), .A1(n1046), .B0(n5579), .C0(n9119), .Y(n9240) );
  NOR2X1 U1143 ( .A(n9013), .B(n444), .Y(n9119) );
  AOI211X1 U1144 ( .A0(n141), .A1(n1130), .B0(n6043), .C0(n7367), .Y(n7488) );
  NOR2X1 U1145 ( .A(n7261), .B(n446), .Y(n7367) );
  AOI211X1 U1146 ( .A0(n139), .A1(n962), .B0(n5073), .C0(n10871), .Y(n10992)
         );
  NOR2X1 U1147 ( .A(n10765), .B(n442), .Y(n10871) );
  AOI211X1 U1148 ( .A0(n138), .A1(n1088), .B0(n5815), .C0(n8243), .Y(n8364) );
  NOR2X1 U1149 ( .A(n8137), .B(n436), .Y(n8243) );
  AOI211X1 U1150 ( .A0(n137), .A1(n948), .B0(n4989), .C0(n11163), .Y(n11284)
         );
  NOR2X1 U1151 ( .A(n11057), .B(n435), .Y(n11163) );
  AOI211X1 U1152 ( .A0(n136), .A1(n1145), .B0(n6139), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n181), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n302) );
  NOR2X1 U1153 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n71), .B(n434), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n181) );
  AOI211X1 U1154 ( .A0(n135), .A1(n1004), .B0(n5343), .C0(n9995), .Y(n10116)
         );
  NOR2X1 U1155 ( .A(n9889), .B(n433), .Y(n9995) );
  NAND2X1 U1156 ( .A(n1094), .B(n7856), .Y(n7912) );
  NAND2X1 U1157 ( .A(n1052), .B(n8732), .Y(n8788) );
  NAND2X1 U1158 ( .A(n1010), .B(n9608), .Y(n9664) );
  NAND2X1 U1159 ( .A(n968), .B(n10484), .Y(n10540) );
  NAND2X1 U1160 ( .A(n926), .B(n11360), .Y(n11416) );
  NAND2X1 U1161 ( .A(n1108), .B(n7564), .Y(n7620) );
  NAND2X1 U1162 ( .A(n1066), .B(n8440), .Y(n8496) );
  NAND2X1 U1163 ( .A(n1024), .B(n9316), .Y(n9372) );
  NAND2X1 U1164 ( .A(n982), .B(n10192), .Y(n10248) );
  NAND2X1 U1165 ( .A(n1122), .B(n7272), .Y(n7328) );
  NAND2X1 U1166 ( .A(n1038), .B(n9024), .Y(n9080) );
  NAND2X1 U1167 ( .A(n954), .B(n10776), .Y(n10832) );
  NAND2X1 U1168 ( .A(n1080), .B(n8148), .Y(n8204) );
  NAND2X1 U1169 ( .A(n940), .B(n11068), .Y(n11124) );
  NAND2X1 U1170 ( .A(n1139), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n141) );
  NAND2X1 U1171 ( .A(n996), .B(n9900), .Y(n9956) );
  AOI222X1 U1172 ( .A0(n1218), .A1(n6897), .B0(n12923), .B1(n12925), .C0(
        n12953), .C1(n6880), .Y(n12950) );
  OAI222XL U1173 ( .A0(n12913), .A1(n75), .B0(n1219), .B1(n13113), .C0(n13040), 
        .C1(n12923), .Y(n13126) );
  AOI222X1 U1174 ( .A0(n1201), .A1(n1272), .B0(n6885), .B1(n12923), .C0(n1197), 
        .C1(n12953), .Y(n13185) );
  CLKINVX3 U1175 ( .A(n612), .Y(n12923) );
  AOI222X1 U1176 ( .A0(n1212), .A1(n6851), .B0(n12608), .B1(n12610), .C0(
        n12638), .C1(n6834), .Y(n12635) );
  OAI222XL U1177 ( .A0(n12598), .A1(n74), .B0(n1213), .B1(n12798), .C0(n12725), 
        .C1(n12608), .Y(n12811) );
  AOI222X1 U1178 ( .A0(n1192), .A1(n1269), .B0(n6839), .B1(n12608), .C0(n1188), 
        .C1(n12638), .Y(n12870) );
  CLKINVX3 U1179 ( .A(n611), .Y(n12608) );
  CLKINVX3 U1180 ( .A(n384), .Y(n1312) );
  CLKINVX3 U1181 ( .A(n382), .Y(n1282) );
  CLKINVX3 U1182 ( .A(n380), .Y(n1300) );
  CLKINVX3 U1183 ( .A(n378), .Y(n1318) );
  CLKINVX3 U1184 ( .A(n376), .Y(n1288) );
  CLKINVX3 U1185 ( .A(n375), .Y(n1306) );
  CLKINVX3 U1186 ( .A(n374), .Y(n1324) );
  CLKINVX3 U1187 ( .A(n373), .Y(n1294) );
  CLKINVX3 U1188 ( .A(n372), .Y(n1291) );
  CLKINVX3 U1189 ( .A(n371), .Y(n1321) );
  CLKINVX3 U1190 ( .A(n370), .Y(n1309) );
  CLKINVX3 U1191 ( .A(n369), .Y(n1279) );
  CLKINVX3 U1192 ( .A(n383), .Y(n1297) );
  CLKINVX3 U1193 ( .A(n379), .Y(n1285) );
  CLKINVX3 U1194 ( .A(n377), .Y(n1303) );
  CLKINVX3 U1195 ( .A(n381), .Y(n1315) );
  OAI32X1 U1196 ( .A0(n12085), .A1(n1359), .A2(n11967), .B0(n12021), .B1(
        n12122), .Y(n12121) );
  AOI221X1 U1197 ( .A0(n6574), .A1(n12021), .B0(n1153), .B1(n11962), .C0(
        n12133), .Y(n12256) );
  OAI32X1 U1198 ( .A0(n12400), .A1(n1358), .A2(n12283), .B0(n12336), .B1(
        n12437), .Y(n12436) );
  AOI221X1 U1199 ( .A0(n6621), .A1(n12336), .B0(n1162), .B1(n12278), .C0(
        n12448), .Y(n12571) );
  OAI32X1 U1200 ( .A0(top_core_KE_sb1_n197), .A1(n1345), .A2(
        top_core_KE_sb1_n76), .B0(top_core_KE_sb1_n130), .B1(
        top_core_KE_sb1_n234), .Y(top_core_KE_sb1_n233) );
  AOI221X1 U1201 ( .A0(n6868), .A1(top_core_KE_sb1_n130), .B0(n1193), .B1(
        top_core_KE_sb1_n71), .C0(top_core_KE_sb1_n245), .Y(
        top_core_KE_sb1_n370) );
  OAI32X1 U1202 ( .A0(n11769), .A1(n1344), .A2(n11651), .B0(n11705), .B1(
        n11806), .Y(n11805) );
  AOI221X1 U1203 ( .A0(n6914), .A1(n11705), .B0(n1202), .B1(n11646), .C0(
        n11817), .Y(n11940) );
  OAI32X1 U1204 ( .A0(n13031), .A1(n1703), .A2(n12913), .B0(n12967), .B1(
        n13067), .Y(n13066) );
  OAI32X1 U1205 ( .A0(n12716), .A1(n1732), .A2(n12598), .B0(n12652), .B1(
        n12752), .Y(n12751) );
  OAI32X1 U1206 ( .A0(n13346), .A1(n1674), .A2(n13228), .B0(n1275), .B1(n13382), .Y(n13381) );
  AOI221X1 U1207 ( .A0(n6549), .A1(n13282), .B0(n1148), .B1(n13223), .C0(
        n13393), .Y(n13516) );
  OAI32X1 U1208 ( .A0(n13661), .A1(top_core_KE_prev_key1_reg_90_), .A2(n13543), 
        .B0(n13597), .B1(n13697), .Y(n13696) );
  AOI222X1 U1209 ( .A0(n5437), .A1(n1308), .B0(n5464), .B1(n1307), .C0(n5441), 
        .C1(n1017), .Y(n16878) );
  AOI222X1 U1210 ( .A0(n5825), .A1(n1293), .B0(n5852), .B1(n1292), .C0(n5829), 
        .C1(n1087), .Y(n15303) );
  AOI222X1 U1211 ( .A0(n4999), .A1(n1323), .B0(n5026), .B1(n1322), .C0(n5003), 
        .C1(n947), .Y(n18453) );
  AOI222X1 U1212 ( .A0(n6121), .A1(n1281), .B0(n6151), .B1(n1280), .C0(n6125), 
        .C1(n1142), .Y(n14043) );
  AOI222X1 U1213 ( .A0(n5353), .A1(n1311), .B0(n5380), .B1(n1310), .C0(n5357), 
        .C1(n1003), .Y(n17193) );
  AOI222X1 U1214 ( .A0(n5665), .A1(n1299), .B0(n5692), .B1(n1298), .C0(n5669), 
        .C1(n1059), .Y(n15933) );
  AOI222X1 U1215 ( .A0(n5977), .A1(n1287), .B0(n6004), .B1(n1286), .C0(n5981), 
        .C1(n1115), .Y(n14673) );
  AOI222X1 U1216 ( .A0(n5513), .A1(n1305), .B0(n5540), .B1(n1304), .C0(n5517), 
        .C1(n1031), .Y(n16563) );
  AOI222X1 U1217 ( .A0(n5191), .A1(n1317), .B0(n5218), .B1(n1316), .C0(n5195), 
        .C1(n975), .Y(n17823) );
  AOI222X1 U1218 ( .A0(n6053), .A1(n1284), .B0(n6080), .B1(n1283), .C0(n6057), 
        .C1(n1129), .Y(n14358) );
  AOI222X1 U1219 ( .A0(n5083), .A1(n1320), .B0(n5110), .B1(n1319), .C0(n5087), 
        .C1(n961), .Y(n18138) );
  AOI222X1 U1220 ( .A0(n5741), .A1(n1296), .B0(n5768), .B1(n1295), .C0(n5745), 
        .C1(n1073), .Y(n15618) );
  AOI222X1 U1221 ( .A0(n5269), .A1(n1314), .B0(n5296), .B1(n1313), .C0(n5273), 
        .C1(n989), .Y(n17508) );
  AOI222X1 U1222 ( .A0(n5589), .A1(n1302), .B0(n5616), .B1(n1301), .C0(n5593), 
        .C1(n1045), .Y(n16248) );
  AOI222X1 U1223 ( .A0(n5901), .A1(n1290), .B0(n5928), .B1(n1289), .C0(n5905), 
        .C1(n1101), .Y(n14988) );
  AOI222X1 U1224 ( .A0(n4883), .A1(n1326), .B0(n4910), .B1(n1325), .C0(n4887), 
        .C1(n933), .Y(n18768) );
  OAI221XL U1225 ( .A0(n675), .A1(n89), .B0(n12349), .B1(n1771), .C0(n12530), 
        .Y(n12525) );
  CLKINVX3 U1226 ( .A(n760), .Y(n12349) );
  OAI221XL U1227 ( .A0(n676), .A1(n53), .B0(n12034), .B1(n1790), .C0(n12215), 
        .Y(n12210) );
  CLKINVX3 U1228 ( .A(n763), .Y(n12034) );
  OAI221XL U1229 ( .A0(n674), .A1(n51), .B0(top_core_KE_sb1_n145), .B1(n1832), 
        .C0(top_core_KE_sb1_n328), .Y(top_core_KE_sb1_n323) );
  CLKINVX3 U1230 ( .A(n762), .Y(top_core_KE_sb1_n145) );
  OAI221XL U1231 ( .A0(n673), .A1(n50), .B0(n11718), .B1(n1811), .C0(n11899), 
        .Y(n11894) );
  CLKINVX3 U1232 ( .A(n761), .Y(n11718) );
  CLKINVX3 U1233 ( .A(n703), .Y(n16760) );
  CLKINVX3 U1234 ( .A(n699), .Y(n13925) );
  CLKINVX3 U1235 ( .A(n701), .Y(n15185) );
  CLKINVX3 U1236 ( .A(n700), .Y(n18335) );
  CLKINVX3 U1237 ( .A(n698), .Y(n17075) );
  CLKINVX3 U1238 ( .A(n712), .Y(n15815) );
  CLKINVX3 U1239 ( .A(n708), .Y(n14555) );
  CLKINVX3 U1240 ( .A(n706), .Y(n16445) );
  CLKINVX3 U1241 ( .A(n710), .Y(n17705) );
  CLKINVX3 U1242 ( .A(n702), .Y(n15500) );
  CLKINVX3 U1243 ( .A(n711), .Y(n14240) );
  CLKINVX3 U1244 ( .A(n707), .Y(n18020) );
  CLKINVX3 U1245 ( .A(n713), .Y(n17390) );
  CLKINVX3 U1246 ( .A(n709), .Y(n16130) );
  CLKINVX3 U1247 ( .A(n705), .Y(n14870) );
  CLKINVX3 U1248 ( .A(n704), .Y(n18650) );
  NAND2X2 U1249 ( .A(top_core_io_n233), .B(n86), .Y(n278) );
  NAND2X2 U1250 ( .A(n86), .B(top_core_io_n27), .Y(n297) );
  NAND2X2 U1251 ( .A(top_core_io_n200), .B(n302), .Y(n289) );
  NAND2X2 U1252 ( .A(top_core_io_n528), .B(n303), .Y(n267) );
  NAND2X2 U1253 ( .A(n304), .B(top_core_io_n38), .Y(n292) );
  NOR2X1 U1254 ( .A(n8728), .B(n367), .Y(n8867) );
  NOR2X1 U1255 ( .A(n10480), .B(n365), .Y(n10619) );
  NOR2X1 U1256 ( .A(n7560), .B(n363), .Y(n7699) );
  NOR2X1 U1257 ( .A(n9312), .B(n361), .Y(n9451) );
  NOR2X1 U1258 ( .A(n7268), .B(n358), .Y(n7407) );
  NOR2X1 U1259 ( .A(n8144), .B(n355), .Y(n8283) );
  NOR2X1 U1260 ( .A(n11064), .B(n356), .Y(n11203) );
  NOR2X1 U1261 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .B(n354), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n221) );
  NOR2X1 U1262 ( .A(n9896), .B(n353), .Y(n10035) );
  NOR2X1 U1263 ( .A(n10772), .B(n357), .Y(n10911) );
  NOR2X1 U1264 ( .A(n10188), .B(n360), .Y(n10327) );
  NOR2X1 U1265 ( .A(n9604), .B(n366), .Y(n9743) );
  NOR2X1 U1266 ( .A(n8436), .B(n362), .Y(n8575) );
  NOR2X1 U1267 ( .A(n7852), .B(n368), .Y(n7991) );
  NOR2X1 U1268 ( .A(n11356), .B(n364), .Y(n11495) );
  NOR2X1 U1269 ( .A(n9020), .B(n359), .Y(n9159) );
  AOI211X1 U1270 ( .A0(n150), .A1(n504), .B0(n7883), .C0(n8000), .Y(n8094) );
  NOR2X1 U1271 ( .A(n105), .B(n456), .Y(n8000) );
  AOI211X1 U1272 ( .A0(n149), .A1(n511), .B0(n8759), .C0(n8876), .Y(n8970) );
  NOR2X1 U1273 ( .A(n104), .B(n463), .Y(n8876) );
  AOI211X1 U1274 ( .A0(n148), .A1(n503), .B0(n9635), .C0(n9752), .Y(n9846) );
  NOR2X1 U1275 ( .A(n103), .B(n455), .Y(n9752) );
  AOI211X1 U1276 ( .A0(n147), .A1(n509), .B0(n10511), .C0(n10628), .Y(n10722)
         );
  NOR2X1 U1277 ( .A(n102), .B(n461), .Y(n10628) );
  AOI211X1 U1278 ( .A0(n146), .A1(n502), .B0(n11387), .C0(n11504), .Y(n11598)
         );
  NOR2X1 U1279 ( .A(n101), .B(n454), .Y(n11504) );
  AOI211X1 U1280 ( .A0(n145), .A1(n507), .B0(n7591), .C0(n7708), .Y(n7802) );
  NOR2X1 U1281 ( .A(n100), .B(n459), .Y(n7708) );
  AOI211X1 U1282 ( .A0(n144), .A1(n499), .B0(n8467), .C0(n8584), .Y(n8678) );
  NOR2X1 U1283 ( .A(n99), .B(n453), .Y(n8584) );
  AOI211X1 U1284 ( .A0(n143), .A1(n505), .B0(n9343), .C0(n9460), .Y(n9554) );
  NOR2X1 U1285 ( .A(n98), .B(n457), .Y(n9460) );
  AOI211X1 U1286 ( .A0(n142), .A1(n512), .B0(n10219), .C0(n10336), .Y(n10430)
         );
  NOR2X1 U1287 ( .A(n97), .B(n464), .Y(n10336) );
  AOI211X1 U1288 ( .A0(n141), .A1(n510), .B0(n7299), .C0(n7416), .Y(n7510) );
  NOR2X1 U1289 ( .A(n95), .B(n462), .Y(n7416) );
  AOI211X1 U1290 ( .A0(n140), .A1(n508), .B0(n9051), .C0(n9168), .Y(n9262) );
  NOR2X1 U1291 ( .A(n96), .B(n460), .Y(n9168) );
  AOI211X1 U1292 ( .A0(n139), .A1(n506), .B0(n10803), .C0(n10920), .Y(n11014)
         );
  NOR2X1 U1293 ( .A(n94), .B(n458), .Y(n10920) );
  AOI211X1 U1294 ( .A0(n138), .A1(n500), .B0(n8175), .C0(n8292), .Y(n8386) );
  NOR2X1 U1295 ( .A(n93), .B(n452), .Y(n8292) );
  AOI211X1 U1296 ( .A0(n137), .A1(n501), .B0(n11095), .C0(n11212), .Y(n11306)
         );
  NOR2X1 U1297 ( .A(n92), .B(n451), .Y(n11212) );
  AOI211X1 U1298 ( .A0(n136), .A1(n497), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n112), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n230), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n324) );
  NOR2X1 U1299 ( .A(n91), .B(n449), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n230) );
  AOI211X1 U1300 ( .A0(n135), .A1(n498), .B0(n9927), .C0(n10044), .Y(n10138)
         );
  NOR2X1 U1301 ( .A(n90), .B(n450), .Y(n10044) );
  NOR2XL U1302 ( .A(n12095), .B(n581), .Y(n240) );
  CLKINVX3 U1303 ( .A(n747), .Y(n12095) );
  NOR2XL U1304 ( .A(n12410), .B(n579), .Y(n241) );
  CLKINVX3 U1305 ( .A(n744), .Y(n12410) );
  NOR2XL U1306 ( .A(top_core_KE_sb1_n207), .B(n578), .Y(n242) );
  CLKINVX3 U1307 ( .A(n746), .Y(top_core_KE_sb1_n207) );
  NOR2XL U1308 ( .A(n11779), .B(n577), .Y(n243) );
  CLKINVX3 U1309 ( .A(n745), .Y(n11779) );
  NOR2XL U1310 ( .A(n72), .B(n352), .Y(n244) );
  NOR2XL U1311 ( .A(n71), .B(n351), .Y(n245) );
  NOR2XL U1312 ( .A(n70), .B(n350), .Y(n246) );
  NOR2XL U1313 ( .A(n69), .B(n349), .Y(n247) );
  NOR2XL U1314 ( .A(n68), .B(n348), .Y(n248) );
  NOR2XL U1315 ( .A(n67), .B(n347), .Y(n249) );
  NOR2XL U1316 ( .A(n66), .B(n346), .Y(n250) );
  NOR2XL U1317 ( .A(n65), .B(n345), .Y(n251) );
  NOR2XL U1318 ( .A(n64), .B(n344), .Y(n252) );
  NOR2XL U1319 ( .A(n63), .B(n343), .Y(n253) );
  NOR2XL U1320 ( .A(n62), .B(n342), .Y(n254) );
  NOR2XL U1321 ( .A(n61), .B(n341), .Y(n255) );
  NOR2XL U1322 ( .A(n60), .B(n340), .Y(n256) );
  NOR2XL U1323 ( .A(n59), .B(n339), .Y(n257) );
  NOR2XL U1324 ( .A(n58), .B(n338), .Y(n258) );
  NOR2XL U1325 ( .A(n57), .B(n337), .Y(n259) );
  NAND2X1 U1326 ( .A(n1161), .B(n13543), .Y(n13561) );
  NAND2X1 U1327 ( .A(n1152), .B(n13228), .Y(n13246) );
  NAND2X1 U1328 ( .A(n1192), .B(n12598), .Y(n12616) );
  NAND2X1 U1329 ( .A(n1201), .B(n12913), .Y(n12931) );
  AOI32X1 U1330 ( .A0(n12085), .A1(n1260), .A2(n11968), .B0(n6502), .B1(n1789), 
        .Y(n12084) );
  AOI221X1 U1331 ( .A0(n6580), .A1(n1260), .B0(n1156), .B1(n11962), .C0(n11978), .Y(n11976) );
  CLKINVX3 U1332 ( .A(n608), .Y(n1260) );
  AOI32X1 U1333 ( .A0(top_core_KE_sb1_n197), .A1(n1329), .A2(
        top_core_KE_sb1_n77), .B0(n6799), .B1(n1831), .Y(top_core_KE_sb1_n196)
         );
  AOI221X1 U1334 ( .A0(n6874), .A1(n1329), .B0(n1196), .B1(top_core_KE_sb1_n71), .C0(top_core_KE_sb1_n87), .Y(top_core_KE_sb1_n85) );
  CLKINVX3 U1335 ( .A(n606), .Y(n1329) );
  AOI32X1 U1336 ( .A0(n11769), .A1(n1257), .A2(n11652), .B0(n6823), .B1(n1810), 
        .Y(n11768) );
  AOI221X1 U1337 ( .A0(n6920), .A1(n1257), .B0(n1205), .B1(n11646), .C0(n11662), .Y(n11660) );
  CLKINVX3 U1338 ( .A(n605), .Y(n1257) );
  AOI32X1 U1339 ( .A0(n12400), .A1(n1263), .A2(n12284), .B0(n6527), .B1(n1768), 
        .Y(n12399) );
  AOI221X1 U1340 ( .A0(n6627), .A1(n1263), .B0(n1165), .B1(n12278), .C0(n12293), .Y(n12292) );
  CLKINVX3 U1341 ( .A(n607), .Y(n1263) );
  AOI211X1 U1342 ( .A0(n747), .A1(n11962), .B0(n11997), .C0(n6572), .Y(n12108)
         );
  CLKINVX3 U1343 ( .A(n693), .Y(n11962) );
  AOI211X1 U1344 ( .A0(n744), .A1(n12278), .B0(n12312), .C0(n6619), .Y(n12423)
         );
  CLKINVX3 U1345 ( .A(n691), .Y(n12278) );
  AOI211X1 U1346 ( .A0(n746), .A1(top_core_KE_sb1_n71), .B0(
        top_core_KE_sb1_n106), .C0(n6866), .Y(top_core_KE_sb1_n220) );
  CLKINVX3 U1347 ( .A(n690), .Y(top_core_KE_sb1_n71) );
  AOI211X1 U1348 ( .A0(n745), .A1(n11646), .B0(n11681), .C0(n6912), .Y(n11792)
         );
  CLKINVX3 U1349 ( .A(n689), .Y(n11646) );
  OAI221XL U1350 ( .A0(n2958), .A1(n16758), .B0(n170), .B1(n1307), .C0(n16894), 
        .Y(n16881) );
  CLKINVX3 U1351 ( .A(n470), .Y(n1307) );
  OAI221XL U1352 ( .A0(n2840), .A1(n17388), .B0(n179), .B1(n1313), .C0(n17524), 
        .Y(n17511) );
  CLKINVX3 U1353 ( .A(n480), .Y(n1313) );
  OAI221XL U1354 ( .A0(n3076), .A1(n16128), .B0(n175), .B1(n1301), .C0(n16264), 
        .Y(n16251) );
  CLKINVX3 U1355 ( .A(n476), .Y(n1301) );
  OAI221XL U1356 ( .A0(n3320), .A1(n14868), .B0(n171), .B1(n1289), .C0(n15004), 
        .Y(n14991) );
  CLKINVX3 U1357 ( .A(n472), .Y(n1289) );
  OAI221XL U1358 ( .A0(n3437), .A1(n14238), .B0(n177), .B1(n1283), .C0(n14374), 
        .Y(n14361) );
  CLKINVX3 U1359 ( .A(n478), .Y(n1283) );
  OAI221XL U1360 ( .A0(n2715), .A1(n18018), .B0(n173), .B1(n1319), .C0(n18154), 
        .Y(n18141) );
  CLKINVX3 U1361 ( .A(n474), .Y(n1319) );
  OAI221XL U1362 ( .A0(n3196), .A1(n15498), .B0(n168), .B1(n1295), .C0(n15634), 
        .Y(n15621) );
  CLKINVX3 U1363 ( .A(n469), .Y(n1295) );
  OAI221XL U1364 ( .A0(n3257), .A1(n15183), .B0(n167), .B1(n1292), .C0(n15319), 
        .Y(n15306) );
  CLKINVX3 U1365 ( .A(n468), .Y(n1292) );
  OAI221XL U1366 ( .A0(n2654), .A1(n18333), .B0(n166), .B1(n1322), .C0(n18469), 
        .Y(n18456) );
  CLKINVX3 U1367 ( .A(n467), .Y(n1322) );
  OAI221XL U1368 ( .A0(n3498), .A1(n13923), .B0(n165), .B1(n1280), .C0(n14059), 
        .Y(n14046) );
  CLKINVX3 U1369 ( .A(n466), .Y(n1280) );
  OAI221XL U1370 ( .A0(n2897), .A1(n17073), .B0(n164), .B1(n1310), .C0(n17209), 
        .Y(n17196) );
  CLKINVX3 U1371 ( .A(n465), .Y(n1310) );
  OAI221XL U1372 ( .A0(n3140), .A1(n15813), .B0(n178), .B1(n1298), .C0(n15949), 
        .Y(n15936) );
  CLKINVX3 U1373 ( .A(n479), .Y(n1298) );
  OAI221XL U1374 ( .A0(n3381), .A1(n14553), .B0(n174), .B1(n1286), .C0(n14689), 
        .Y(n14676) );
  CLKINVX3 U1375 ( .A(n475), .Y(n1286) );
  OAI221XL U1376 ( .A0(n3021), .A1(n16443), .B0(n172), .B1(n1304), .C0(n16579), 
        .Y(n16566) );
  CLKINVX3 U1377 ( .A(n473), .Y(n1304) );
  OAI221XL U1378 ( .A0(n2780), .A1(n17703), .B0(n176), .B1(n1316), .C0(n17839), 
        .Y(n17826) );
  CLKINVX3 U1379 ( .A(n477), .Y(n1316) );
  OAI221XL U1380 ( .A0(n2593), .A1(n18648), .B0(n169), .B1(n1325), .C0(n18784), 
        .Y(n18771) );
  CLKINVX3 U1381 ( .A(n471), .Y(n1325) );
  CLKINVX3 U1382 ( .A(n496), .Y(n1231) );
  CLKINVX3 U1383 ( .A(n495), .Y(n1237) );
  CLKINVX3 U1384 ( .A(n494), .Y(n1243) );
  CLKINVX3 U1385 ( .A(n493), .Y(n1249) );
  CLKINVX3 U1386 ( .A(n492), .Y(n1255) );
  CLKINVX3 U1387 ( .A(n491), .Y(n1229) );
  CLKINVX3 U1388 ( .A(n490), .Y(n1235) );
  CLKINVX3 U1389 ( .A(n489), .Y(n1241) );
  CLKINVX3 U1390 ( .A(n488), .Y(n1247) );
  CLKINVX3 U1391 ( .A(n487), .Y(n1227) );
  CLKINVX3 U1392 ( .A(n486), .Y(n1239) );
  CLKINVX3 U1393 ( .A(n485), .Y(n1251) );
  CLKINVX3 U1394 ( .A(n484), .Y(n1233) );
  CLKINVX3 U1395 ( .A(n483), .Y(n1253) );
  CLKINVX3 U1396 ( .A(n482), .Y(n1327) );
  CLKINVX3 U1397 ( .A(n481), .Y(n1245) );
  CLKINVX3 U1398 ( .A(n670), .Y(n1275) );
  CLKINVX3 U1399 ( .A(n672), .Y(n1272) );
  CLKINVX3 U1400 ( .A(n671), .Y(n1269) );
  CLKINVX3 U1401 ( .A(n669), .Y(n1278) );
  AOI211X1 U1402 ( .A0(n150), .A1(n3320), .B0(n5920), .C0(n5913), .Y(n8092) );
  AOI211X1 U1403 ( .A0(n149), .A1(n3142), .B0(n5684), .C0(n5677), .Y(n8968) );
  AOI211X1 U1404 ( .A0(n148), .A1(n2962), .B0(n5456), .C0(n5449), .Y(n9844) );
  AOI211X1 U1405 ( .A0(n147), .A1(n2779), .B0(n5210), .C0(n5203), .Y(n10720)
         );
  AOI211X1 U1406 ( .A0(n146), .A1(n2603), .B0(n4902), .C0(n4895), .Y(n11596)
         );
  AOI211X1 U1407 ( .A0(n145), .A1(n3383), .B0(n5996), .C0(n5989), .Y(n7800) );
  AOI211X1 U1408 ( .A0(n144), .A1(n3200), .B0(n5760), .C0(n5753), .Y(n8676) );
  AOI211X1 U1409 ( .A0(n143), .A1(n3023), .B0(n5532), .C0(n5525), .Y(n9552) );
  AOI211X1 U1410 ( .A0(n142), .A1(n2841), .B0(n5288), .C0(n5281), .Y(n10428)
         );
  AOI211X1 U1411 ( .A0(n141), .A1(n3436), .B0(n6072), .C0(n6065), .Y(n7508) );
  AOI211X1 U1412 ( .A0(n140), .A1(n3086), .B0(n5608), .C0(n5601), .Y(n9260) );
  AOI211X1 U1413 ( .A0(n139), .A1(n2714), .B0(n5102), .C0(n5095), .Y(n11012)
         );
  AOI211X1 U1414 ( .A0(n138), .A1(n3261), .B0(n5844), .C0(n5837), .Y(n8384) );
  AOI211X1 U1415 ( .A0(n137), .A1(n2664), .B0(n5018), .C0(n5011), .Y(n11304)
         );
  AOI211X1 U1416 ( .A0(n136), .A1(n3502), .B0(n6162), .C0(n6155), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n322) );
  AOI211X1 U1417 ( .A0(n135), .A1(n2901), .B0(n5372), .C0(n5365), .Y(n10136)
         );
  OAI221XL U1418 ( .A0(n13355), .A1(n13228), .B0(n1688), .B1(n52), .C0(n13350), 
        .Y(n13518) );
  CLKINVX3 U1419 ( .A(n748), .Y(n13355) );
  CLKINVX3 U1420 ( .A(n752), .Y(n12409) );
  CLKINVX3 U1421 ( .A(n755), .Y(n12094) );
  CLKINVX3 U1422 ( .A(n753), .Y(n11778) );
  CLKINVX3 U1423 ( .A(n754), .Y(top_core_KE_sb1_n206) );
  CLKINVX3 U1424 ( .A(n663), .Y(n15866) );
  CLKINVX3 U1425 ( .A(n661), .Y(n17756) );
  CLKINVX3 U1426 ( .A(n659), .Y(n14606) );
  CLKINVX3 U1427 ( .A(n657), .Y(n16496) );
  CLKINVX3 U1428 ( .A(n655), .Y(n16811) );
  CLKINVX3 U1429 ( .A(n652), .Y(n15236) );
  CLKINVX3 U1430 ( .A(n651), .Y(n18386) );
  CLKINVX3 U1431 ( .A(n650), .Y(n17126) );
  CLKINVX3 U1432 ( .A(n649), .Y(n13976) );
  CLKINVX3 U1433 ( .A(n664), .Y(n17441) );
  CLKINVX3 U1434 ( .A(n660), .Y(n16181) );
  CLKINVX3 U1435 ( .A(n662), .Y(n14291) );
  CLKINVX3 U1436 ( .A(n658), .Y(n18071) );
  CLKINVX3 U1437 ( .A(n656), .Y(n14921) );
  CLKINVX3 U1438 ( .A(n653), .Y(n15551) );
  CLKINVX3 U1439 ( .A(n654), .Y(n18701) );
  OAI221XL U1440 ( .A0(n677), .A1(n52), .B0(n13295), .B1(n1690), .C0(n13475), 
        .Y(n13470) );
  CLKINVX3 U1441 ( .A(n756), .Y(n13295) );
  NAND2X2 U1442 ( .A(n86), .B(top_core_io_n38), .Y(n296) );
  NAND2X2 U1443 ( .A(top_core_io_n211), .B(n302), .Y(n288) );
  NAND2X2 U1444 ( .A(n304), .B(top_core_io_n49), .Y(n291) );
  NAND2X2 U1445 ( .A(top_core_io_n495), .B(n303), .Y(n270) );
  NOR2X1 U1446 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n71), .B(n3500), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n241) );
  NAND2X1 U1447 ( .A(n564), .B(n8139), .Y(n8258) );
  NAND2X1 U1448 ( .A(n561), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n196) );
  NAND2X1 U1449 ( .A(n7844), .B(n7843), .Y(n7944) );
  NAND2X1 U1450 ( .A(n8720), .B(n8719), .Y(n8820) );
  NAND2X1 U1451 ( .A(n9596), .B(n9595), .Y(n9696) );
  NAND2X1 U1452 ( .A(n10472), .B(n10471), .Y(n10572) );
  NAND2X1 U1453 ( .A(n11348), .B(n11347), .Y(n11448) );
  NAND2X1 U1454 ( .A(n7552), .B(n7551), .Y(n7652) );
  NAND2X1 U1455 ( .A(n8428), .B(n8427), .Y(n8528) );
  NAND2X1 U1456 ( .A(n9304), .B(n9303), .Y(n9404) );
  NAND2X1 U1457 ( .A(n10180), .B(n10179), .Y(n10280) );
  NAND2X1 U1458 ( .A(n7260), .B(n7259), .Y(n7360) );
  NAND2X1 U1459 ( .A(n9012), .B(n9011), .Y(n9112) );
  NAND2X1 U1460 ( .A(n10764), .B(n10763), .Y(n10864) );
  NAND2X1 U1461 ( .A(n8136), .B(n8135), .Y(n8236) );
  NAND2X1 U1462 ( .A(n11056), .B(n11055), .Y(n11156) );
  NAND2X1 U1463 ( .A(n9888), .B(n9887), .Y(n9988) );
  NAND2X1 U1464 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n70), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n69), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n174) );
  NOR2XL U1465 ( .A(n5), .B(n582), .Y(n260) );
  NOR2XL U1466 ( .A(n6), .B(n583), .Y(n261) );
  NOR2XL U1467 ( .A(n4), .B(n584), .Y(n262) );
  NOR2XL U1468 ( .A(n3), .B(n580), .Y(n263) );
  NOR2X1 U1469 ( .A(n29), .B(n368), .Y(n7942) );
  NOR2X1 U1470 ( .A(n28), .B(n367), .Y(n8818) );
  NOR2X1 U1471 ( .A(n27), .B(n366), .Y(n9694) );
  NOR2X1 U1472 ( .A(n26), .B(n365), .Y(n10570) );
  NOR2X1 U1473 ( .A(n25), .B(n364), .Y(n11446) );
  NOR2X1 U1474 ( .A(n24), .B(n363), .Y(n7650) );
  NOR2X1 U1475 ( .A(n23), .B(n362), .Y(n8526) );
  NOR2X1 U1476 ( .A(n22), .B(n361), .Y(n9402) );
  NOR2X1 U1477 ( .A(n21), .B(n360), .Y(n10278) );
  NOR2X1 U1478 ( .A(n20), .B(n358), .Y(n7358) );
  NOR2X1 U1479 ( .A(n19), .B(n359), .Y(n9110) );
  NOR2X1 U1480 ( .A(n18), .B(n357), .Y(n10862) );
  NOR2X1 U1481 ( .A(n17), .B(n355), .Y(n8234) );
  NOR2X1 U1482 ( .A(n16), .B(n356), .Y(n11154) );
  NOR2X1 U1483 ( .A(n14), .B(n354), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n172) );
  NOR2X1 U1484 ( .A(n15), .B(n353), .Y(n9986) );
  AOI221X1 U1485 ( .A0(n6151), .A1(n3483), .B0(n6117), .B1(n1280), .C0(n13853), 
        .Y(n13852) );
  AOI221X1 U1486 ( .A0(n5464), .A1(n2943), .B0(n5418), .B1(n1307), .C0(n16688), 
        .Y(n16687) );
  AOI221X1 U1487 ( .A0(n5296), .A1(n2822), .B0(n5250), .B1(n1313), .C0(n17318), 
        .Y(n17317) );
  AOI221X1 U1488 ( .A0(n5616), .A1(n3062), .B0(n5570), .B1(n1301), .C0(n16058), 
        .Y(n16057) );
  AOI221X1 U1489 ( .A0(n5928), .A1(n3303), .B0(n5882), .B1(n1289), .C0(n14798), 
        .Y(n14797) );
  AOI221X1 U1490 ( .A0(n6080), .A1(n3422), .B0(n6034), .B1(n1283), .C0(n14168), 
        .Y(n14167) );
  AOI221X1 U1491 ( .A0(n5110), .A1(n2701), .B0(n5064), .B1(n1319), .C0(n17948), 
        .Y(n17947) );
  AOI221X1 U1492 ( .A0(n5026), .A1(n2640), .B0(n4980), .B1(n1322), .C0(n18263), 
        .Y(n18262) );
  AOI221X1 U1493 ( .A0(n5852), .A1(n3242), .B0(n5806), .B1(n1292), .C0(n15113), 
        .Y(n15112) );
  AOI221X1 U1494 ( .A0(n5380), .A1(n2882), .B0(n5334), .B1(n1310), .C0(n17003), 
        .Y(n17002) );
  AOI221X1 U1495 ( .A0(n5768), .A1(n3181), .B0(n5722), .B1(n1295), .C0(n15428), 
        .Y(n15427) );
  AOI221X1 U1496 ( .A0(n5692), .A1(n3123), .B0(n5646), .B1(n1298), .C0(n15743), 
        .Y(n15742) );
  AOI221X1 U1497 ( .A0(n6004), .A1(n3364), .B0(n5958), .B1(n1286), .C0(n14483), 
        .Y(n14482) );
  AOI221X1 U1498 ( .A0(n5540), .A1(n3004), .B0(n5494), .B1(n1304), .C0(n16373), 
        .Y(n16372) );
  AOI221X1 U1499 ( .A0(n4910), .A1(n2579), .B0(n4864), .B1(n1325), .C0(n18578), 
        .Y(n18577) );
  AOI221X1 U1500 ( .A0(n5218), .A1(n2761), .B0(n5172), .B1(n1316), .C0(n17633), 
        .Y(n17632) );
  AOI211X1 U1501 ( .A0(n1151), .A1(n13223), .B0(n13258), .C0(n6547), .Y(n13368) );
  CLKINVX3 U1502 ( .A(n692), .Y(n13223) );
  OAI211X1 U1503 ( .A0(n13228), .A1(n73), .B0(n13266), .C0(n13453), .Y(n13448)
         );
  OAI211X1 U1504 ( .A0(n12913), .A1(n75), .B0(n12951), .C0(n13138), .Y(n13133)
         );
  OAI211X1 U1505 ( .A0(n12598), .A1(n74), .B0(n12636), .C0(n12823), .Y(n12818)
         );
  OAI211X1 U1506 ( .A0(n13543), .A1(n76), .B0(n13581), .C0(n13768), .Y(n13763)
         );
  CLKINVX3 U1507 ( .A(n721), .Y(n13031) );
  CLKINVX3 U1508 ( .A(n719), .Y(n12716) );
  CLKINVX3 U1509 ( .A(n717), .Y(n13346) );
  CLKINVX3 U1510 ( .A(n720), .Y(n13661) );
  NAND2X2 U1511 ( .A(n86), .B(top_core_io_n49), .Y(n295) );
  NAND2X2 U1512 ( .A(top_core_io_n222), .B(n302), .Y(n287) );
  NAND2X2 U1513 ( .A(top_core_io_n200), .B(n304), .Y(n273) );
  NAND2X2 U1514 ( .A(top_core_io_n506), .B(n303), .Y(n269) );
  AOI222X1 U1515 ( .A0(n760), .A1(n12322), .B0(n1182), .B1(n752), .C0(n683), 
        .C1(n6622), .Y(n12397) );
  CLKINVX3 U1516 ( .A(n627), .Y(n12322) );
  AOI222X1 U1517 ( .A0(n763), .A1(n12007), .B0(n1177), .B1(n755), .C0(n684), 
        .C1(n6575), .Y(n12082) );
  CLKINVX3 U1518 ( .A(n628), .Y(n12007) );
  AOI222X1 U1519 ( .A0(n762), .A1(top_core_KE_sb1_n116), .B0(n1217), .B1(n754), 
        .C0(n682), .C1(n6869), .Y(top_core_KE_sb1_n194) );
  CLKINVX3 U1520 ( .A(n626), .Y(top_core_KE_sb1_n116) );
  AOI222X1 U1521 ( .A0(n761), .A1(n11691), .B0(n1223), .B1(n753), .C0(n681), 
        .C1(n6915), .Y(n11766) );
  CLKINVX3 U1522 ( .A(n625), .Y(n11691) );
  CLKINVX3 U1523 ( .A(n434), .Y(n13897) );
  CLKINVX3 U1524 ( .A(n447), .Y(n15787) );
  CLKINVX3 U1525 ( .A(n445), .Y(n17677) );
  CLKINVX3 U1526 ( .A(n443), .Y(n14527) );
  CLKINVX3 U1527 ( .A(n441), .Y(n16417) );
  CLKINVX3 U1528 ( .A(n438), .Y(n16732) );
  CLKINVX3 U1529 ( .A(n436), .Y(n15157) );
  CLKINVX3 U1530 ( .A(n435), .Y(n18307) );
  CLKINVX3 U1531 ( .A(n433), .Y(n17047) );
  CLKINVX3 U1532 ( .A(n437), .Y(n15472) );
  CLKINVX3 U1533 ( .A(n446), .Y(n14212) );
  CLKINVX3 U1534 ( .A(n442), .Y(n17992) );
  CLKINVX3 U1535 ( .A(n440), .Y(n14842) );
  CLKINVX3 U1536 ( .A(n448), .Y(n17362) );
  CLKINVX3 U1537 ( .A(n444), .Y(n16102) );
  CLKINVX3 U1538 ( .A(n439), .Y(n18622) );
  CLKINVX3 U1539 ( .A(n423), .Y(n7285) );
  CLKINVX3 U1540 ( .A(n420), .Y(n8161) );
  CLKINVX3 U1541 ( .A(n419), .Y(n11081) );
  CLKINVX3 U1542 ( .A(n418), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n97) );
  CLKINVX3 U1543 ( .A(n417), .Y(n9913) );
  CLKINVX3 U1544 ( .A(n431), .Y(n8745) );
  CLKINVX3 U1545 ( .A(n427), .Y(n7577) );
  CLKINVX3 U1546 ( .A(n425), .Y(n9329) );
  CLKINVX3 U1547 ( .A(n429), .Y(n10497) );
  CLKINVX3 U1548 ( .A(n424), .Y(n10205) );
  CLKINVX3 U1549 ( .A(n432), .Y(n7869) );
  CLKINVX3 U1550 ( .A(n428), .Y(n11373) );
  CLKINVX3 U1551 ( .A(n421), .Y(n10789) );
  CLKINVX3 U1552 ( .A(n430), .Y(n9621) );
  CLKINVX3 U1553 ( .A(n426), .Y(n8453) );
  CLKINVX3 U1554 ( .A(n422), .Y(n9037) );
  NAND2X1 U1555 ( .A(n5678), .B(n8802), .Y(n8793) );
  INVX4 U1556 ( .A(n415), .Y(n8802) );
  NAND2X1 U1557 ( .A(n5204), .B(n10554), .Y(n10545) );
  INVX4 U1558 ( .A(n413), .Y(n10554) );
  NAND2X1 U1559 ( .A(n5990), .B(n7634), .Y(n7625) );
  INVX4 U1560 ( .A(n411), .Y(n7634) );
  NAND2X1 U1561 ( .A(n5526), .B(n9386), .Y(n9377) );
  INVX4 U1562 ( .A(n409), .Y(n9386) );
  NAND2X1 U1563 ( .A(n6066), .B(n7342), .Y(n7333) );
  INVX4 U1564 ( .A(n407), .Y(n7342) );
  NAND2X1 U1565 ( .A(n5838), .B(n8218), .Y(n8209) );
  INVX4 U1566 ( .A(n404), .Y(n8218) );
  NAND2X1 U1567 ( .A(n5012), .B(n11138), .Y(n11129) );
  INVX4 U1568 ( .A(n403), .Y(n11138) );
  NAND2X1 U1569 ( .A(n6156), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n146) );
  INVX4 U1570 ( .A(n402), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n156) );
  NAND2X1 U1571 ( .A(n5366), .B(n9970), .Y(n9961) );
  INVX4 U1572 ( .A(n401), .Y(n9970) );
  NAND2X1 U1573 ( .A(n5096), .B(n10846), .Y(n10837) );
  INVX4 U1574 ( .A(n405), .Y(n10846) );
  NAND2X1 U1575 ( .A(n5282), .B(n10262), .Y(n10253) );
  INVX4 U1576 ( .A(n408), .Y(n10262) );
  NAND2X1 U1577 ( .A(n5450), .B(n9678), .Y(n9669) );
  INVX4 U1578 ( .A(n414), .Y(n9678) );
  NAND2X1 U1579 ( .A(n5754), .B(n8510), .Y(n8501) );
  INVX4 U1580 ( .A(n410), .Y(n8510) );
  NAND2X1 U1581 ( .A(n5914), .B(n7926), .Y(n7917) );
  INVX4 U1582 ( .A(n416), .Y(n7926) );
  NAND2X1 U1583 ( .A(n4896), .B(n11430), .Y(n11421) );
  INVX4 U1584 ( .A(n412), .Y(n11430) );
  NAND2X1 U1585 ( .A(n5602), .B(n9094), .Y(n9085) );
  INVX4 U1586 ( .A(n406), .Y(n9094) );
  NOR2X1 U1587 ( .A(n29), .B(n3320), .Y(n7877) );
  NOR2X1 U1588 ( .A(n28), .B(n3140), .Y(n8753) );
  NOR2X1 U1589 ( .A(n27), .B(n2958), .Y(n9629) );
  NOR2X1 U1590 ( .A(n26), .B(n2780), .Y(n10505) );
  NOR2X1 U1591 ( .A(n25), .B(n2593), .Y(n11381) );
  NOR2X1 U1592 ( .A(n24), .B(n3381), .Y(n7585) );
  NOR2X1 U1593 ( .A(n23), .B(n3196), .Y(n8461) );
  NOR2X1 U1594 ( .A(n22), .B(n3021), .Y(n9337) );
  NOR2X1 U1595 ( .A(n21), .B(n2840), .Y(n10213) );
  NOR2X1 U1596 ( .A(n20), .B(n3437), .Y(n7293) );
  NOR2X1 U1597 ( .A(n19), .B(n3076), .Y(n9045) );
  NOR2X1 U1598 ( .A(n18), .B(n2715), .Y(n10797) );
  NOR2X1 U1599 ( .A(n17), .B(n3257), .Y(n8169) );
  NOR2X1 U1600 ( .A(n16), .B(n2654), .Y(n11089) );
  NOR2X1 U1601 ( .A(n14), .B(n3502), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n106) );
  NOR2X1 U1602 ( .A(n15), .B(n2897), .Y(n9921) );
  NOR2X1 U1603 ( .A(n7847), .B(n7844), .Y(n7956) );
  CLKINVX3 U1604 ( .A(n600), .Y(n7844) );
  NOR2X1 U1605 ( .A(n9599), .B(n9596), .Y(n9708) );
  CLKINVX3 U1606 ( .A(n598), .Y(n9596) );
  NOR2X1 U1607 ( .A(n11351), .B(n11348), .Y(n11460) );
  CLKINVX3 U1608 ( .A(n596), .Y(n11348) );
  NOR2X1 U1609 ( .A(n8431), .B(n8428), .Y(n8540) );
  CLKINVX3 U1610 ( .A(n594), .Y(n8428) );
  NOR2X1 U1611 ( .A(n10183), .B(n10180), .Y(n10292) );
  CLKINVX3 U1612 ( .A(n592), .Y(n10180) );
  NOR2X1 U1613 ( .A(n7263), .B(n7260), .Y(n7372) );
  CLKINVX3 U1614 ( .A(n591), .Y(n7260) );
  NOR2X1 U1615 ( .A(n9015), .B(n9012), .Y(n9124) );
  CLKINVX3 U1616 ( .A(n590), .Y(n9012) );
  NOR2X1 U1617 ( .A(n10767), .B(n10764), .Y(n10876) );
  CLKINVX3 U1618 ( .A(n589), .Y(n10764) );
  NOR2XL U1619 ( .A(n8139), .B(n8136), .Y(n264) );
  CLKINVX3 U1620 ( .A(n588), .Y(n8136) );
  CLKINVX3 U1621 ( .A(n355), .Y(n8139) );
  NOR2X1 U1622 ( .A(n11059), .B(n11056), .Y(n11168) );
  CLKINVX3 U1623 ( .A(n587), .Y(n11056) );
  NOR2XL U1624 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n70), .Y(n265) );
  CLKINVX3 U1625 ( .A(n585), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n70) );
  CLKINVX3 U1626 ( .A(n354), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n74) );
  NOR2X1 U1627 ( .A(n9891), .B(n9888), .Y(n10000) );
  CLKINVX3 U1628 ( .A(n586), .Y(n9888) );
  NOR2X1 U1629 ( .A(n8723), .B(n8720), .Y(n8832) );
  CLKINVX3 U1630 ( .A(n599), .Y(n8720) );
  NOR2X1 U1631 ( .A(n7555), .B(n7552), .Y(n7664) );
  CLKINVX3 U1632 ( .A(n595), .Y(n7552) );
  NOR2X1 U1633 ( .A(n9307), .B(n9304), .Y(n9416) );
  CLKINVX3 U1634 ( .A(n593), .Y(n9304) );
  NOR2X1 U1635 ( .A(n10475), .B(n10472), .Y(n10584) );
  CLKINVX3 U1636 ( .A(n597), .Y(n10472) );
  NOR2X1 U1637 ( .A(n7845), .B(n3313), .Y(n7994) );
  CLKINVX3 U1638 ( .A(n576), .Y(n7845) );
  NOR2X1 U1639 ( .A(n8721), .B(n3133), .Y(n8870) );
  CLKINVX3 U1640 ( .A(n575), .Y(n8721) );
  NOR2X1 U1641 ( .A(n9597), .B(n2953), .Y(n9746) );
  CLKINVX3 U1642 ( .A(n574), .Y(n9597) );
  NOR2X1 U1643 ( .A(n10473), .B(n2771), .Y(n10622) );
  CLKINVX3 U1644 ( .A(n573), .Y(n10473) );
  NOR2X1 U1645 ( .A(n11349), .B(n2589), .Y(n11498) );
  CLKINVX3 U1646 ( .A(n572), .Y(n11349) );
  NOR2X1 U1647 ( .A(n7553), .B(n3374), .Y(n7702) );
  CLKINVX3 U1648 ( .A(n571), .Y(n7553) );
  NOR2X1 U1649 ( .A(n8429), .B(n3191), .Y(n8578) );
  CLKINVX3 U1650 ( .A(n570), .Y(n8429) );
  NOR2X1 U1651 ( .A(n9305), .B(n3014), .Y(n9454) );
  CLKINVX3 U1652 ( .A(n569), .Y(n9305) );
  NOR2X1 U1653 ( .A(n10181), .B(n2832), .Y(n10330) );
  CLKINVX3 U1654 ( .A(n568), .Y(n10181) );
  NOR2X1 U1655 ( .A(n7261), .B(n3432), .Y(n7410) );
  CLKINVX3 U1656 ( .A(n567), .Y(n7261) );
  NOR2X1 U1657 ( .A(n9013), .B(n3081), .Y(n9162) );
  CLKINVX3 U1658 ( .A(n566), .Y(n9013) );
  NOR2X1 U1659 ( .A(n10765), .B(n2710), .Y(n10914) );
  CLKINVX3 U1660 ( .A(n565), .Y(n10765) );
  NOR2X1 U1661 ( .A(n8137), .B(n3252), .Y(n8286) );
  CLKINVX3 U1662 ( .A(n564), .Y(n8137) );
  NOR2X1 U1663 ( .A(n11057), .B(n2659), .Y(n11206) );
  CLKINVX3 U1664 ( .A(n563), .Y(n11057) );
  NOR2X1 U1665 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n71), .B(n3493), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n224) );
  CLKINVX3 U1666 ( .A(n561), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n71) );
  NOR2X1 U1667 ( .A(n9889), .B(n2892), .Y(n10038) );
  CLKINVX3 U1668 ( .A(n562), .Y(n9889) );
  NAND2X1 U1669 ( .A(n576), .B(n7847), .Y(n7966) );
  CLKINVX3 U1670 ( .A(n368), .Y(n7847) );
  NAND2X1 U1671 ( .A(n575), .B(n8723), .Y(n8842) );
  CLKINVX3 U1672 ( .A(n367), .Y(n8723) );
  NAND2X1 U1673 ( .A(n574), .B(n9599), .Y(n9718) );
  CLKINVX3 U1674 ( .A(n366), .Y(n9599) );
  NAND2X1 U1675 ( .A(n573), .B(n10475), .Y(n10594) );
  CLKINVX3 U1676 ( .A(n365), .Y(n10475) );
  NAND2X1 U1677 ( .A(n572), .B(n11351), .Y(n11470) );
  CLKINVX3 U1678 ( .A(n364), .Y(n11351) );
  NAND2X1 U1679 ( .A(n571), .B(n7555), .Y(n7674) );
  CLKINVX3 U1680 ( .A(n363), .Y(n7555) );
  NAND2X1 U1681 ( .A(n570), .B(n8431), .Y(n8550) );
  CLKINVX3 U1682 ( .A(n362), .Y(n8431) );
  NAND2X1 U1683 ( .A(n569), .B(n9307), .Y(n9426) );
  CLKINVX3 U1684 ( .A(n361), .Y(n9307) );
  NAND2X1 U1685 ( .A(n568), .B(n10183), .Y(n10302) );
  CLKINVX3 U1686 ( .A(n360), .Y(n10183) );
  NAND2X1 U1687 ( .A(n567), .B(n7263), .Y(n7382) );
  CLKINVX3 U1688 ( .A(n358), .Y(n7263) );
  NAND2X1 U1689 ( .A(n566), .B(n9015), .Y(n9134) );
  CLKINVX3 U1690 ( .A(n359), .Y(n9015) );
  NAND2X1 U1691 ( .A(n565), .B(n10767), .Y(n10886) );
  CLKINVX3 U1692 ( .A(n357), .Y(n10767) );
  NAND2X1 U1693 ( .A(n563), .B(n11059), .Y(n11178) );
  CLKINVX3 U1694 ( .A(n356), .Y(n11059) );
  NAND2X1 U1695 ( .A(n562), .B(n9891), .Y(n10010) );
  CLKINVX3 U1696 ( .A(n353), .Y(n9891) );
  NAND2X1 U1697 ( .A(n105), .B(n7900), .Y(n7952) );
  NAND2X1 U1698 ( .A(n104), .B(n8776), .Y(n8828) );
  NAND2X1 U1699 ( .A(n103), .B(n9652), .Y(n9704) );
  NAND2X1 U1700 ( .A(n102), .B(n10528), .Y(n10580) );
  NAND2X1 U1701 ( .A(n101), .B(n11404), .Y(n11456) );
  NAND2X1 U1702 ( .A(n100), .B(n7608), .Y(n7660) );
  NAND2X1 U1703 ( .A(n99), .B(n8484), .Y(n8536) );
  NAND2X1 U1704 ( .A(n98), .B(n9360), .Y(n9412) );
  NAND2X1 U1705 ( .A(n97), .B(n10236), .Y(n10288) );
  NAND2X1 U1706 ( .A(n96), .B(n9068), .Y(n9120) );
  NAND2X1 U1707 ( .A(n95), .B(n7316), .Y(n7368) );
  NAND2X1 U1708 ( .A(n94), .B(n10820), .Y(n10872) );
  NAND2X1 U1709 ( .A(n92), .B(n11112), .Y(n11164) );
  NAND2X1 U1710 ( .A(n93), .B(n8192), .Y(n8244) );
  NAND2X1 U1711 ( .A(n91), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n129), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n182) );
  NAND2X1 U1712 ( .A(n90), .B(n9944), .Y(n9996) );
  CLKINVX3 U1713 ( .A(n667), .Y(n1266) );
  CLKINVX3 U1714 ( .A(n668), .Y(n1262) );
  CLKINVX3 U1715 ( .A(n666), .Y(n1331) );
  CLKINVX3 U1716 ( .A(n665), .Y(n1259) );
  NOR2BX2 U1717 ( .AN(top_core_KE_n2700), .B(top_core_KE_n918), .Y(
        top_core_KE_n1873) );
  NOR2X1 U1718 ( .A(n180), .B(n1683), .Y(n13393) );
  NOR2X1 U1719 ( .A(n183), .B(n1654), .Y(n13708) );
  NOR2X1 U1720 ( .A(n182), .B(n1712), .Y(n13078) );
  NOR2X1 U1721 ( .A(n181), .B(n1741), .Y(n12763) );
  NOR2X1 U1722 ( .A(n170), .B(n2945), .Y(n16858) );
  NOR2X1 U1723 ( .A(n79), .B(n1784), .Y(n12133) );
  NOR2X1 U1724 ( .A(n77), .B(n1805), .Y(n11817) );
  NOR2X1 U1725 ( .A(n184), .B(n1763), .Y(n12448) );
  NOR2X1 U1726 ( .A(n78), .B(n1826), .Y(top_core_KE_sb1_n245) );
  NOR2X1 U1727 ( .A(n165), .B(n3485), .Y(n14023) );
  NOR2X1 U1728 ( .A(n167), .B(n3244), .Y(n15283) );
  NOR2X1 U1729 ( .A(n166), .B(n2644), .Y(n18433) );
  NOR2X1 U1730 ( .A(n164), .B(n2886), .Y(n17173) );
  NOR2X1 U1731 ( .A(n178), .B(n3124), .Y(n15913) );
  NOR2X1 U1732 ( .A(n174), .B(n3365), .Y(n14653) );
  NOR2X1 U1733 ( .A(n172), .B(n3006), .Y(n16543) );
  NOR2X1 U1734 ( .A(n176), .B(n2762), .Y(n17803) );
  NOR2X1 U1735 ( .A(n168), .B(n3182), .Y(n15598) );
  NOR2X1 U1736 ( .A(n171), .B(n3305), .Y(n14968) );
  NOR2X1 U1737 ( .A(n177), .B(n3426), .Y(n14338) );
  NOR2X1 U1738 ( .A(n173), .B(n2702), .Y(n18118) );
  NOR2X1 U1739 ( .A(n179), .B(n2824), .Y(n17488) );
  NOR2X1 U1740 ( .A(n175), .B(n3064), .Y(n16228) );
  NOR2X1 U1741 ( .A(n169), .B(n2580), .Y(n18748) );
  CLKINVX3 U1742 ( .A(n750), .Y(n13040) );
  CLKINVX3 U1743 ( .A(n749), .Y(n12725) );
  CLKINVX3 U1744 ( .A(n639), .Y(n16820) );
  CLKINVX3 U1745 ( .A(n751), .Y(n13670) );
  CLKINVX3 U1746 ( .A(n636), .Y(n15245) );
  CLKINVX3 U1747 ( .A(n635), .Y(n18395) );
  CLKINVX3 U1748 ( .A(n634), .Y(n13985) );
  CLKINVX3 U1749 ( .A(n633), .Y(n17135) );
  CLKINVX3 U1750 ( .A(n647), .Y(n15875) );
  CLKINVX3 U1751 ( .A(n643), .Y(n14615) );
  CLKINVX3 U1752 ( .A(n641), .Y(n16505) );
  CLKINVX3 U1753 ( .A(n645), .Y(n17765) );
  CLKINVX3 U1754 ( .A(n646), .Y(n14300) );
  CLKINVX3 U1755 ( .A(n642), .Y(n18080) );
  CLKINVX3 U1756 ( .A(n637), .Y(n15560) );
  CLKINVX3 U1757 ( .A(n648), .Y(n17450) );
  CLKINVX3 U1758 ( .A(n644), .Y(n16190) );
  CLKINVX3 U1759 ( .A(n640), .Y(n14930) );
  CLKINVX3 U1760 ( .A(n638), .Y(n18710) );
  CLKINVX3 U1761 ( .A(n716), .Y(n12400) );
  CLKINVX3 U1762 ( .A(n714), .Y(n11769) );
  CLKINVX3 U1763 ( .A(n715), .Y(top_core_KE_sb1_n197) );
  CLKINVX3 U1764 ( .A(n718), .Y(n12085) );
  NAND2X2 U1765 ( .A(n86), .B(top_core_io_n60), .Y(n294) );
  NAND2X2 U1766 ( .A(top_core_io_n233), .B(n302), .Y(n286) );
  NAND2X2 U1767 ( .A(top_core_io_n211), .B(n304), .Y(n272) );
  NAND2X2 U1768 ( .A(top_core_io_n517), .B(n303), .Y(n268) );
  CLKINVX3 U1769 ( .A(n743), .Y(top_core_KE_n1865) );
  NAND3X1 U1770 ( .A(n6308), .B(n4256), .C(n1), .Y(top_core_EC_n1011) );
  CLKINVX3 U1771 ( .A(n551), .Y(n7268) );
  CLKINVX3 U1772 ( .A(n552), .Y(n10188) );
  CLKINVX3 U1773 ( .A(n560), .Y(n7852) );
  CLKINVX3 U1774 ( .A(n556), .Y(n11356) );
  CLKINVX3 U1775 ( .A(n548), .Y(n8144) );
  CLKINVX3 U1776 ( .A(n547), .Y(n11064) );
  CLKINVX3 U1777 ( .A(n546), .Y(n9896) );
  CLKINVX3 U1778 ( .A(n545), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n79) );
  CLKINVX3 U1779 ( .A(n559), .Y(n8728) );
  CLKINVX3 U1780 ( .A(n555), .Y(n7560) );
  CLKINVX3 U1781 ( .A(n553), .Y(n9312) );
  CLKINVX3 U1782 ( .A(n550), .Y(n9020) );
  CLKINVX3 U1783 ( .A(n557), .Y(n10480) );
  CLKINVX3 U1784 ( .A(n558), .Y(n9604) );
  CLKINVX3 U1785 ( .A(n554), .Y(n8436) );
  CLKINVX3 U1786 ( .A(n549), .Y(n10772) );
  AOI222X1 U1787 ( .A0(n756), .A1(n13268), .B0(n610), .B1(n748), .C0(n686), 
        .C1(n6550), .Y(n13343) );
  CLKINVX3 U1788 ( .A(n629), .Y(n13268) );
  AOI222X1 U1789 ( .A0(n758), .A1(n12953), .B0(n612), .B1(n750), .C0(n687), 
        .C1(n6891), .Y(n13028) );
  CLKINVX3 U1790 ( .A(n632), .Y(n12953) );
  AOI222X1 U1791 ( .A0(n757), .A1(n12638), .B0(n611), .B1(n749), .C0(n688), 
        .C1(n6845), .Y(n12713) );
  CLKINVX3 U1792 ( .A(n630), .Y(n12638) );
  AOI222X1 U1793 ( .A0(n759), .A1(n13583), .B0(n616), .B1(n751), .C0(n685), 
        .C1(n6598), .Y(n13658) );
  CLKINVX3 U1794 ( .A(n631), .Y(n13583) );
  CLKINVX3 U1795 ( .A(n580), .Y(n13228) );
  CLKINVX3 U1796 ( .A(n582), .Y(n12913) );
  CLKINVX3 U1797 ( .A(n584), .Y(n12598) );
  CLKINVX3 U1798 ( .A(n583), .Y(n13543) );
  CLKINVX3 U1799 ( .A(n342), .Y(n16692) );
  CLKINVX3 U1800 ( .A(n352), .Y(n17322) );
  CLKINVX3 U1801 ( .A(n348), .Y(n16062) );
  CLKINVX3 U1802 ( .A(n344), .Y(n14802) );
  CLKINVX3 U1803 ( .A(n350), .Y(n14172) );
  CLKINVX3 U1804 ( .A(n346), .Y(n17952) );
  CLKINVX3 U1805 ( .A(n341), .Y(n15432) );
  CLKINVX3 U1806 ( .A(n340), .Y(n15117) );
  CLKINVX3 U1807 ( .A(n339), .Y(n18267) );
  CLKINVX3 U1808 ( .A(n338), .Y(n13857) );
  CLKINVX3 U1809 ( .A(n337), .Y(n17007) );
  CLKINVX3 U1810 ( .A(n351), .Y(n15747) );
  CLKINVX3 U1811 ( .A(n347), .Y(n14487) );
  CLKINVX3 U1812 ( .A(n345), .Y(n16377) );
  CLKINVX3 U1813 ( .A(n349), .Y(n17637) );
  CLKINVX3 U1814 ( .A(n343), .Y(n18582) );
  CLKINVX3 U1815 ( .A(n581), .Y(n11967) );
  CLKINVX3 U1816 ( .A(n578), .Y(top_core_KE_sb1_n76) );
  CLKINVX3 U1817 ( .A(n577), .Y(n11651) );
  CLKINVX3 U1818 ( .A(n579), .Y(n12283) );
  INVX4 U1819 ( .A(n326), .Y(n7272) );
  INVX4 U1820 ( .A(n328), .Y(n10192) );
  INVX4 U1821 ( .A(n327), .Y(n9024) );
  INVX4 U1822 ( .A(n336), .Y(n7856) );
  INVX4 U1823 ( .A(n332), .Y(n11360) );
  INVX4 U1824 ( .A(n325), .Y(n10776) );
  INVX4 U1825 ( .A(n334), .Y(n9608) );
  INVX4 U1826 ( .A(n330), .Y(n8440) );
  INVX4 U1827 ( .A(n323), .Y(n11068) );
  INVX4 U1828 ( .A(n322), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n83) );
  INVX4 U1829 ( .A(n324), .Y(n8148) );
  INVX4 U1830 ( .A(n321), .Y(n9900) );
  INVX4 U1831 ( .A(n335), .Y(n8732) );
  INVX4 U1832 ( .A(n331), .Y(n7564) );
  INVX4 U1833 ( .A(n329), .Y(n9316) );
  INVX4 U1834 ( .A(n333), .Y(n10484) );
  AOI222XL U1835 ( .A0(n5341), .A1(n2884), .B0(n5350), .B1(n9913), .C0(n5366), 
        .C1(n9891), .Y(n10037) );
  AOI222XL U1836 ( .A0(n6137), .A1(n3487), .B0(n6146), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .C0(n6156), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n74), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n223) );
  AOI222XL U1837 ( .A0(n4987), .A1(n2643), .B0(n4996), .B1(n11081), .C0(n5012), 
        .C1(n11059), .Y(n11205) );
  AOI222XL U1838 ( .A0(n5813), .A1(n3245), .B0(n5822), .B1(n8161), .C0(n5838), 
        .C1(n8139), .Y(n8285) );
  AOI222XL U1839 ( .A0(n5071), .A1(n2705), .B0(n5080), .B1(n10789), .C0(n5096), 
        .C1(n10767), .Y(n10913) );
  AOI222XL U1840 ( .A0(n5577), .A1(n3063), .B0(n5586), .B1(n9037), .C0(n5602), 
        .C1(n9015), .Y(n9161) );
  AOI222XL U1841 ( .A0(n6041), .A1(n3425), .B0(n6050), .B1(n7285), .C0(n6066), 
        .C1(n7263), .Y(n7409) );
  AOI222XL U1842 ( .A0(n5257), .A1(n2823), .B0(n5266), .B1(n10205), .C0(n5282), 
        .C1(n10183), .Y(n10329) );
  AOI222XL U1843 ( .A0(n5501), .A1(n3007), .B0(n5510), .B1(n9329), .C0(n5526), 
        .C1(n9307), .Y(n9453) );
  AOI222XL U1844 ( .A0(n5729), .A1(n3185), .B0(n5738), .B1(n8453), .C0(n5754), 
        .C1(n8431), .Y(n8577) );
  AOI222XL U1845 ( .A0(n5965), .A1(n3368), .B0(n5974), .B1(n7577), .C0(n5990), 
        .C1(n7555), .Y(n7701) );
  AOI222XL U1846 ( .A0(n4871), .A1(n2583), .B0(n4880), .B1(n11373), .C0(n4896), 
        .C1(n11351), .Y(n11497) );
  AOI222XL U1847 ( .A0(n5179), .A1(n2765), .B0(n5188), .B1(n10497), .C0(n5204), 
        .C1(n10475), .Y(n10621) );
  AOI222XL U1848 ( .A0(n5425), .A1(n2947), .B0(n5434), .B1(n9621), .C0(n5450), 
        .C1(n9599), .Y(n9745) );
  AOI222XL U1849 ( .A0(n5653), .A1(n3127), .B0(n5662), .B1(n8745), .C0(n5678), 
        .C1(n8723), .Y(n8869) );
  AOI222XL U1850 ( .A0(n5889), .A1(n3306), .B0(n5898), .B1(n7869), .C0(n5914), 
        .C1(n7847), .Y(n7993) );
  AOI22XL U1851 ( .A0(n6169), .A1(n3495), .B0(n545), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n113) );
  AOI22XL U1852 ( .A0(n5384), .A1(n2901), .B0(n546), .B1(n9900), .Y(n9928) );
  AOI22XL U1853 ( .A0(n5030), .A1(n2663), .B0(n547), .B1(n11068), .Y(n11096)
         );
  AOI22XL U1854 ( .A0(n5856), .A1(n3261), .B0(n548), .B1(n8148), .Y(n8176) );
  AOI22XL U1855 ( .A0(n5114), .A1(n2713), .B0(n549), .B1(n10776), .Y(n10804)
         );
  AOI22XL U1856 ( .A0(n5620), .A1(n3085), .B0(n550), .B1(n9024), .Y(n9052) );
  AOI22XL U1857 ( .A0(n6084), .A1(n3435), .B0(n551), .B1(n7272), .Y(n7300) );
  AOI22XL U1858 ( .A0(n5300), .A1(n2835), .B0(n552), .B1(n10192), .Y(n10220)
         );
  AOI22XL U1859 ( .A0(n5544), .A1(n3025), .B0(n553), .B1(n9316), .Y(n9344) );
  AOI22XL U1860 ( .A0(n5772), .A1(n3200), .B0(n554), .B1(n8440), .Y(n8468) );
  AOI22XL U1861 ( .A0(n6008), .A1(n3385), .B0(n555), .B1(n7564), .Y(n7592) );
  AOI22XL U1862 ( .A0(n4914), .A1(n2602), .B0(n556), .B1(n11360), .Y(n11388)
         );
  AOI22XL U1863 ( .A0(n5222), .A1(n2774), .B0(n557), .B1(n10484), .Y(n10512)
         );
  AOI22XL U1864 ( .A0(n5468), .A1(n2962), .B0(n558), .B1(n9608), .Y(n9636) );
  AOI22XL U1865 ( .A0(n5696), .A1(n3144), .B0(n559), .B1(n8732), .Y(n8760) );
  AOI22XL U1866 ( .A0(n5932), .A1(n3315), .B0(n560), .B1(n7856), .Y(n7884) );
  AOI211XL U1867 ( .A0(n1615), .A1(n2872), .B0(n5339), .C0(n9921), .Y(n9920)
         );
  AOI211XL U1868 ( .A0(n1621), .A1(n3231), .B0(n5811), .C0(n8169), .Y(n8168)
         );
  AOI211XL U1869 ( .A0(n1618), .A1(n3052), .B0(n5575), .C0(n9045), .Y(n9044)
         );
  AOI211XL U1870 ( .A0(n1614), .A1(n2811), .B0(n5255), .C0(n10213), .Y(n10212)
         );
  AOI211XL U1871 ( .A0(n1611), .A1(n2630), .B0(n4985), .C0(n11089), .Y(n11088)
         );
  AOI211XL U1872 ( .A0(n1612), .A1(n2698), .B0(n5069), .C0(n10797), .Y(n10796)
         );
  AOI211XL U1873 ( .A0(n1624), .A1(n3419), .B0(n6039), .C0(n7293), .Y(n7292)
         );
  AOI211XL U1874 ( .A0(n1617), .A1(n3001), .B0(n5499), .C0(n9337), .Y(n9336)
         );
  AOI211XL U1875 ( .A0(n1620), .A1(n3170), .B0(n5727), .C0(n8461), .Y(n8460)
         );
  AOI211XL U1876 ( .A0(n1623), .A1(n3353), .B0(n5963), .C0(n7585), .Y(n7584)
         );
  AOI211XL U1877 ( .A0(n1610), .A1(n2569), .B0(n4869), .C0(n11381), .Y(n11380)
         );
  AOI211XL U1878 ( .A0(n1613), .A1(n2750), .B0(n5177), .C0(n10505), .Y(n10504)
         );
  AOI211XL U1879 ( .A0(n1616), .A1(n2940), .B0(n5423), .C0(n9629), .Y(n9628)
         );
  AOI211XL U1880 ( .A0(n1619), .A1(n3113), .B0(n5651), .C0(n8753), .Y(n8752)
         );
  AOI211XL U1881 ( .A0(n1622), .A1(n3292), .B0(n5887), .C0(n7877), .Y(n7876)
         );
  AOI31XL U1882 ( .A0(n13561), .A1(n13562), .A2(n13563), .B0(n1638), .Y(n13560) );
  NAND3XL U1883 ( .A(n1258), .B(n1204), .C(n11849), .Y(n11851) );
  NAND3XL U1884 ( .A(n1330), .B(n1195), .C(top_core_KE_sb1_n278), .Y(
        top_core_KE_sb1_n280) );
  NAND3XL U1885 ( .A(n1265), .B(n1164), .C(n12480), .Y(n12482) );
  NAND3XL U1886 ( .A(n1261), .B(n1155), .C(n12165), .Y(n12167) );
  NAND3XL U1887 ( .A(n1268), .B(n1190), .C(n12795), .Y(n12797) );
  NAND3XL U1888 ( .A(n1277), .B(n1159), .C(n13740), .Y(n13742) );
  NAND3XL U1889 ( .A(n1271), .B(n1199), .C(n13110), .Y(n13112) );
  INVX1 U1890 ( .A(n_ADDR[1]), .Y(n4137) );
  CLKINVX3 U1891 ( .A(n4140), .Y(n4138) );
  CLKINVX3 U1892 ( .A(n4143), .Y(n4142) );
  NAND2X2 U1893 ( .A(top_core_io_n49), .B(n85), .Y(n266) );
  NOR4BXL U1894 ( .AN(n10010), .B(n993), .C(n5339), .D(n5365), .Y(n10009) );
  NOR4BXL U1895 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n196), .B(n1135), .C(
        n6135), .D(n6155), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n195) );
  NOR4BXL U1896 ( .AN(n11178), .B(n937), .C(n4985), .D(n5011), .Y(n11177) );
  NOR4BXL U1897 ( .AN(n8258), .B(n1077), .C(n5811), .D(n5837), .Y(n8257) );
  NOR4BXL U1898 ( .AN(n10886), .B(n951), .C(n5069), .D(n5095), .Y(n10885) );
  NOR4BXL U1899 ( .AN(n9134), .B(n1035), .C(n5575), .D(n5601), .Y(n9133) );
  NOR4BXL U1900 ( .AN(n7382), .B(n1119), .C(n6039), .D(n6065), .Y(n7381) );
  NOR4BXL U1901 ( .AN(n10302), .B(n979), .C(n5255), .D(n5281), .Y(n10301) );
  NOR4BXL U1902 ( .AN(n9426), .B(n1021), .C(n5499), .D(n5525), .Y(n9425) );
  NOR4BXL U1903 ( .AN(n8550), .B(n1063), .C(n5727), .D(n5753), .Y(n8549) );
  NOR4BXL U1904 ( .AN(n7674), .B(n1105), .C(n5963), .D(n5989), .Y(n7673) );
  NOR4BXL U1905 ( .AN(n11470), .B(n923), .C(n4869), .D(n4895), .Y(n11469) );
  NOR4BXL U1906 ( .AN(n10594), .B(n965), .C(n5177), .D(n5203), .Y(n10593) );
  NOR4BXL U1907 ( .AN(n9718), .B(n1007), .C(n5423), .D(n5449), .Y(n9717) );
  NOR4BXL U1908 ( .AN(n8842), .B(n1049), .C(n5651), .D(n5677), .Y(n8841) );
  NOR4BXL U1909 ( .AN(n7966), .B(n1091), .C(n5887), .D(n5913), .Y(n7965) );
  AND2X1 U1910 ( .A(n10497), .B(n1250), .Y(n333) );
  AND2X1 U1911 ( .A(n9329), .B(n1242), .Y(n329) );
  AND2X1 U1912 ( .A(n7577), .B(n1230), .Y(n331) );
  AND2X1 U1913 ( .A(n8745), .B(n1238), .Y(n335) );
  AND2X1 U1914 ( .A(n9913), .B(n1246), .Y(n321) );
  AND2X1 U1915 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .B(n1328), .Y(
        n322) );
  AND2X1 U1916 ( .A(n11081), .B(n1254), .Y(n323) );
  AND2X1 U1917 ( .A(n8161), .B(n1234), .Y(n324) );
  AND2X1 U1918 ( .A(n10789), .B(n1252), .Y(n325) );
  AND2X1 U1919 ( .A(n7285), .B(n1228), .Y(n326) );
  AND2X1 U1920 ( .A(n9037), .B(n1240), .Y(n327) );
  AND2X1 U1921 ( .A(n10205), .B(n1248), .Y(n328) );
  AND2X1 U1922 ( .A(n8453), .B(n1236), .Y(n330) );
  AND2X1 U1923 ( .A(n11373), .B(n1256), .Y(n332) );
  AND2X1 U1924 ( .A(n9621), .B(n1244), .Y(n334) );
  AND2X1 U1925 ( .A(n7869), .B(n1232), .Y(n336) );
  AOI21XL U1926 ( .A0(n9900), .A1(n5350), .B0(n9986), .Y(n10021) );
  AOI21XL U1927 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .A1(n6146), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n172), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n207) );
  AOI21XL U1928 ( .A0(n11068), .A1(n4996), .B0(n11154), .Y(n11189) );
  AOI21XL U1929 ( .A0(n8148), .A1(n5822), .B0(n8234), .Y(n8269) );
  AOI21XL U1930 ( .A0(n10776), .A1(n5080), .B0(n10862), .Y(n10897) );
  AOI21XL U1931 ( .A0(n9024), .A1(n5586), .B0(n9110), .Y(n9145) );
  AOI21XL U1932 ( .A0(n7272), .A1(n6050), .B0(n7358), .Y(n7393) );
  AOI21XL U1933 ( .A0(n10192), .A1(n5266), .B0(n10278), .Y(n10313) );
  AOI21XL U1934 ( .A0(n9316), .A1(n5510), .B0(n9402), .Y(n9437) );
  AOI21XL U1935 ( .A0(n8440), .A1(n5738), .B0(n8526), .Y(n8561) );
  AOI21XL U1936 ( .A0(n7564), .A1(n5974), .B0(n7650), .Y(n7685) );
  AOI21XL U1937 ( .A0(n11360), .A1(n4880), .B0(n11446), .Y(n11481) );
  AOI21XL U1938 ( .A0(n10484), .A1(n5188), .B0(n10570), .Y(n10605) );
  AOI21XL U1939 ( .A0(n9608), .A1(n5434), .B0(n9694), .Y(n9729) );
  AOI21XL U1940 ( .A0(n8732), .A1(n5662), .B0(n8818), .Y(n8853) );
  AOI21XL U1941 ( .A0(n7856), .A1(n5898), .B0(n7942), .Y(n7977) );
  AOI21XL U1942 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), .A1(n6137), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n198), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n91) );
  AOI21XL U1943 ( .A0(n9891), .A1(n5341), .B0(n10012), .Y(n9907) );
  AOI21XL U1944 ( .A0(n11059), .A1(n4987), .B0(n11180), .Y(n11075) );
  AOI21XL U1945 ( .A0(n8139), .A1(n5813), .B0(n8260), .Y(n8155) );
  AOI21XL U1946 ( .A0(n10767), .A1(n5071), .B0(n10888), .Y(n10783) );
  AOI21XL U1947 ( .A0(n7263), .A1(n6041), .B0(n7384), .Y(n7279) );
  AOI21XL U1948 ( .A0(n9015), .A1(n5577), .B0(n9136), .Y(n9031) );
  AOI21XL U1949 ( .A0(n10183), .A1(n5257), .B0(n10304), .Y(n10199) );
  AOI21XL U1950 ( .A0(n9307), .A1(n5501), .B0(n9428), .Y(n9323) );
  AOI21XL U1951 ( .A0(n8431), .A1(n5729), .B0(n8552), .Y(n8447) );
  AOI21XL U1952 ( .A0(n7555), .A1(n5965), .B0(n7676), .Y(n7571) );
  AOI21XL U1953 ( .A0(n11351), .A1(n4871), .B0(n11472), .Y(n11367) );
  AOI21XL U1954 ( .A0(n10475), .A1(n5179), .B0(n10596), .Y(n10491) );
  AOI21XL U1955 ( .A0(n9599), .A1(n5425), .B0(n9720), .Y(n9615) );
  AOI21XL U1956 ( .A0(n8723), .A1(n5653), .B0(n8844), .Y(n8739) );
  AOI21XL U1957 ( .A0(n7847), .A1(n5889), .B0(n7968), .Y(n7863) );
  AOI21XL U1958 ( .A0(n5350), .A1(n9970), .B0(n10012), .Y(n10046) );
  AOI21XL U1959 ( .A0(n6146), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n198), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n232) );
  AOI21XL U1960 ( .A0(n4996), .A1(n11138), .B0(n11180), .Y(n11214) );
  AOI21XL U1961 ( .A0(n5822), .A1(n8218), .B0(n8260), .Y(n8294) );
  AOI21XL U1962 ( .A0(n5080), .A1(n10846), .B0(n10888), .Y(n10922) );
  AOI21XL U1963 ( .A0(n5586), .A1(n9094), .B0(n9136), .Y(n9170) );
  AOI21XL U1964 ( .A0(n6050), .A1(n7342), .B0(n7384), .Y(n7418) );
  AOI21XL U1965 ( .A0(n5266), .A1(n10262), .B0(n10304), .Y(n10338) );
  AOI21XL U1966 ( .A0(n5510), .A1(n9386), .B0(n9428), .Y(n9462) );
  AOI21XL U1967 ( .A0(n5738), .A1(n8510), .B0(n8552), .Y(n8586) );
  AOI21XL U1968 ( .A0(n5974), .A1(n7634), .B0(n7676), .Y(n7710) );
  AOI21XL U1969 ( .A0(n4880), .A1(n11430), .B0(n11472), .Y(n11506) );
  AOI21XL U1970 ( .A0(n5188), .A1(n10554), .B0(n10596), .Y(n10630) );
  AOI21XL U1971 ( .A0(n5434), .A1(n9678), .B0(n9720), .Y(n9754) );
  AOI21XL U1972 ( .A0(n5662), .A1(n8802), .B0(n8844), .Y(n8878) );
  AOI21XL U1973 ( .A0(n5898), .A1(n7926), .B0(n7968), .Y(n8002) );
  AOI222XL U1974 ( .A0(n5341), .A1(n9891), .B0(n481), .B1(n993), .C0(n996), 
        .C1(n2881), .Y(n10002) );
  AOI222XL U1975 ( .A0(n6137), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), 
        .B0(n482), .B1(n1135), .C0(n1139), .C1(n3490), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n188) );
  AOI222XL U1976 ( .A0(n4987), .A1(n11059), .B0(n483), .B1(n937), .C0(n940), 
        .C1(n2639), .Y(n11170) );
  AOI222XL U1977 ( .A0(n5813), .A1(n8139), .B0(n484), .B1(n1077), .C0(n1080), 
        .C1(n3241), .Y(n8250) );
  AOI222XL U1978 ( .A0(n5071), .A1(n10767), .B0(n485), .B1(n951), .C0(n954), 
        .C1(n2700), .Y(n10878) );
  AOI222XL U1979 ( .A0(n5577), .A1(n9015), .B0(n486), .B1(n1035), .C0(n1038), 
        .C1(n3061), .Y(n9126) );
  AOI222XL U1980 ( .A0(n6041), .A1(n7263), .B0(n487), .B1(n1119), .C0(n1122), 
        .C1(n3421), .Y(n7374) );
  AOI222XL U1981 ( .A0(n5257), .A1(n10183), .B0(n488), .B1(n979), .C0(n982), 
        .C1(n2821), .Y(n10294) );
  AOI222XL U1982 ( .A0(n5501), .A1(n9307), .B0(n489), .B1(n1021), .C0(n1024), 
        .C1(n3003), .Y(n9418) );
  AOI222XL U1983 ( .A0(n5729), .A1(n8431), .B0(n490), .B1(n1063), .C0(n1066), 
        .C1(n3180), .Y(n8542) );
  AOI222XL U1984 ( .A0(n5965), .A1(n7555), .B0(n491), .B1(n1105), .C0(n1108), 
        .C1(n3363), .Y(n7666) );
  AOI222XL U1985 ( .A0(n4871), .A1(n11351), .B0(n492), .B1(n923), .C0(n926), 
        .C1(n2578), .Y(n11462) );
  AOI222XL U1986 ( .A0(n5179), .A1(n10475), .B0(n493), .B1(n965), .C0(n968), 
        .C1(n2760), .Y(n10586) );
  AOI222XL U1987 ( .A0(n5425), .A1(n9599), .B0(n494), .B1(n1007), .C0(n1010), 
        .C1(n2942), .Y(n9710) );
  AOI222XL U1988 ( .A0(n5653), .A1(n8723), .B0(n495), .B1(n1049), .C0(n1052), 
        .C1(n3122), .Y(n8834) );
  AOI222XL U1989 ( .A0(n5889), .A1(n7847), .B0(n496), .B1(n1091), .C0(n1094), 
        .C1(n3302), .Y(n7958) );
  NOR4BXL U1990 ( .AN(n9950), .B(n5372), .C(n10044), .D(n10064), .Y(n10063) );
  NOR4BXL U1991 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n135), .B(n6162), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n230), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n250), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n249) );
  NOR4BXL U1992 ( .AN(n11118), .B(n5018), .C(n11212), .D(n11232), .Y(n11231)
         );
  NOR4BXL U1993 ( .AN(n8198), .B(n5844), .C(n8292), .D(n8312), .Y(n8311) );
  NOR4BXL U1994 ( .AN(n10826), .B(n5102), .C(n10920), .D(n10940), .Y(n10939)
         );
  NOR4BXL U1995 ( .AN(n7322), .B(n6072), .C(n7416), .D(n7436), .Y(n7435) );
  NOR4BXL U1996 ( .AN(n9074), .B(n5608), .C(n9168), .D(n9188), .Y(n9187) );
  NOR4BXL U1997 ( .AN(n10242), .B(n5288), .C(n10336), .D(n10356), .Y(n10355)
         );
  NOR4BXL U1998 ( .AN(n9366), .B(n5532), .C(n9460), .D(n9480), .Y(n9479) );
  NOR4BXL U1999 ( .AN(n8490), .B(n5760), .C(n8584), .D(n8604), .Y(n8603) );
  NOR4BXL U2000 ( .AN(n7614), .B(n5996), .C(n7708), .D(n7728), .Y(n7727) );
  NOR4BXL U2001 ( .AN(n11410), .B(n4902), .C(n11504), .D(n11524), .Y(n11523)
         );
  NOR4BXL U2002 ( .AN(n10534), .B(n5210), .C(n10628), .D(n10648), .Y(n10647)
         );
  NOR4BXL U2003 ( .AN(n9658), .B(n5456), .C(n9752), .D(n9772), .Y(n9771) );
  NOR4BXL U2004 ( .AN(n8782), .B(n5684), .C(n8876), .D(n8896), .Y(n8895) );
  NOR4BXL U2005 ( .AN(n7906), .B(n5920), .C(n8000), .D(n8020), .Y(n8019) );
  AOI211XL U2006 ( .A0(n481), .A1(n586), .B0(n5345), .C0(n10038), .Y(n10072)
         );
  AOI211XL U2007 ( .A0(n482), .A1(n585), .B0(n6141), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n224), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n258) );
  AOI211XL U2008 ( .A0(n483), .A1(n587), .B0(n4991), .C0(n11206), .Y(n11240)
         );
  AOI211XL U2009 ( .A0(n484), .A1(n588), .B0(n5817), .C0(n8286), .Y(n8320) );
  AOI211XL U2010 ( .A0(n485), .A1(n589), .B0(n5075), .C0(n10914), .Y(n10948)
         );
  AOI211XL U2011 ( .A0(n487), .A1(n591), .B0(n6045), .C0(n7410), .Y(n7444) );
  AOI211XL U2012 ( .A0(n486), .A1(n590), .B0(n5581), .C0(n9162), .Y(n9196) );
  AOI211XL U2013 ( .A0(n488), .A1(n592), .B0(n5261), .C0(n10330), .Y(n10364)
         );
  AOI211XL U2014 ( .A0(n489), .A1(n593), .B0(n5505), .C0(n9454), .Y(n9488) );
  AOI211XL U2015 ( .A0(n490), .A1(n594), .B0(n5733), .C0(n8578), .Y(n8612) );
  AOI211XL U2016 ( .A0(n491), .A1(n595), .B0(n5969), .C0(n7702), .Y(n7736) );
  AOI211XL U2017 ( .A0(n492), .A1(n596), .B0(n4875), .C0(n11498), .Y(n11532)
         );
  AOI211XL U2018 ( .A0(n493), .A1(n597), .B0(n5183), .C0(n10622), .Y(n10656)
         );
  AOI211XL U2019 ( .A0(n494), .A1(n598), .B0(n5429), .C0(n9746), .Y(n9780) );
  AOI211XL U2020 ( .A0(n495), .A1(n599), .B0(n5657), .C0(n8870), .Y(n8904) );
  AOI211XL U2021 ( .A0(n496), .A1(n600), .B0(n5893), .C0(n7994), .Y(n8028) );
  NOR2XL U2022 ( .A(n10064), .B(n9921), .Y(n10117) );
  NOR2XL U2023 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n250), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n106), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n303) );
  NOR2XL U2024 ( .A(n8312), .B(n8169), .Y(n8365) );
  NOR2XL U2025 ( .A(n11232), .B(n11089), .Y(n11285) );
  NOR2XL U2026 ( .A(n10940), .B(n10797), .Y(n10993) );
  NOR2XL U2027 ( .A(n7436), .B(n7293), .Y(n7489) );
  NOR2XL U2028 ( .A(n9188), .B(n9045), .Y(n9241) );
  NOR2XL U2029 ( .A(n10356), .B(n10213), .Y(n10409) );
  NOR2XL U2030 ( .A(n9480), .B(n9337), .Y(n9533) );
  NOR2XL U2031 ( .A(n8604), .B(n8461), .Y(n8657) );
  NOR2XL U2032 ( .A(n7728), .B(n7585), .Y(n7781) );
  NOR2XL U2033 ( .A(n11524), .B(n11381), .Y(n11577) );
  NOR2XL U2034 ( .A(n10648), .B(n10505), .Y(n10701) );
  NOR2XL U2035 ( .A(n9772), .B(n9629), .Y(n9825) );
  NOR2XL U2036 ( .A(n8896), .B(n8753), .Y(n8949) );
  NOR2XL U2037 ( .A(n8020), .B(n7877), .Y(n8073) );
  AOI22XL U2038 ( .A0(n3492), .A1(n1136), .B0(n13857), .B1(n1133), .Y(n13896)
         );
  AOI22XL U2039 ( .A0(n2891), .A1(n997), .B0(n17007), .B1(n994), .Y(n17046) );
  AOI22XL U2040 ( .A0(n2649), .A1(n941), .B0(n18267), .B1(n938), .Y(n18306) );
  AOI22XL U2041 ( .A0(n3251), .A1(n1081), .B0(n15117), .B1(n1078), .Y(n15156)
         );
  AOI22XL U2042 ( .A0(n3183), .A1(n1067), .B0(n15432), .B1(n1064), .Y(n15471)
         );
  AOI22XL U2043 ( .A0(n2581), .A1(n927), .B0(n18582), .B1(n924), .Y(n18621) );
  AOI22XL U2044 ( .A0(n2952), .A1(n1011), .B0(n16692), .B1(n1008), .Y(n16731)
         );
  AOI22XL U2045 ( .A0(n3312), .A1(n1095), .B0(n14802), .B1(n1092), .Y(n14841)
         );
  AOI22XL U2046 ( .A0(n3013), .A1(n1025), .B0(n16377), .B1(n1022), .Y(n16416)
         );
  AOI22XL U2047 ( .A0(n2703), .A1(n955), .B0(n17952), .B1(n952), .Y(n17991) );
  AOI22XL U2048 ( .A0(n3366), .A1(n1109), .B0(n14487), .B1(n1106), .Y(n14526)
         );
  AOI22XL U2049 ( .A0(n3071), .A1(n1039), .B0(n16062), .B1(n1036), .Y(n16101)
         );
  AOI22XL U2050 ( .A0(n2763), .A1(n969), .B0(n17637), .B1(n966), .Y(n17676) );
  AOI22XL U2051 ( .A0(n3431), .A1(n1123), .B0(n14172), .B1(n1120), .Y(n14211)
         );
  AOI22XL U2052 ( .A0(n3125), .A1(n1053), .B0(n15747), .B1(n1050), .Y(n15786)
         );
  AOI22XL U2053 ( .A0(n2831), .A1(n983), .B0(n17322), .B1(n980), .Y(n17361) );
  AOI22XL U2054 ( .A0(n13867), .A1(n3474), .B0(n3472), .B1(n13897), .Y(n13868)
         );
  AOI22XL U2055 ( .A0(n5384), .A1(n9900), .B0(n5336), .B1(n2892), .Y(n10007)
         );
  AOI22XL U2056 ( .A0(n6169), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), 
        .B0(n6132), .B1(n3493), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n193) );
  AOI22XL U2057 ( .A0(n5030), .A1(n11068), .B0(n4982), .B1(n2651), .Y(n11175)
         );
  AOI22XL U2058 ( .A0(n5856), .A1(n8148), .B0(n5808), .B1(n3252), .Y(n8255) );
  AOI22XL U2059 ( .A0(n5114), .A1(n10776), .B0(n5066), .B1(n2710), .Y(n10883)
         );
  AOI22XL U2060 ( .A0(n5620), .A1(n9024), .B0(n5572), .B1(n3073), .Y(n9131) );
  AOI22XL U2061 ( .A0(n6084), .A1(n7272), .B0(n6036), .B1(n3432), .Y(n7379) );
  AOI22XL U2062 ( .A0(n5300), .A1(n10192), .B0(n5252), .B1(n2832), .Y(n10299)
         );
  AOI22XL U2063 ( .A0(n5544), .A1(n9316), .B0(n5496), .B1(n3014), .Y(n9423) );
  AOI22XL U2064 ( .A0(n5772), .A1(n8440), .B0(n5724), .B1(n3191), .Y(n8547) );
  AOI22XL U2065 ( .A0(n6008), .A1(n7564), .B0(n5960), .B1(n3374), .Y(n7671) );
  AOI22XL U2066 ( .A0(n4914), .A1(n11360), .B0(n4866), .B1(n2589), .Y(n11467)
         );
  AOI22XL U2067 ( .A0(n5222), .A1(n10484), .B0(n5174), .B1(n2771), .Y(n10591)
         );
  AOI22XL U2068 ( .A0(n5468), .A1(n9608), .B0(n5420), .B1(n2953), .Y(n9715) );
  AOI22XL U2069 ( .A0(n5696), .A1(n8732), .B0(n5648), .B1(n3133), .Y(n8839) );
  AOI22XL U2070 ( .A0(n5932), .A1(n7856), .B0(n5884), .B1(n3313), .Y(n7963) );
  AOI211XL U2071 ( .A0(n5383), .A1(n9913), .B0(n5339), .C0(n5342), .Y(n9959)
         );
  AOI211XL U2072 ( .A0(n6168), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n97), 
        .B0(n6135), .C0(n6138), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n144) );
  AOI211XL U2073 ( .A0(n5029), .A1(n11081), .B0(n4985), .C0(n4988), .Y(n11127)
         );
  AOI211XL U2074 ( .A0(n5855), .A1(n8161), .B0(n5811), .C0(n5814), .Y(n8207)
         );
  AOI211XL U2075 ( .A0(n5113), .A1(n10789), .B0(n5069), .C0(n5072), .Y(n10835)
         );
  AOI211XL U2076 ( .A0(n5619), .A1(n9037), .B0(n5575), .C0(n5578), .Y(n9083)
         );
  AOI211XL U2077 ( .A0(n6083), .A1(n7285), .B0(n6039), .C0(n6042), .Y(n7331)
         );
  AOI211XL U2078 ( .A0(n5299), .A1(n10205), .B0(n5255), .C0(n5258), .Y(n10251)
         );
  AOI211XL U2079 ( .A0(n5543), .A1(n9329), .B0(n5499), .C0(n5502), .Y(n9375)
         );
  AOI211XL U2080 ( .A0(n5771), .A1(n8453), .B0(n5727), .C0(n5730), .Y(n8499)
         );
  AOI211XL U2081 ( .A0(n6007), .A1(n7577), .B0(n5963), .C0(n5966), .Y(n7623)
         );
  AOI211XL U2082 ( .A0(n4913), .A1(n11373), .B0(n4869), .C0(n4872), .Y(n11419)
         );
  AOI211XL U2083 ( .A0(n5221), .A1(n10497), .B0(n5177), .C0(n5180), .Y(n10543)
         );
  AOI211XL U2084 ( .A0(n5467), .A1(n9621), .B0(n5423), .C0(n5426), .Y(n9667)
         );
  AOI211XL U2085 ( .A0(n5695), .A1(n8745), .B0(n5651), .C0(n5654), .Y(n8791)
         );
  AOI211XL U2086 ( .A0(n5931), .A1(n7869), .B0(n5887), .C0(n5890), .Y(n7915)
         );
  AOI222XL U2087 ( .A0(n1002), .A1(n5385), .B0(n17175), .B1(n2897), .C0(n5357), 
        .C1(n17047), .Y(n17204) );
  AOI222XL U2088 ( .A0(n1141), .A1(n6167), .B0(n14025), .B1(n3496), .C0(n6125), 
        .C1(n13897), .Y(n14054) );
  AOI222XL U2089 ( .A0(n946), .A1(n5031), .B0(n18435), .B1(n2658), .C0(n5003), 
        .C1(n18307), .Y(n18464) );
  AOI222XL U2090 ( .A0(n1086), .A1(n5857), .B0(n15285), .B1(n3257), .C0(n5829), 
        .C1(n15157), .Y(n15314) );
  AOI222XL U2091 ( .A0(n1072), .A1(n5773), .B0(n15600), .B1(n3196), .C0(n5745), 
        .C1(n15472), .Y(n15629) );
  AOI222XL U2092 ( .A0(n1016), .A1(n5469), .B0(n16860), .B1(n2958), .C0(n5441), 
        .C1(n16732), .Y(n16889) );
  AOI222XL U2093 ( .A0(n932), .A1(n4915), .B0(n18750), .B1(n2597), .C0(n4887), 
        .C1(n18622), .Y(n18779) );
  AOI222XL U2094 ( .A0(n1100), .A1(n5933), .B0(n14970), .B1(n3317), .C0(n5905), 
        .C1(n14842), .Y(n14999) );
  AOI222XL U2095 ( .A0(n1030), .A1(n5545), .B0(n16545), .B1(n3022), .C0(n5517), 
        .C1(n16417), .Y(n16574) );
  AOI222XL U2096 ( .A0(n960), .A1(n5115), .B0(n18120), .B1(n2716), .C0(n5087), 
        .C1(n17992), .Y(n18149) );
  AOI222XL U2097 ( .A0(n1114), .A1(n6009), .B0(n14655), .B1(n3382), .C0(n5981), 
        .C1(n14527), .Y(n14684) );
  AOI222XL U2098 ( .A0(n1044), .A1(n5621), .B0(n16230), .B1(n3080), .C0(n5593), 
        .C1(n16102), .Y(n16259) );
  AOI222XL U2099 ( .A0(n974), .A1(n5223), .B0(n17805), .B1(n2782), .C0(n5195), 
        .C1(n17677), .Y(n17834) );
  AOI222XL U2100 ( .A0(n1128), .A1(n6085), .B0(n14340), .B1(n3438), .C0(n6057), 
        .C1(n14212), .Y(n14369) );
  AOI222XL U2101 ( .A0(n1058), .A1(n5697), .B0(n15915), .B1(n3141), .C0(n5669), 
        .C1(n15787), .Y(n15944) );
  AOI222XL U2102 ( .A0(n988), .A1(n5301), .B0(n17490), .B1(n2835), .C0(n5273), 
        .C1(n17362), .Y(n17519) );
  AOI222XL U2103 ( .A0(n6137), .A1(n1327), .B0(n6169), .B1(n530), .C0(n6146), 
        .C1(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n316) );
  AOI2BB1XL U2104 ( .A0N(n3497), .A1N(top_core_EC_ss_gen_tbox_0__sboxs_r_n255), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n287), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n315) );
  AOI222XL U2105 ( .A0(n5341), .A1(n1245), .B0(n5384), .B1(n529), .C0(n5350), 
        .C1(n9970), .Y(n10130) );
  AOI2BB1XL U2106 ( .A0N(n2904), .A1N(n10069), .B0(n10101), .Y(n10129) );
  AOI222XL U2107 ( .A0(n4987), .A1(n1253), .B0(n5030), .B1(n531), .C0(n4996), 
        .C1(n11138), .Y(n11298) );
  AOI2BB1XL U2108 ( .A0N(n2658), .A1N(n11237), .B0(n11269), .Y(n11297) );
  AOI222XL U2109 ( .A0(n5813), .A1(n1233), .B0(n5856), .B1(n532), .C0(n5822), 
        .C1(n8218), .Y(n8378) );
  AOI2BB1XL U2110 ( .A0N(n3264), .A1N(n8317), .B0(n8349), .Y(n8377) );
  AOI222XL U2111 ( .A0(n5071), .A1(n1251), .B0(n5114), .B1(n533), .C0(n5080), 
        .C1(n10846), .Y(n11006) );
  AOI2BB1XL U2112 ( .A0N(n2714), .A1N(n10945), .B0(n10977), .Y(n11005) );
  AOI222XL U2113 ( .A0(n5577), .A1(n1239), .B0(n5620), .B1(n534), .C0(n5586), 
        .C1(n9094), .Y(n9254) );
  AOI2BB1XL U2114 ( .A0N(n3080), .A1N(n9193), .B0(n9225), .Y(n9253) );
  AOI222XL U2115 ( .A0(n6041), .A1(n1227), .B0(n6084), .B1(n535), .C0(n6050), 
        .C1(n7342), .Y(n7502) );
  AOI2BB1XL U2116 ( .A0N(n3436), .A1N(n7441), .B0(n7473), .Y(n7501) );
  AOI222XL U2117 ( .A0(n5257), .A1(n1247), .B0(n5300), .B1(n536), .C0(n5266), 
        .C1(n10262), .Y(n10422) );
  AOI2BB1XL U2118 ( .A0N(n2837), .A1N(n10361), .B0(n10393), .Y(n10421) );
  AOI222XL U2119 ( .A0(n5501), .A1(n1241), .B0(n5544), .B1(n537), .C0(n5510), 
        .C1(n9386), .Y(n9546) );
  AOI2BB1XL U2120 ( .A0N(n3025), .A1N(n9485), .B0(n9517), .Y(n9545) );
  AOI222XL U2121 ( .A0(n5729), .A1(n1235), .B0(n5772), .B1(n538), .C0(n5738), 
        .C1(n8510), .Y(n8670) );
  AOI2BB1XL U2122 ( .A0N(n3203), .A1N(n8609), .B0(n8641), .Y(n8669) );
  AOI222XL U2123 ( .A0(n5965), .A1(n1229), .B0(n6008), .B1(n539), .C0(n5974), 
        .C1(n7634), .Y(n7794) );
  AOI2BB1XL U2124 ( .A0N(n3385), .A1N(n7733), .B0(n7765), .Y(n7793) );
  AOI222XL U2125 ( .A0(n4871), .A1(n1255), .B0(n4914), .B1(n540), .C0(n4880), 
        .C1(n11430), .Y(n11590) );
  AOI2BB1XL U2126 ( .A0N(n2597), .A1N(n11529), .B0(n11561), .Y(n11589) );
  AOI222XL U2127 ( .A0(n5179), .A1(n1249), .B0(n5222), .B1(n541), .C0(n5188), 
        .C1(n10554), .Y(n10714) );
  AOI2BB1XL U2128 ( .A0N(n2782), .A1N(n10653), .B0(n10685), .Y(n10713) );
  AOI222XL U2129 ( .A0(n5425), .A1(n1243), .B0(n5468), .B1(n542), .C0(n5434), 
        .C1(n9678), .Y(n9838) );
  AOI2BB1XL U2130 ( .A0N(n2965), .A1N(n9777), .B0(n9809), .Y(n9837) );
  AOI222XL U2131 ( .A0(n5653), .A1(n1237), .B0(n5696), .B1(n543), .C0(n5662), 
        .C1(n8802), .Y(n8962) );
  AOI2BB1XL U2132 ( .A0N(n3144), .A1N(n8901), .B0(n8933), .Y(n8961) );
  AOI222XL U2133 ( .A0(n5889), .A1(n1231), .B0(n5932), .B1(n544), .C0(n5898), 
        .C1(n7926), .Y(n8086) );
  AOI2BB1XL U2134 ( .A0N(n3320), .A1N(n8025), .B0(n8057), .Y(n8085) );
  AOI22XL U2135 ( .A0(n5375), .A1(n9913), .B0(n1245), .B1(n2871), .Y(n9975) );
  AOI22XL U2136 ( .A0(n6165), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n97), 
        .B0(n1327), .B1(n3472), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n161) );
  AOI22XL U2137 ( .A0(n5021), .A1(n11081), .B0(n1253), .B1(n2629), .Y(n11143)
         );
  AOI22XL U2138 ( .A0(n5847), .A1(n8161), .B0(n1233), .B1(n3231), .Y(n8223) );
  AOI22XL U2139 ( .A0(n5105), .A1(n10789), .B0(n1251), .B1(n2690), .Y(n10851)
         );
  AOI22XL U2140 ( .A0(n5611), .A1(n9037), .B0(n1239), .B1(n3051), .Y(n9099) );
  AOI22XL U2141 ( .A0(n6075), .A1(n7285), .B0(n1227), .B1(n3411), .Y(n7347) );
  AOI22XL U2142 ( .A0(n5291), .A1(n10205), .B0(n1247), .B1(n2811), .Y(n10267)
         );
  AOI22XL U2143 ( .A0(n5535), .A1(n9329), .B0(n1241), .B1(n2993), .Y(n9391) );
  AOI22XL U2144 ( .A0(n5763), .A1(n8453), .B0(n1235), .B1(n3170), .Y(n8515) );
  AOI22XL U2145 ( .A0(n5999), .A1(n7577), .B0(n1229), .B1(n3353), .Y(n7639) );
  AOI22XL U2146 ( .A0(n4905), .A1(n11373), .B0(n1255), .B1(n2568), .Y(n11435)
         );
  AOI22XL U2147 ( .A0(n5213), .A1(n10497), .B0(n1249), .B1(n2750), .Y(n10559)
         );
  AOI22XL U2148 ( .A0(n5459), .A1(n9621), .B0(n1243), .B1(n2932), .Y(n9683) );
  AOI22XL U2149 ( .A0(n5687), .A1(n8745), .B0(n1237), .B1(n3112), .Y(n8807) );
  AOI22XL U2150 ( .A0(n5923), .A1(n7869), .B0(n1231), .B1(n3292), .Y(n7931) );
  NOR4BXL U2151 ( .AN(n9993), .B(n9994), .C(n9903), .D(n9995), .Y(n9991) );
  AOI22XL U2152 ( .A0(n353), .A1(n9996), .B0(n5350), .B1(n2900), .Y(n9993) );
  NOR4BXL U2153 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n179), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n180), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n86), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n181), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n177) );
  AOI22XL U2154 ( .A0(n354), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n182), 
        .B0(n6146), .B1(n3507), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n179) );
  NOR4BXL U2155 ( .AN(n11161), .B(n11162), .C(n11071), .D(n11163), .Y(n11159)
         );
  AOI22XL U2156 ( .A0(n356), .A1(n11164), .B0(n4996), .B1(n2664), .Y(n11161)
         );
  NOR4BXL U2157 ( .AN(n8241), .B(n8242), .C(n8151), .D(n8243), .Y(n8239) );
  AOI22XL U2158 ( .A0(n355), .A1(n8244), .B0(n5822), .B1(n3260), .Y(n8241) );
  NOR4BXL U2159 ( .AN(n10869), .B(n10870), .C(n10779), .D(n10871), .Y(n10867)
         );
  AOI22XL U2160 ( .A0(n357), .A1(n10872), .B0(n5080), .B1(n2713), .Y(n10869)
         );
  NOR4BXL U2161 ( .AN(n9117), .B(n9118), .C(n9027), .D(n9119), .Y(n9115) );
  AOI22XL U2162 ( .A0(n359), .A1(n9120), .B0(n5586), .B1(n3086), .Y(n9117) );
  NOR4BXL U2163 ( .AN(n7365), .B(n7366), .C(n7275), .D(n7367), .Y(n7363) );
  AOI22XL U2164 ( .A0(n358), .A1(n7368), .B0(n6050), .B1(n3435), .Y(n7365) );
  NOR4BXL U2165 ( .AN(n10285), .B(n10286), .C(n10195), .D(n10287), .Y(n10283)
         );
  AOI22XL U2166 ( .A0(n360), .A1(n10288), .B0(n5266), .B1(n2837), .Y(n10285)
         );
  NOR4BXL U2167 ( .AN(n9409), .B(n9410), .C(n9319), .D(n9411), .Y(n9407) );
  AOI22XL U2168 ( .A0(n361), .A1(n9412), .B0(n5510), .B1(n3018), .Y(n9409) );
  NOR4BXL U2169 ( .AN(n8533), .B(n8534), .C(n8443), .D(n8535), .Y(n8531) );
  AOI22XL U2170 ( .A0(n362), .A1(n8536), .B0(n5738), .B1(n3199), .Y(n8533) );
  NOR4BXL U2171 ( .AN(n7657), .B(n7658), .C(n7567), .D(n7659), .Y(n7655) );
  AOI22XL U2172 ( .A0(n363), .A1(n7660), .B0(n5974), .B1(n3378), .Y(n7657) );
  NOR4BXL U2173 ( .AN(n11453), .B(n11454), .C(n11363), .D(n11455), .Y(n11451)
         );
  AOI22XL U2174 ( .A0(n364), .A1(n11456), .B0(n4880), .B1(n2603), .Y(n11453)
         );
  NOR4BXL U2175 ( .AN(n10577), .B(n10578), .C(n10487), .D(n10579), .Y(n10575)
         );
  AOI22XL U2176 ( .A0(n365), .A1(n10580), .B0(n5188), .B1(n2776), .Y(n10577)
         );
  NOR4BXL U2177 ( .AN(n9701), .B(n9702), .C(n9611), .D(n9703), .Y(n9699) );
  AOI22XL U2178 ( .A0(n366), .A1(n9704), .B0(n5434), .B1(n2961), .Y(n9701) );
  NOR4BXL U2179 ( .AN(n8825), .B(n8826), .C(n8735), .D(n8827), .Y(n8823) );
  AOI22XL U2180 ( .A0(n367), .A1(n8828), .B0(n5662), .B1(n3137), .Y(n8825) );
  NOR4BXL U2181 ( .AN(n7949), .B(n7950), .C(n7859), .D(n7951), .Y(n7947) );
  AOI22XL U2182 ( .A0(n368), .A1(n7952), .B0(n5898), .B1(n3317), .Y(n7949) );
  AOI21XL U2183 ( .A0(n11430), .A1(n4908), .B0(n18633), .Y(n18868) );
  AOI21XL U2184 ( .A0(n7926), .A1(n5926), .B0(n14853), .Y(n15088) );
  AOI21XL U2185 ( .A0(n9094), .A1(n5614), .B0(n16113), .Y(n16348) );
  AOI21XL U2186 ( .A0(n10262), .A1(n5294), .B0(n17373), .Y(n17608) );
  AOI21XL U2187 ( .A0(n8510), .A1(n5766), .B0(n15483), .Y(n15718) );
  AOI21XL U2188 ( .A0(n10846), .A1(n5108), .B0(n18003), .Y(n18238) );
  AOI21XL U2189 ( .A0(n7342), .A1(n6078), .B0(n14223), .Y(n14458) );
  AOI21XL U2190 ( .A0(n9970), .A1(n5378), .B0(n17058), .Y(n17293) );
  AOI21XL U2191 ( .A0(n8218), .A1(n5850), .B0(n15168), .Y(n15403) );
  AOI21XL U2192 ( .A0(n11138), .A1(n5024), .B0(n18318), .Y(n18553) );
  AOI21XL U2193 ( .A0(n9678), .A1(n5462), .B0(n16743), .Y(n16978) );
  AOI21XL U2194 ( .A0(n9386), .A1(n5538), .B0(n16428), .Y(n16663) );
  AOI21XL U2195 ( .A0(n7634), .A1(n6002), .B0(n14538), .Y(n14773) );
  AOI21XL U2196 ( .A0(n10554), .A1(n5216), .B0(n17688), .Y(n17923) );
  AOI21XL U2197 ( .A0(n8802), .A1(n5690), .B0(n15798), .Y(n16033) );
  AOI21XL U2198 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .A1(n6149), 
        .B0(n13908), .Y(n14143) );
  AOI222XL U2199 ( .A0(n18649), .A1(n638), .B0(n924), .B1(n374), .C0(n928), 
        .C1(n1325), .Y(n18761) );
  AOI222XL U2200 ( .A0(n16129), .A1(n644), .B0(n1036), .B1(n380), .C0(n1040), 
        .C1(n1301), .Y(n16241) );
  AOI222XL U2201 ( .A0(n17389), .A1(n648), .B0(n980), .B1(n384), .C0(n984), 
        .C1(n1313), .Y(n17501) );
  AOI222XL U2202 ( .A0(n18019), .A1(n642), .B0(n952), .B1(n378), .C0(n956), 
        .C1(n1319), .Y(n18131) );
  AOI222XL U2203 ( .A0(n14239), .A1(n646), .B0(n1120), .B1(n382), .C0(n1124), 
        .C1(n1283), .Y(n14351) );
  AOI222XL U2204 ( .A0(n14869), .A1(n640), .B0(n1092), .B1(n376), .C0(n1096), 
        .C1(n1289), .Y(n14981) );
  AOI222XL U2205 ( .A0(n15499), .A1(n637), .B0(n1064), .B1(n373), .C0(n1068), 
        .C1(n1295), .Y(n15611) );
  AOI222XL U2206 ( .A0(n17074), .A1(n633), .B0(n994), .B1(n370), .C0(n998), 
        .C1(n1310), .Y(n17186) );
  AOI222XL U2207 ( .A0(n13924), .A1(n634), .B0(n1133), .B1(n369), .C0(n1137), 
        .C1(n1280), .Y(n14036) );
  AOI222XL U2208 ( .A0(n18334), .A1(n635), .B0(n938), .B1(n371), .C0(n942), 
        .C1(n1322), .Y(n18446) );
  AOI222XL U2209 ( .A0(n15184), .A1(n636), .B0(n1078), .B1(n372), .C0(n1082), 
        .C1(n1292), .Y(n15296) );
  AOI222XL U2210 ( .A0(n16759), .A1(n639), .B0(n1008), .B1(n375), .C0(n1012), 
        .C1(n1307), .Y(n16871) );
  AOI222XL U2211 ( .A0(n16444), .A1(n641), .B0(n1022), .B1(n377), .C0(n1026), 
        .C1(n1304), .Y(n16556) );
  AOI222XL U2212 ( .A0(n14554), .A1(n643), .B0(n1106), .B1(n379), .C0(n1110), 
        .C1(n1286), .Y(n14666) );
  AOI222XL U2213 ( .A0(n17704), .A1(n645), .B0(n966), .B1(n381), .C0(n970), 
        .C1(n1316), .Y(n17816) );
  AOI222XL U2214 ( .A0(n15814), .A1(n647), .B0(n1050), .B1(n383), .C0(n1054), 
        .C1(n1298), .Y(n15926) );
  NAND2XL U2215 ( .A(n17195), .B(n1311), .Y(n17085) );
  NAND2XL U2216 ( .A(n14045), .B(n1281), .Y(n13935) );
  NAND2XL U2217 ( .A(n15305), .B(n1293), .Y(n15195) );
  NAND2XL U2218 ( .A(n18455), .B(n1323), .Y(n18345) );
  NAND2XL U2219 ( .A(n15620), .B(n1296), .Y(n15510) );
  NAND2XL U2220 ( .A(n16880), .B(n1308), .Y(n16770) );
  NAND2XL U2221 ( .A(n18770), .B(n1326), .Y(n18660) );
  NAND2XL U2222 ( .A(n14990), .B(n1290), .Y(n14880) );
  NAND2XL U2223 ( .A(n16565), .B(n1305), .Y(n16455) );
  NAND2XL U2224 ( .A(n18140), .B(n1320), .Y(n18030) );
  NAND2XL U2225 ( .A(n14675), .B(n1287), .Y(n14565) );
  NAND2XL U2226 ( .A(n16250), .B(n1302), .Y(n16140) );
  NAND2XL U2227 ( .A(n17825), .B(n1317), .Y(n17715) );
  NAND2XL U2228 ( .A(n14360), .B(n1284), .Y(n14250) );
  NAND2XL U2229 ( .A(n15935), .B(n1299), .Y(n15825) );
  NAND2XL U2230 ( .A(n17510), .B(n1314), .Y(n17400) );
  OAI211XL U2231 ( .A0(n2881), .A1(n57), .B0(n17091), .C0(n17220), .Y(n17236)
         );
  OAI211XL U2232 ( .A0(n3482), .A1(n58), .B0(n13941), .C0(n14070), .Y(n14086)
         );
  OAI211XL U2233 ( .A0(n3241), .A1(n60), .B0(n15201), .C0(n15330), .Y(n15346)
         );
  OAI211XL U2234 ( .A0(n2639), .A1(n59), .B0(n18351), .C0(n18480), .Y(n18496)
         );
  OAI211XL U2235 ( .A0(n3180), .A1(n61), .B0(n15516), .C0(n15645), .Y(n15661)
         );
  OAI211XL U2236 ( .A0(n2942), .A1(n62), .B0(n16776), .C0(n16905), .Y(n16921)
         );
  OAI211XL U2237 ( .A0(n2578), .A1(n63), .B0(n18666), .C0(n18795), .Y(n18811)
         );
  OAI211XL U2238 ( .A0(n3302), .A1(n64), .B0(n14886), .C0(n15015), .Y(n15031)
         );
  OAI211XL U2239 ( .A0(n3003), .A1(n65), .B0(n16461), .C0(n16590), .Y(n16606)
         );
  OAI211XL U2240 ( .A0(n2700), .A1(n66), .B0(n18036), .C0(n18165), .Y(n18181)
         );
  OAI211XL U2241 ( .A0(n3363), .A1(n67), .B0(n14571), .C0(n14700), .Y(n14716)
         );
  OAI211XL U2242 ( .A0(n3061), .A1(n68), .B0(n16146), .C0(n16275), .Y(n16291)
         );
  OAI211XL U2243 ( .A0(n2760), .A1(n69), .B0(n17721), .C0(n17850), .Y(n17866)
         );
  OAI211XL U2244 ( .A0(n3421), .A1(n70), .B0(n14256), .C0(n14385), .Y(n14401)
         );
  OAI211XL U2245 ( .A0(n3122), .A1(n71), .B0(n15831), .C0(n15960), .Y(n15976)
         );
  OAI211XL U2246 ( .A0(n2821), .A1(n72), .B0(n17406), .C0(n17535), .Y(n17551)
         );
  NAND3XL U2247 ( .A(n10013), .B(n9956), .C(n9948), .Y(n10104) );
  NAND3XL U2248 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n199), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n141), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n133), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n290) );
  NAND3XL U2249 ( .A(n8261), .B(n8204), .C(n8196), .Y(n8352) );
  NAND3XL U2250 ( .A(n11181), .B(n11124), .C(n11116), .Y(n11272) );
  NAND3XL U2251 ( .A(n10889), .B(n10832), .C(n10824), .Y(n10980) );
  NAND3XL U2252 ( .A(n7385), .B(n7328), .C(n7320), .Y(n7476) );
  NAND3XL U2253 ( .A(n9137), .B(n9080), .C(n9072), .Y(n9228) );
  NAND3XL U2254 ( .A(n10305), .B(n10248), .C(n10240), .Y(n10396) );
  NAND3XL U2255 ( .A(n9429), .B(n9372), .C(n9364), .Y(n9520) );
  NAND3XL U2256 ( .A(n8553), .B(n8496), .C(n8488), .Y(n8644) );
  NAND3XL U2257 ( .A(n7677), .B(n7620), .C(n7612), .Y(n7768) );
  NAND3XL U2258 ( .A(n11473), .B(n11416), .C(n11408), .Y(n11564) );
  NAND3XL U2259 ( .A(n10597), .B(n10540), .C(n10532), .Y(n10688) );
  NAND3XL U2260 ( .A(n9721), .B(n9664), .C(n9656), .Y(n9812) );
  NAND3XL U2261 ( .A(n8845), .B(n8788), .C(n8780), .Y(n8936) );
  NAND3XL U2262 ( .A(n7969), .B(n7912), .C(n7904), .Y(n8060) );
  AOI22XL U2263 ( .A0(n5384), .A1(n401), .B0(n5336), .B1(n1245), .Y(n9962) );
  AOI22XL U2264 ( .A0(n6169), .A1(n402), .B0(n6132), .B1(n1327), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n147) );
  AOI22XL U2265 ( .A0(n5030), .A1(n403), .B0(n4982), .B1(n1253), .Y(n11130) );
  AOI22XL U2266 ( .A0(n5856), .A1(n404), .B0(n5808), .B1(n1233), .Y(n8210) );
  AOI22XL U2267 ( .A0(n5114), .A1(n405), .B0(n5066), .B1(n1251), .Y(n10838) );
  AOI22XL U2268 ( .A0(n5620), .A1(n406), .B0(n5572), .B1(n1239), .Y(n9086) );
  AOI22XL U2269 ( .A0(n6084), .A1(n407), .B0(n6036), .B1(n1227), .Y(n7334) );
  AOI22XL U2270 ( .A0(n5300), .A1(n408), .B0(n5252), .B1(n1247), .Y(n10254) );
  AOI22XL U2271 ( .A0(n5544), .A1(n409), .B0(n5496), .B1(n1241), .Y(n9378) );
  AOI22XL U2272 ( .A0(n5772), .A1(n410), .B0(n5724), .B1(n1235), .Y(n8502) );
  AOI22XL U2273 ( .A0(n6008), .A1(n411), .B0(n5960), .B1(n1229), .Y(n7626) );
  AOI22XL U2274 ( .A0(n4914), .A1(n412), .B0(n4866), .B1(n1255), .Y(n11422) );
  AOI22XL U2275 ( .A0(n5222), .A1(n413), .B0(n5174), .B1(n1249), .Y(n10546) );
  AOI22XL U2276 ( .A0(n5468), .A1(n414), .B0(n5420), .B1(n1243), .Y(n9670) );
  AOI22XL U2277 ( .A0(n5696), .A1(n415), .B0(n5648), .B1(n1237), .Y(n8794) );
  AOI22XL U2278 ( .A0(n5932), .A1(n416), .B0(n5884), .B1(n1231), .Y(n7918) );
  AOI21XL U2279 ( .A0(n17061), .A1(n5380), .B0(n17098), .Y(n17219) );
  AOI21XL U2280 ( .A0(n13911), .A1(n6151), .B0(n13948), .Y(n14069) );
  AOI21XL U2281 ( .A0(n15171), .A1(n5852), .B0(n15208), .Y(n15329) );
  AOI21XL U2282 ( .A0(n18321), .A1(n5026), .B0(n18358), .Y(n18479) );
  AOI21XL U2283 ( .A0(n15486), .A1(n5768), .B0(n15523), .Y(n15644) );
  AOI21XL U2284 ( .A0(n16746), .A1(n5464), .B0(n16783), .Y(n16904) );
  AOI21XL U2285 ( .A0(n18636), .A1(n4910), .B0(n18673), .Y(n18794) );
  AOI21XL U2286 ( .A0(n14856), .A1(n5928), .B0(n14893), .Y(n15014) );
  AOI21XL U2287 ( .A0(n16431), .A1(n5540), .B0(n16468), .Y(n16589) );
  AOI21XL U2288 ( .A0(n18006), .A1(n5110), .B0(n18043), .Y(n18164) );
  AOI21XL U2289 ( .A0(n14541), .A1(n6004), .B0(n14578), .Y(n14699) );
  AOI21XL U2290 ( .A0(n16116), .A1(n5616), .B0(n16153), .Y(n16274) );
  AOI21XL U2291 ( .A0(n17691), .A1(n5218), .B0(n17728), .Y(n17849) );
  AOI21XL U2292 ( .A0(n14226), .A1(n6080), .B0(n14263), .Y(n14384) );
  AOI21XL U2293 ( .A0(n15801), .A1(n5692), .B0(n15838), .Y(n15959) );
  AOI21XL U2294 ( .A0(n17376), .A1(n5296), .B0(n17413), .Y(n17534) );
  AOI21XL U2295 ( .A0(n5384), .A1(n450), .B0(n10038), .Y(n10036) );
  AOI21XL U2296 ( .A0(n6169), .A1(n449), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n224), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n222) );
  AOI21XL U2297 ( .A0(n5030), .A1(n451), .B0(n11206), .Y(n11204) );
  AOI21XL U2298 ( .A0(n5856), .A1(n452), .B0(n8286), .Y(n8284) );
  AOI21XL U2299 ( .A0(n5114), .A1(n458), .B0(n10914), .Y(n10912) );
  AOI21XL U2300 ( .A0(n5620), .A1(n460), .B0(n9162), .Y(n9160) );
  AOI21XL U2301 ( .A0(n6084), .A1(n462), .B0(n7410), .Y(n7408) );
  AOI21XL U2302 ( .A0(n5300), .A1(n464), .B0(n10330), .Y(n10328) );
  AOI21XL U2303 ( .A0(n5544), .A1(n457), .B0(n9454), .Y(n9452) );
  AOI21XL U2304 ( .A0(n5772), .A1(n453), .B0(n8578), .Y(n8576) );
  AOI21XL U2305 ( .A0(n6008), .A1(n459), .B0(n7702), .Y(n7700) );
  AOI21XL U2306 ( .A0(n4914), .A1(n454), .B0(n11498), .Y(n11496) );
  AOI21XL U2307 ( .A0(n5222), .A1(n461), .B0(n10622), .Y(n10620) );
  AOI21XL U2308 ( .A0(n5468), .A1(n455), .B0(n9746), .Y(n9744) );
  AOI21XL U2309 ( .A0(n5696), .A1(n463), .B0(n8870), .Y(n8868) );
  AOI21XL U2310 ( .A0(n5932), .A1(n456), .B0(n7994), .Y(n7992) );
  AOI21XL U2311 ( .A0(n5380), .A1(n17007), .B0(n5361), .Y(n17199) );
  AOI21XL U2312 ( .A0(n6151), .A1(n13857), .B0(n6129), .Y(n14049) );
  AOI21XL U2313 ( .A0(n5026), .A1(n18267), .B0(n5007), .Y(n18459) );
  AOI21XL U2314 ( .A0(n5852), .A1(n15117), .B0(n5833), .Y(n15309) );
  AOI21XL U2315 ( .A0(n5768), .A1(n15432), .B0(n5749), .Y(n15624) );
  AOI21XL U2316 ( .A0(n5464), .A1(n16692), .B0(n5445), .Y(n16884) );
  AOI21XL U2317 ( .A0(n4910), .A1(n18582), .B0(n4891), .Y(n18774) );
  AOI21XL U2318 ( .A0(n5928), .A1(n14802), .B0(n5909), .Y(n14994) );
  AOI21XL U2319 ( .A0(n5540), .A1(n16377), .B0(n5521), .Y(n16569) );
  AOI21XL U2320 ( .A0(n5110), .A1(n17952), .B0(n5091), .Y(n18144) );
  AOI21XL U2321 ( .A0(n6004), .A1(n14487), .B0(n5985), .Y(n14679) );
  AOI21XL U2322 ( .A0(n5616), .A1(n16062), .B0(n5597), .Y(n16254) );
  AOI21XL U2323 ( .A0(n5218), .A1(n17637), .B0(n5199), .Y(n17829) );
  AOI21XL U2324 ( .A0(n6080), .A1(n14172), .B0(n6061), .Y(n14364) );
  AOI21XL U2325 ( .A0(n5692), .A1(n15747), .B0(n5673), .Y(n15939) );
  AOI21XL U2326 ( .A0(n5296), .A1(n17322), .B0(n5277), .Y(n17514) );
  AOI222XL U2327 ( .A0(n586), .A1(n2896), .B0(n5384), .B1(n1245), .C0(n5350), 
        .C1(n529), .Y(n10015) );
  AOI222XL U2328 ( .A0(n585), .A1(n3496), .B0(n6169), .B1(n1327), .C0(n6146), 
        .C1(n530), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n201) );
  AOI222XL U2329 ( .A0(n587), .A1(n2653), .B0(n5030), .B1(n1253), .C0(n4996), 
        .C1(n531), .Y(n11183) );
  AOI222XL U2330 ( .A0(n588), .A1(n3256), .B0(n5856), .B1(n1233), .C0(n5822), 
        .C1(n532), .Y(n8263) );
  AOI222XL U2331 ( .A0(n589), .A1(n2719), .B0(n5114), .B1(n1251), .C0(n5080), 
        .C1(n533), .Y(n10891) );
  AOI222XL U2332 ( .A0(n590), .A1(n3075), .B0(n5620), .B1(n1239), .C0(n5586), 
        .C1(n534), .Y(n9139) );
  AOI222XL U2333 ( .A0(n591), .A1(n3441), .B0(n6084), .B1(n1227), .C0(n6050), 
        .C1(n535), .Y(n7387) );
  AOI222XL U2334 ( .A0(n592), .A1(n2841), .B0(n5300), .B1(n1247), .C0(n5266), 
        .C1(n536), .Y(n10307) );
  AOI222XL U2335 ( .A0(n593), .A1(n3020), .B0(n5544), .B1(n1241), .C0(n5510), 
        .C1(n537), .Y(n9431) );
  AOI222XL U2336 ( .A0(n594), .A1(n3195), .B0(n5772), .B1(n1235), .C0(n5738), 
        .C1(n538), .Y(n8555) );
  AOI222XL U2337 ( .A0(n595), .A1(n3380), .B0(n6008), .B1(n1229), .C0(n5974), 
        .C1(n539), .Y(n7679) );
  AOI222XL U2338 ( .A0(n596), .A1(n2592), .B0(n4914), .B1(n1255), .C0(n4880), 
        .C1(n540), .Y(n11475) );
  AOI222XL U2339 ( .A0(n597), .A1(n2775), .B0(n5222), .B1(n1249), .C0(n5188), 
        .C1(n541), .Y(n10599) );
  AOI222XL U2340 ( .A0(n598), .A1(n2957), .B0(n5468), .B1(n1243), .C0(n5434), 
        .C1(n542), .Y(n9723) );
  AOI222XL U2341 ( .A0(n599), .A1(n3139), .B0(n5696), .B1(n1237), .C0(n5662), 
        .C1(n543), .Y(n8847) );
  AOI222XL U2342 ( .A0(n600), .A1(n3318), .B0(n5932), .B1(n1231), .C0(n5898), 
        .C1(n544), .Y(n7971) );
  AOI22XL U2343 ( .A0(n17017), .A1(n2876), .B0(n2871), .B1(n17047), .Y(n17018)
         );
  AOI22XL U2344 ( .A0(n18277), .A1(n2634), .B0(n2629), .B1(n18307), .Y(n18278)
         );
  AOI22XL U2345 ( .A0(n15127), .A1(n3233), .B0(n3231), .B1(n15157), .Y(n15128)
         );
  AOI22XL U2346 ( .A0(n15442), .A1(n3172), .B0(n3170), .B1(n15472), .Y(n15443)
         );
  AOI22XL U2347 ( .A0(n18592), .A1(n2573), .B0(n2568), .B1(n18622), .Y(n18593)
         );
  AOI22XL U2348 ( .A0(n16702), .A1(n2936), .B0(n2932), .B1(n16732), .Y(n16703)
         );
  AOI22XL U2349 ( .A0(n14812), .A1(n3295), .B0(n3292), .B1(n14842), .Y(n14813)
         );
  AOI22XL U2350 ( .A0(n16387), .A1(n2997), .B0(n2993), .B1(n16417), .Y(n16388)
         );
  AOI22XL U2351 ( .A0(n17962), .A1(n2694), .B0(n2690), .B1(n17992), .Y(n17963)
         );
  AOI22XL U2352 ( .A0(n14497), .A1(n3355), .B0(n3353), .B1(n14527), .Y(n14498)
         );
  AOI22XL U2353 ( .A0(n16072), .A1(n3056), .B0(n3051), .B1(n16102), .Y(n16073)
         );
  AOI22XL U2354 ( .A0(n17647), .A1(n2752), .B0(n2750), .B1(n17677), .Y(n17648)
         );
  AOI22XL U2355 ( .A0(n14182), .A1(n3415), .B0(n3411), .B1(n14212), .Y(n14183)
         );
  AOI22XL U2356 ( .A0(n15757), .A1(n3117), .B0(n3112), .B1(n15787), .Y(n15758)
         );
  AOI22XL U2357 ( .A0(n17332), .A1(n2814), .B0(n2811), .B1(n17362), .Y(n17333)
         );
  AOI222XL U2358 ( .A0(n5375), .A1(n2898), .B0(n10067), .B1(n9900), .C0(n498), 
        .C1(n9988), .Y(n10066) );
  AOI222XL U2359 ( .A0(n6165), .A1(n3507), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n253), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .C0(n497), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n174), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n252) );
  AOI222XL U2360 ( .A0(n5021), .A1(n2658), .B0(n11235), .B1(n11068), .C0(n501), 
        .C1(n11156), .Y(n11234) );
  AOI222XL U2361 ( .A0(n5847), .A1(n3258), .B0(n8315), .B1(n8148), .C0(n500), 
        .C1(n8236), .Y(n8314) );
  AOI222XL U2362 ( .A0(n5105), .A1(n2717), .B0(n10943), .B1(n10776), .C0(n506), 
        .C1(n10864), .Y(n10942) );
  AOI222XL U2363 ( .A0(n6075), .A1(n3439), .B0(n7439), .B1(n7272), .C0(n510), 
        .C1(n7360), .Y(n7438) );
  AOI222XL U2364 ( .A0(n5611), .A1(n3080), .B0(n9191), .B1(n9024), .C0(n508), 
        .C1(n9112), .Y(n9190) );
  AOI222XL U2365 ( .A0(n5291), .A1(n2843), .B0(n10359), .B1(n10192), .C0(n512), 
        .C1(n10280), .Y(n10358) );
  AOI222XL U2366 ( .A0(n5535), .A1(n3022), .B0(n9483), .B1(n9316), .C0(n505), 
        .C1(n9404), .Y(n9482) );
  AOI222XL U2367 ( .A0(n5763), .A1(n3197), .B0(n8607), .B1(n8440), .C0(n499), 
        .C1(n8528), .Y(n8606) );
  AOI222XL U2368 ( .A0(n5999), .A1(n3382), .B0(n7731), .B1(n7564), .C0(n507), 
        .C1(n7652), .Y(n7730) );
  AOI222XL U2369 ( .A0(n4905), .A1(n2597), .B0(n11527), .B1(n11360), .C0(n502), 
        .C1(n11448), .Y(n11526) );
  AOI222XL U2370 ( .A0(n5213), .A1(n2782), .B0(n10651), .B1(n10484), .C0(n509), 
        .C1(n10572), .Y(n10650) );
  AOI222XL U2371 ( .A0(n5459), .A1(n2959), .B0(n9775), .B1(n9608), .C0(n503), 
        .C1(n9696), .Y(n9774) );
  AOI222XL U2372 ( .A0(n5687), .A1(n3141), .B0(n8899), .B1(n8732), .C0(n511), 
        .C1(n8820), .Y(n8898) );
  AOI222XL U2373 ( .A0(n5923), .A1(n3321), .B0(n8023), .B1(n7856), .C0(n504), 
        .C1(n7944), .Y(n8022) );
  AOI222XL U2374 ( .A0(n993), .A1(n498), .B0(n10040), .B1(n9970), .C0(n10041), 
        .C1(n698), .Y(n10039) );
  AOI222XL U2375 ( .A0(n1135), .A1(n497), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n226), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n227), .C1(n699), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n225) );
  AOI222XL U2376 ( .A0(n937), .A1(n501), .B0(n11208), .B1(n11138), .C0(n11209), 
        .C1(n700), .Y(n11207) );
  AOI222XL U2377 ( .A0(n1077), .A1(n500), .B0(n8288), .B1(n8218), .C0(n8289), 
        .C1(n701), .Y(n8287) );
  AOI222XL U2378 ( .A0(n951), .A1(n506), .B0(n10916), .B1(n10846), .C0(n10917), 
        .C1(n707), .Y(n10915) );
  AOI222XL U2379 ( .A0(n1035), .A1(n508), .B0(n9164), .B1(n9094), .C0(n9165), 
        .C1(n709), .Y(n9163) );
  AOI222XL U2380 ( .A0(n1119), .A1(n510), .B0(n7412), .B1(n7342), .C0(n7413), 
        .C1(n711), .Y(n7411) );
  AOI222XL U2381 ( .A0(n979), .A1(n512), .B0(n10332), .B1(n10262), .C0(n10333), 
        .C1(n713), .Y(n10331) );
  AOI222XL U2382 ( .A0(n1021), .A1(n505), .B0(n9456), .B1(n9386), .C0(n9457), 
        .C1(n706), .Y(n9455) );
  AOI222XL U2383 ( .A0(n1063), .A1(n499), .B0(n8580), .B1(n8510), .C0(n8581), 
        .C1(n702), .Y(n8579) );
  AOI222XL U2384 ( .A0(n1105), .A1(n507), .B0(n7704), .B1(n7634), .C0(n7705), 
        .C1(n708), .Y(n7703) );
  AOI222XL U2385 ( .A0(n923), .A1(n502), .B0(n11500), .B1(n11430), .C0(n11501), 
        .C1(n704), .Y(n11499) );
  AOI222XL U2386 ( .A0(n965), .A1(n509), .B0(n10624), .B1(n10554), .C0(n10625), 
        .C1(n710), .Y(n10623) );
  AOI222XL U2387 ( .A0(n1007), .A1(n503), .B0(n9748), .B1(n9678), .C0(n9749), 
        .C1(n703), .Y(n9747) );
  AOI222XL U2388 ( .A0(n1049), .A1(n511), .B0(n8872), .B1(n8802), .C0(n8873), 
        .C1(n712), .Y(n8871) );
  AOI222XL U2389 ( .A0(n1091), .A1(n504), .B0(n7996), .B1(n7926), .C0(n7997), 
        .C1(n705), .Y(n7995) );
  AOI211XL U2390 ( .A0(n5926), .A1(n14842), .B0(n14893), .C0(n15029), .Y(
        n15028) );
  AOI211XL U2391 ( .A0(n5614), .A1(n16102), .B0(n16153), .C0(n16289), .Y(
        n16288) );
  AOI211XL U2392 ( .A0(n5294), .A1(n17362), .B0(n17413), .C0(n17549), .Y(
        n17548) );
  AOI211XL U2393 ( .A0(n4908), .A1(n18622), .B0(n18673), .C0(n18809), .Y(
        n18808) );
  AOI211XL U2394 ( .A0(n5378), .A1(n17047), .B0(n17098), .C0(n17234), .Y(
        n17233) );
  AOI211XL U2395 ( .A0(n6149), .A1(n13897), .B0(n13948), .C0(n14084), .Y(
        n14083) );
  AOI211XL U2396 ( .A0(n5850), .A1(n15157), .B0(n15208), .C0(n15344), .Y(
        n15343) );
  AOI211XL U2397 ( .A0(n5024), .A1(n18307), .B0(n18358), .C0(n18494), .Y(
        n18493) );
  AOI211XL U2398 ( .A0(n5766), .A1(n15472), .B0(n15523), .C0(n15659), .Y(
        n15658) );
  AOI211XL U2399 ( .A0(n5462), .A1(n16732), .B0(n16783), .C0(n16919), .Y(
        n16918) );
  AOI211XL U2400 ( .A0(n5538), .A1(n16417), .B0(n16468), .C0(n16604), .Y(
        n16603) );
  AOI211XL U2401 ( .A0(n5108), .A1(n17992), .B0(n18043), .C0(n18179), .Y(
        n18178) );
  AOI211XL U2402 ( .A0(n6002), .A1(n14527), .B0(n14578), .C0(n14714), .Y(
        n14713) );
  AOI211XL U2403 ( .A0(n5216), .A1(n17677), .B0(n17728), .C0(n17864), .Y(
        n17863) );
  AOI211XL U2404 ( .A0(n6078), .A1(n14212), .B0(n14263), .C0(n14399), .Y(
        n14398) );
  AOI211XL U2405 ( .A0(n5690), .A1(n15787), .B0(n15838), .C0(n15974), .Y(
        n15973) );
  AOI211XL U2406 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n82), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n84), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n85), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n81) );
  AOI211XL U2407 ( .A0(n9899), .A1(n9900), .B0(n9901), .C0(n9902), .Y(n9898)
         );
  AOI211XL U2408 ( .A0(n11067), .A1(n11068), .B0(n11069), .C0(n11070), .Y(
        n11066) );
  AOI211XL U2409 ( .A0(n8147), .A1(n8148), .B0(n8149), .C0(n8150), .Y(n8146)
         );
  AOI211XL U2410 ( .A0(n10775), .A1(n10776), .B0(n10777), .C0(n10778), .Y(
        n10774) );
  AOI211XL U2411 ( .A0(n9023), .A1(n9024), .B0(n9025), .C0(n9026), .Y(n9022)
         );
  AOI211XL U2412 ( .A0(n7271), .A1(n7272), .B0(n7273), .C0(n7274), .Y(n7270)
         );
  AOI211XL U2413 ( .A0(n10191), .A1(n10192), .B0(n10193), .C0(n10194), .Y(
        n10190) );
  AOI211XL U2414 ( .A0(n9315), .A1(n9316), .B0(n9317), .C0(n9318), .Y(n9314)
         );
  AOI211XL U2415 ( .A0(n8439), .A1(n8440), .B0(n8441), .C0(n8442), .Y(n8438)
         );
  AOI211XL U2416 ( .A0(n7563), .A1(n7564), .B0(n7565), .C0(n7566), .Y(n7562)
         );
  AOI211XL U2417 ( .A0(n11359), .A1(n11360), .B0(n11361), .C0(n11362), .Y(
        n11358) );
  AOI211XL U2418 ( .A0(n10483), .A1(n10484), .B0(n10485), .C0(n10486), .Y(
        n10482) );
  AOI211XL U2419 ( .A0(n9607), .A1(n9608), .B0(n9609), .C0(n9610), .Y(n9606)
         );
  AOI211XL U2420 ( .A0(n8731), .A1(n8732), .B0(n8733), .C0(n8734), .Y(n8730)
         );
  AOI211XL U2421 ( .A0(n7855), .A1(n7856), .B0(n7857), .C0(n7858), .Y(n7854)
         );
  AOI22XL U2422 ( .A0(n698), .A1(n9900), .B0(n546), .B1(n9970), .Y(n10158) );
  AOI22XL U2423 ( .A0(n699), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .B0(
        n545), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n344) );
  AOI22XL U2424 ( .A0(n701), .A1(n8148), .B0(n548), .B1(n8218), .Y(n8406) );
  AOI22XL U2425 ( .A0(n700), .A1(n11068), .B0(n547), .B1(n11138), .Y(n11326)
         );
  AOI22XL U2426 ( .A0(n707), .A1(n10776), .B0(n549), .B1(n10846), .Y(n11034)
         );
  AOI22XL U2427 ( .A0(n711), .A1(n7272), .B0(n551), .B1(n7342), .Y(n7530) );
  AOI22XL U2428 ( .A0(n709), .A1(n9024), .B0(n550), .B1(n9094), .Y(n9282) );
  AOI22XL U2429 ( .A0(n713), .A1(n10192), .B0(n552), .B1(n10262), .Y(n10450)
         );
  AOI22XL U2430 ( .A0(n706), .A1(n9316), .B0(n553), .B1(n9386), .Y(n9574) );
  AOI22XL U2431 ( .A0(n702), .A1(n8440), .B0(n554), .B1(n8510), .Y(n8698) );
  AOI22XL U2432 ( .A0(n708), .A1(n7564), .B0(n555), .B1(n7634), .Y(n7822) );
  AOI22XL U2433 ( .A0(n704), .A1(n11360), .B0(n556), .B1(n11430), .Y(n11618)
         );
  AOI22XL U2434 ( .A0(n710), .A1(n10484), .B0(n557), .B1(n10554), .Y(n10742)
         );
  AOI22XL U2435 ( .A0(n703), .A1(n9608), .B0(n558), .B1(n9678), .Y(n9866) );
  AOI22XL U2436 ( .A0(n712), .A1(n8732), .B0(n559), .B1(n8802), .Y(n8990) );
  AOI22XL U2437 ( .A0(n705), .A1(n7856), .B0(n560), .B1(n7926), .Y(n8114) );
  AOI22XL U2438 ( .A0(n1001), .A1(n722), .B0(n993), .B1(n9970), .Y(n10153) );
  AOI22XL U2439 ( .A0(n1143), .A1(n723), .B0(n1135), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n339) );
  AOI22XL U2440 ( .A0(n1085), .A1(n725), .B0(n1077), .B1(n8218), .Y(n8401) );
  AOI22XL U2441 ( .A0(n945), .A1(n724), .B0(n937), .B1(n11138), .Y(n11321) );
  AOI22XL U2442 ( .A0(n959), .A1(n731), .B0(n951), .B1(n10846), .Y(n11029) );
  AOI22XL U2443 ( .A0(n1127), .A1(n735), .B0(n1119), .B1(n7342), .Y(n7525) );
  AOI22XL U2444 ( .A0(n1043), .A1(n733), .B0(n1035), .B1(n9094), .Y(n9277) );
  AOI22XL U2445 ( .A0(n987), .A1(n737), .B0(n979), .B1(n10262), .Y(n10445) );
  AOI22XL U2446 ( .A0(n1029), .A1(n730), .B0(n1021), .B1(n9386), .Y(n9569) );
  AOI22XL U2447 ( .A0(n1071), .A1(n726), .B0(n1063), .B1(n8510), .Y(n8693) );
  AOI22XL U2448 ( .A0(n1113), .A1(n732), .B0(n1105), .B1(n7634), .Y(n7817) );
  AOI22XL U2449 ( .A0(n931), .A1(n728), .B0(n923), .B1(n11430), .Y(n11613) );
  AOI22XL U2450 ( .A0(n973), .A1(n734), .B0(n965), .B1(n10554), .Y(n10737) );
  AOI22XL U2451 ( .A0(n1015), .A1(n727), .B0(n1007), .B1(n9678), .Y(n9861) );
  AOI22XL U2452 ( .A0(n1057), .A1(n736), .B0(n1049), .B1(n8802), .Y(n8985) );
  AOI22XL U2453 ( .A0(n1099), .A1(n729), .B0(n1091), .B1(n7926), .Y(n8109) );
  AOI222XL U2454 ( .A0(n5624), .A1(n9015), .B0(n1618), .B1(n9205), .C0(n5572), 
        .C1(n9037), .Y(n9204) );
  AOI222XL U2455 ( .A0(n4918), .A1(n11351), .B0(n1610), .B1(n11541), .C0(n4866), .C1(n11373), .Y(n11540) );
  AOI222XL U2456 ( .A0(n5936), .A1(n7847), .B0(n1622), .B1(n8037), .C0(n5884), 
        .C1(n7869), .Y(n8036) );
  AOI222XL U2457 ( .A0(n5776), .A1(n8431), .B0(n1620), .B1(n8621), .C0(n5724), 
        .C1(n8453), .Y(n8620) );
  AOI222XL U2458 ( .A0(n5472), .A1(n9599), .B0(n1616), .B1(n9789), .C0(n5420), 
        .C1(n9621), .Y(n9788) );
  AOI222XL U2459 ( .A0(n5304), .A1(n10183), .B0(n1614), .B1(n10373), .C0(n5252), .C1(n10205), .Y(n10372) );
  AOI222XL U2460 ( .A0(n5118), .A1(n10767), .B0(n1612), .B1(n10957), .C0(n5066), .C1(n10789), .Y(n10956) );
  AOI222XL U2461 ( .A0(n5388), .A1(n9891), .B0(n1615), .B1(n10081), .C0(n5336), 
        .C1(n9913), .Y(n10080) );
  AOI222XL U2462 ( .A0(n6175), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), 
        .B0(n1625), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n267), .C0(n6132), 
        .C1(top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n266) );
  AOI222XL U2463 ( .A0(n5034), .A1(n11059), .B0(n1611), .B1(n11249), .C0(n4982), .C1(n11081), .Y(n11248) );
  AOI222XL U2464 ( .A0(n5860), .A1(n8139), .B0(n1621), .B1(n8329), .C0(n5808), 
        .C1(n8161), .Y(n8328) );
  AOI222XL U2465 ( .A0(n6088), .A1(n7263), .B0(n1624), .B1(n7453), .C0(n6036), 
        .C1(n7285), .Y(n7452) );
  AOI222XL U2466 ( .A0(n5548), .A1(n9307), .B0(n1617), .B1(n9497), .C0(n5496), 
        .C1(n9329), .Y(n9496) );
  AOI222XL U2467 ( .A0(n6012), .A1(n7555), .B0(n1623), .B1(n7745), .C0(n5960), 
        .C1(n7577), .Y(n7744) );
  AOI222XL U2468 ( .A0(n5226), .A1(n10475), .B0(n1613), .B1(n10665), .C0(n5174), .C1(n10497), .Y(n10664) );
  AOI222XL U2469 ( .A0(n5700), .A1(n8723), .B0(n1619), .B1(n8913), .C0(n5648), 
        .C1(n8745), .Y(n8912) );
  AOI222XL U2470 ( .A0(n999), .A1(n2883), .B0(n997), .B1(n1003), .C0(n5362), 
        .C1(n17007), .Y(n17064) );
  AOI222XL U2471 ( .A0(n1138), .A1(n3487), .B0(n1136), .B1(n1142), .C0(n6130), 
        .C1(n13857), .Y(n13914) );
  AOI222XL U2472 ( .A0(n943), .A1(n2644), .B0(n941), .B1(n947), .C0(n5008), 
        .C1(n18267), .Y(n18324) );
  AOI222XL U2473 ( .A0(n1083), .A1(n3246), .B0(n1081), .B1(n1087), .C0(n5834), 
        .C1(n15117), .Y(n15174) );
  AOI222XL U2474 ( .A0(n1069), .A1(n3186), .B0(n1067), .B1(n1073), .C0(n5750), 
        .C1(n15432), .Y(n15489) );
  AOI222XL U2475 ( .A0(n929), .A1(n2584), .B0(n927), .B1(n933), .C0(n4892), 
        .C1(n18582), .Y(n18639) );
  AOI222XL U2476 ( .A0(n1013), .A1(n2944), .B0(n1011), .B1(n1017), .C0(n5446), 
        .C1(n16692), .Y(n16749) );
  AOI222XL U2477 ( .A0(n1097), .A1(n3307), .B0(n1095), .B1(n1101), .C0(n5910), 
        .C1(n14802), .Y(n14859) );
  AOI222XL U2478 ( .A0(n1027), .A1(n3008), .B0(n1025), .B1(n1031), .C0(n5522), 
        .C1(n16377), .Y(n16434) );
  AOI222XL U2479 ( .A0(n957), .A1(n2706), .B0(n955), .B1(n961), .C0(n5092), 
        .C1(n17952), .Y(n18009) );
  AOI222XL U2480 ( .A0(n1111), .A1(n3369), .B0(n1109), .B1(n1115), .C0(n5986), 
        .C1(n14487), .Y(n14544) );
  AOI222XL U2481 ( .A0(n1041), .A1(n3066), .B0(n1039), .B1(n1045), .C0(n5598), 
        .C1(n16062), .Y(n16119) );
  AOI222XL U2482 ( .A0(n971), .A1(n2766), .B0(n969), .B1(n975), .C0(n5200), 
        .C1(n17637), .Y(n17694) );
  AOI222XL U2483 ( .A0(n1125), .A1(n3426), .B0(n1123), .B1(n1129), .C0(n6062), 
        .C1(n14172), .Y(n14229) );
  AOI222XL U2484 ( .A0(n1055), .A1(n3128), .B0(n1053), .B1(n1059), .C0(n5674), 
        .C1(n15747), .Y(n15804) );
  AOI222XL U2485 ( .A0(n985), .A1(n2826), .B0(n983), .B1(n989), .C0(n5278), 
        .C1(n17322), .Y(n17379) );
  AOI222XL U2486 ( .A0(n999), .A1(n17047), .B0(n370), .B1(n633), .C0(n417), 
        .C1(n5363), .Y(n17123) );
  AOI222XL U2487 ( .A0(n1138), .A1(n13897), .B0(n369), .B1(n634), .C0(n418), 
        .C1(n6131), .Y(n13973) );
  AOI222XL U2488 ( .A0(n943), .A1(n18307), .B0(n371), .B1(n635), .C0(n419), 
        .C1(n5009), .Y(n18383) );
  AOI222XL U2489 ( .A0(n1083), .A1(n15157), .B0(n372), .B1(n636), .C0(n420), 
        .C1(n5835), .Y(n15233) );
  AOI222XL U2490 ( .A0(n1069), .A1(n15472), .B0(n373), .B1(n637), .C0(n426), 
        .C1(n5751), .Y(n15548) );
  AOI222XL U2491 ( .A0(n929), .A1(n18622), .B0(n374), .B1(n638), .C0(n428), 
        .C1(n4893), .Y(n18698) );
  AOI222XL U2492 ( .A0(n1013), .A1(n16732), .B0(n375), .B1(n639), .C0(n430), 
        .C1(n5447), .Y(n16808) );
  AOI222XL U2493 ( .A0(n1097), .A1(n14842), .B0(n376), .B1(n640), .C0(n432), 
        .C1(n5911), .Y(n14918) );
  AOI222XL U2494 ( .A0(n1027), .A1(n16417), .B0(n377), .B1(n641), .C0(n425), 
        .C1(n5523), .Y(n16493) );
  AOI222XL U2495 ( .A0(n957), .A1(n17992), .B0(n378), .B1(n642), .C0(n421), 
        .C1(n5093), .Y(n18068) );
  AOI222XL U2496 ( .A0(n1111), .A1(n14527), .B0(n379), .B1(n643), .C0(n427), 
        .C1(n5987), .Y(n14603) );
  AOI222XL U2497 ( .A0(n1041), .A1(n16102), .B0(n380), .B1(n644), .C0(n422), 
        .C1(n5599), .Y(n16178) );
  AOI222XL U2498 ( .A0(n971), .A1(n17677), .B0(n381), .B1(n645), .C0(n429), 
        .C1(n5201), .Y(n17753) );
  AOI222XL U2499 ( .A0(n1125), .A1(n14212), .B0(n382), .B1(n646), .C0(n423), 
        .C1(n6063), .Y(n14288) );
  AOI222XL U2500 ( .A0(n1055), .A1(n15787), .B0(n383), .B1(n647), .C0(n431), 
        .C1(n5675), .Y(n15863) );
  AOI222XL U2501 ( .A0(n985), .A1(n17362), .B0(n384), .B1(n648), .C0(n424), 
        .C1(n5279), .Y(n17438) );
  AOI211XL U2502 ( .A0(n1065), .A1(n1294), .B0(n15462), .C0(n15445), .Y(n15459) );
  AOI211XL U2503 ( .A0(n953), .A1(n1318), .B0(n17982), .C0(n17965), .Y(n17979)
         );
  AOI211XL U2504 ( .A0(n1121), .A1(n1282), .B0(n14202), .C0(n14185), .Y(n14199) );
  AOI211XL U2505 ( .A0(n925), .A1(n1324), .B0(n18612), .C0(n18595), .Y(n18609)
         );
  AOI211XL U2506 ( .A0(n1093), .A1(n1288), .B0(n14832), .C0(n14815), .Y(n14829) );
  AOI211XL U2507 ( .A0(n1037), .A1(n1300), .B0(n16092), .C0(n16075), .Y(n16089) );
  AOI211XL U2508 ( .A0(n981), .A1(n1312), .B0(n17352), .C0(n17335), .Y(n17349)
         );
  AOI211XL U2509 ( .A0(n1134), .A1(n1279), .B0(n13887), .C0(n13870), .Y(n13884) );
  AOI211XL U2510 ( .A0(n995), .A1(n1309), .B0(n17037), .C0(n17020), .Y(n17034)
         );
  AOI211XL U2511 ( .A0(n939), .A1(n1321), .B0(n18297), .C0(n18280), .Y(n18294)
         );
  AOI211XL U2512 ( .A0(n1079), .A1(n1291), .B0(n15147), .C0(n15130), .Y(n15144) );
  AOI211XL U2513 ( .A0(n1009), .A1(n1306), .B0(n16722), .C0(n16705), .Y(n16719) );
  AOI211XL U2514 ( .A0(n1023), .A1(n1303), .B0(n16407), .C0(n16390), .Y(n16404) );
  AOI211XL U2515 ( .A0(n1107), .A1(n1285), .B0(n14517), .C0(n14500), .Y(n14514) );
  AOI211XL U2516 ( .A0(n967), .A1(n1315), .B0(n17667), .C0(n17650), .Y(n17664)
         );
  AOI211XL U2517 ( .A0(n1051), .A1(n1297), .B0(n15777), .C0(n15760), .Y(n15774) );
  AND4X1 U2518 ( .A(n9961), .B(n10072), .C(n9999), .D(n10045), .Y(n10071) );
  AND4X1 U2519 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n146), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n258), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n185), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n231), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n257) );
  AND4X1 U2520 ( .A(n11129), .B(n11240), .C(n11167), .D(n11213), .Y(n11239) );
  AND4X1 U2521 ( .A(n8209), .B(n8320), .C(n8247), .D(n8293), .Y(n8319) );
  AND4X1 U2522 ( .A(n10837), .B(n10948), .C(n10875), .D(n10921), .Y(n10947) );
  AND4X1 U2523 ( .A(n7333), .B(n7444), .C(n7371), .D(n7417), .Y(n7443) );
  AND4X1 U2524 ( .A(n9085), .B(n9196), .C(n9123), .D(n9169), .Y(n9195) );
  AND4X1 U2525 ( .A(n10253), .B(n10364), .C(n10291), .D(n10337), .Y(n10363) );
  AND4X1 U2526 ( .A(n9377), .B(n9488), .C(n9415), .D(n9461), .Y(n9487) );
  AND4X1 U2527 ( .A(n8501), .B(n8612), .C(n8539), .D(n8585), .Y(n8611) );
  AND4X1 U2528 ( .A(n7625), .B(n7736), .C(n7663), .D(n7709), .Y(n7735) );
  AND4X1 U2529 ( .A(n11421), .B(n11532), .C(n11459), .D(n11505), .Y(n11531) );
  AND4X1 U2530 ( .A(n10545), .B(n10656), .C(n10583), .D(n10629), .Y(n10655) );
  AND4X1 U2531 ( .A(n9669), .B(n9780), .C(n9707), .D(n9753), .Y(n9779) );
  AND4X1 U2532 ( .A(n8793), .B(n8904), .C(n8831), .D(n8877), .Y(n8903) );
  AND4X1 U2533 ( .A(n7917), .B(n8028), .C(n7955), .D(n8001), .Y(n8027) );
  AOI31XL U2534 ( .A0(n932), .A1(n2566), .A2(n18780), .B0(n253), .Y(n18784) );
  AOI31XL U2535 ( .A0(n1044), .A1(n3049), .A2(n16260), .B0(n248), .Y(n16264)
         );
  AOI31XL U2536 ( .A0(n988), .A1(n2809), .A2(n17520), .B0(n244), .Y(n17524) );
  AOI31XL U2537 ( .A0(n960), .A1(n2687), .A2(n18150), .B0(n250), .Y(n18154) );
  AOI31XL U2538 ( .A0(n1128), .A1(n3409), .A2(n14370), .B0(n246), .Y(n14374)
         );
  AOI31XL U2539 ( .A0(n1100), .A1(n3290), .A2(n15000), .B0(n252), .Y(n15004)
         );
  AOI31XL U2540 ( .A0(n1072), .A1(n3168), .A2(n15630), .B0(n255), .Y(n15634)
         );
  AOI31XL U2541 ( .A0(n1002), .A1(n2869), .A2(n17205), .B0(n259), .Y(n17209)
         );
  AOI31XL U2542 ( .A0(n1141), .A1(n3470), .A2(n14055), .B0(n258), .Y(n14059)
         );
  AOI31XL U2543 ( .A0(n946), .A1(n2627), .A2(n18465), .B0(n257), .Y(n18469) );
  AOI31XL U2544 ( .A0(n1086), .A1(n3229), .A2(n15315), .B0(n256), .Y(n15319)
         );
  AOI31XL U2545 ( .A0(n1016), .A1(n2930), .A2(n16890), .B0(n254), .Y(n16894)
         );
  AOI31XL U2546 ( .A0(n1030), .A1(n2991), .A2(n16575), .B0(n251), .Y(n16579)
         );
  AOI31XL U2547 ( .A0(n1114), .A1(n3351), .A2(n14685), .B0(n249), .Y(n14689)
         );
  AOI31XL U2548 ( .A0(n974), .A1(n2749), .A2(n17835), .B0(n247), .Y(n17839) );
  AOI31XL U2549 ( .A0(n1058), .A1(n3110), .A2(n15945), .B0(n245), .Y(n15949)
         );
  AOI221XL U2550 ( .A0(n1615), .A1(n698), .B0(n10112), .B1(n9891), .C0(n5376), 
        .Y(n10111) );
  AOI221XL U2551 ( .A0(n1625), .A1(n699), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n298), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n74), .C0(n6166), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n297) );
  AOI221XL U2552 ( .A0(n1621), .A1(n701), .B0(n8360), .B1(n8139), .C0(n5848), 
        .Y(n8359) );
  AOI221XL U2553 ( .A0(n1611), .A1(n700), .B0(n11280), .B1(n11059), .C0(n5022), 
        .Y(n11279) );
  AOI221XL U2554 ( .A0(n1612), .A1(n707), .B0(n10988), .B1(n10767), .C0(n5106), 
        .Y(n10987) );
  AOI221XL U2555 ( .A0(n1624), .A1(n711), .B0(n7484), .B1(n7263), .C0(n6076), 
        .Y(n7483) );
  AOI221XL U2556 ( .A0(n1618), .A1(n709), .B0(n9236), .B1(n9015), .C0(n5612), 
        .Y(n9235) );
  AOI221XL U2557 ( .A0(n1614), .A1(n713), .B0(n10404), .B1(n10183), .C0(n5292), 
        .Y(n10403) );
  AOI221XL U2558 ( .A0(n1617), .A1(n706), .B0(n9528), .B1(n9307), .C0(n5536), 
        .Y(n9527) );
  AOI221XL U2559 ( .A0(n1620), .A1(n702), .B0(n8652), .B1(n8431), .C0(n5764), 
        .Y(n8651) );
  AOI221XL U2560 ( .A0(n1623), .A1(n708), .B0(n7776), .B1(n7555), .C0(n6000), 
        .Y(n7775) );
  AOI221XL U2561 ( .A0(n1610), .A1(n704), .B0(n11572), .B1(n11351), .C0(n4906), 
        .Y(n11571) );
  AOI221XL U2562 ( .A0(n1613), .A1(n710), .B0(n10696), .B1(n10475), .C0(n5214), 
        .Y(n10695) );
  AOI221XL U2563 ( .A0(n1616), .A1(n703), .B0(n9820), .B1(n9599), .C0(n5460), 
        .Y(n9819) );
  AOI221XL U2564 ( .A0(n1619), .A1(n712), .B0(n8944), .B1(n8723), .C0(n5688), 
        .Y(n8943) );
  AOI221XL U2565 ( .A0(n1622), .A1(n705), .B0(n8068), .B1(n7847), .C0(n5924), 
        .Y(n8067) );
  AOI21XL U2566 ( .A0(n5363), .A1(n1310), .B0(n5352), .Y(n17169) );
  AOI21XL U2567 ( .A0(n6131), .A1(n1280), .B0(n6120), .Y(n14019) );
  AOI21XL U2568 ( .A0(n5009), .A1(n1322), .B0(n4998), .Y(n18429) );
  AOI21XL U2569 ( .A0(n5835), .A1(n1292), .B0(n5824), .Y(n15279) );
  AOI21XL U2570 ( .A0(n5751), .A1(n1295), .B0(n5740), .Y(n15594) );
  AOI21XL U2571 ( .A0(n4893), .A1(n1325), .B0(n4882), .Y(n18744) );
  AOI21XL U2572 ( .A0(n5447), .A1(n1307), .B0(n5436), .Y(n16854) );
  AOI21XL U2573 ( .A0(n5911), .A1(n1289), .B0(n5900), .Y(n14964) );
  AOI21XL U2574 ( .A0(n5523), .A1(n1304), .B0(n5512), .Y(n16539) );
  AOI21XL U2575 ( .A0(n5093), .A1(n1319), .B0(n5082), .Y(n18114) );
  AOI21XL U2576 ( .A0(n5987), .A1(n1286), .B0(n5976), .Y(n14649) );
  AOI21XL U2577 ( .A0(n5599), .A1(n1301), .B0(n5588), .Y(n16224) );
  AOI21XL U2578 ( .A0(n5201), .A1(n1316), .B0(n5190), .Y(n17799) );
  AOI21XL U2579 ( .A0(n6063), .A1(n1283), .B0(n6052), .Y(n14334) );
  AOI21XL U2580 ( .A0(n5675), .A1(n1298), .B0(n5664), .Y(n15909) );
  AOI21XL U2581 ( .A0(n5279), .A1(n1313), .B0(n5268), .Y(n17484) );
  AOI211XL U2582 ( .A0(n9030), .A1(n9024), .B0(n9291), .C0(n9292), .Y(n9290)
         );
  AOI22XL U2583 ( .A0(n5612), .A1(n9015), .B0(n5624), .B1(n3063), .Y(n9289) );
  AOI211XL U2584 ( .A0(n10198), .A1(n10192), .B0(n10459), .C0(n10460), .Y(
        n10458) );
  AOI22XL U2585 ( .A0(n5292), .A1(n10183), .B0(n5304), .B1(n2823), .Y(n10457)
         );
  AOI211XL U2586 ( .A0(n11366), .A1(n11360), .B0(n11627), .C0(n11628), .Y(
        n11626) );
  AOI22XL U2587 ( .A0(n4906), .A1(n11351), .B0(n4918), .B1(n2580), .Y(n11625)
         );
  AOI211XL U2588 ( .A0(n7862), .A1(n7856), .B0(n8123), .C0(n8124), .Y(n8122)
         );
  AOI22XL U2589 ( .A0(n5924), .A1(n7847), .B0(n5936), .B1(n3307), .Y(n8121) );
  AOI211XL U2590 ( .A0(n10782), .A1(n10776), .B0(n11043), .C0(n11044), .Y(
        n11042) );
  AOI22XL U2591 ( .A0(n5106), .A1(n10767), .B0(n5118), .B1(n2702), .Y(n11041)
         );
  AOI211XL U2592 ( .A0(n8446), .A1(n8440), .B0(n8707), .C0(n8708), .Y(n8706)
         );
  AOI22XL U2593 ( .A0(n5764), .A1(n8431), .B0(n5776), .B1(n3182), .Y(n8705) );
  AOI211XL U2594 ( .A0(n9614), .A1(n9608), .B0(n9875), .C0(n9876), .Y(n9874)
         );
  AOI22XL U2595 ( .A0(n5460), .A1(n9599), .B0(n5472), .B1(n2944), .Y(n9873) );
  AOI211XL U2596 ( .A0(n9906), .A1(n9900), .B0(n10167), .C0(n10168), .Y(n10166) );
  AOI22XL U2597 ( .A0(n5376), .A1(n9891), .B0(n5388), .B1(n2883), .Y(n10165)
         );
  AOI211XL U2598 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n89), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n353), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n354), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n352) );
  AOI22XL U2599 ( .A0(n6166), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), 
        .B0(n6175), .B1(n3486), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n351) );
  AOI211XL U2600 ( .A0(n8154), .A1(n8148), .B0(n8415), .C0(n8416), .Y(n8414)
         );
  AOI22XL U2601 ( .A0(n5848), .A1(n8139), .B0(n5860), .B1(n3246), .Y(n8413) );
  AOI211XL U2602 ( .A0(n11074), .A1(n11068), .B0(n11335), .C0(n11336), .Y(
        n11334) );
  AOI22XL U2603 ( .A0(n5022), .A1(n11059), .B0(n5034), .B1(n2641), .Y(n11333)
         );
  AOI211XL U2604 ( .A0(n7278), .A1(n7272), .B0(n7539), .C0(n7540), .Y(n7538)
         );
  AOI22XL U2605 ( .A0(n6076), .A1(n7263), .B0(n6088), .B1(n3423), .Y(n7537) );
  AOI211XL U2606 ( .A0(n9322), .A1(n9316), .B0(n9583), .C0(n9584), .Y(n9582)
         );
  AOI22XL U2607 ( .A0(n5536), .A1(n9307), .B0(n5548), .B1(n3008), .Y(n9581) );
  AOI211XL U2608 ( .A0(n7570), .A1(n7564), .B0(n7831), .C0(n7832), .Y(n7830)
         );
  AOI22XL U2609 ( .A0(n6000), .A1(n7555), .B0(n6012), .B1(n3365), .Y(n7829) );
  AOI211XL U2610 ( .A0(n10490), .A1(n10484), .B0(n10751), .C0(n10752), .Y(
        n10750) );
  AOI22XL U2611 ( .A0(n5214), .A1(n10475), .B0(n5226), .B1(n2762), .Y(n10749)
         );
  AOI211XL U2612 ( .A0(n8738), .A1(n8732), .B0(n8999), .C0(n9000), .Y(n8998)
         );
  AOI22XL U2613 ( .A0(n5688), .A1(n8723), .B0(n5700), .B1(n3124), .Y(n8997) );
  AOI211XL U2614 ( .A0(n723), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), 
        .B0(n6137), .C0(n6155), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n73) );
  AOI211XL U2615 ( .A0(n722), .A1(n9891), .B0(n5341), .C0(n5365), .Y(n9890) );
  AOI211XL U2616 ( .A0(n724), .A1(n11059), .B0(n4987), .C0(n5011), .Y(n11058)
         );
  AOI211XL U2617 ( .A0(n725), .A1(n8139), .B0(n5813), .C0(n5837), .Y(n8138) );
  AOI211XL U2618 ( .A0(n731), .A1(n10767), .B0(n5071), .C0(n5095), .Y(n10766)
         );
  AOI211XL U2619 ( .A0(n733), .A1(n9015), .B0(n5577), .C0(n5601), .Y(n9014) );
  AOI211XL U2620 ( .A0(n735), .A1(n7263), .B0(n6041), .C0(n6065), .Y(n7262) );
  AOI211XL U2621 ( .A0(n737), .A1(n10183), .B0(n5257), .C0(n5281), .Y(n10182)
         );
  AOI211XL U2622 ( .A0(n730), .A1(n9307), .B0(n5501), .C0(n5525), .Y(n9306) );
  AOI211XL U2623 ( .A0(n726), .A1(n8431), .B0(n5729), .C0(n5753), .Y(n8430) );
  AOI211XL U2624 ( .A0(n732), .A1(n7555), .B0(n5965), .C0(n5989), .Y(n7554) );
  AOI211XL U2625 ( .A0(n728), .A1(n11351), .B0(n4871), .C0(n4895), .Y(n11350)
         );
  AOI211XL U2626 ( .A0(n734), .A1(n10475), .B0(n5179), .C0(n5203), .Y(n10474)
         );
  AOI211XL U2627 ( .A0(n727), .A1(n9599), .B0(n5425), .C0(n5449), .Y(n9598) );
  AOI211XL U2628 ( .A0(n736), .A1(n8723), .B0(n5653), .C0(n5677), .Y(n8722) );
  AOI211XL U2629 ( .A0(n729), .A1(n7847), .B0(n5889), .C0(n5913), .Y(n7846) );
  AOI211XL U2630 ( .A0(n997), .A1(n1310), .B0(n17037), .C0(n5360), .Y(n17148)
         );
  AOI211XL U2631 ( .A0(n1136), .A1(n1280), .B0(n13887), .C0(n6128), .Y(n13998)
         );
  AOI211XL U2632 ( .A0(n941), .A1(n1322), .B0(n18297), .C0(n5006), .Y(n18408)
         );
  AOI211XL U2633 ( .A0(n1081), .A1(n1292), .B0(n15147), .C0(n5832), .Y(n15258)
         );
  AOI211XL U2634 ( .A0(n1067), .A1(n1295), .B0(n15462), .C0(n5748), .Y(n15573)
         );
  AOI211XL U2635 ( .A0(n927), .A1(n1325), .B0(n18612), .C0(n4890), .Y(n18723)
         );
  AOI211XL U2636 ( .A0(n1011), .A1(n1307), .B0(n16722), .C0(n5444), .Y(n16833)
         );
  AOI211XL U2637 ( .A0(n1095), .A1(n1289), .B0(n14832), .C0(n5908), .Y(n14943)
         );
  AOI211XL U2638 ( .A0(n1025), .A1(n1304), .B0(n16407), .C0(n5520), .Y(n16518)
         );
  AOI211XL U2639 ( .A0(n955), .A1(n1319), .B0(n17982), .C0(n5090), .Y(n18093)
         );
  AOI211XL U2640 ( .A0(n1109), .A1(n1286), .B0(n14517), .C0(n5984), .Y(n14628)
         );
  AOI211XL U2641 ( .A0(n1039), .A1(n1301), .B0(n16092), .C0(n5596), .Y(n16203)
         );
  AOI211XL U2642 ( .A0(n969), .A1(n1316), .B0(n17667), .C0(n5198), .Y(n17778)
         );
  AOI211XL U2643 ( .A0(n1123), .A1(n1283), .B0(n14202), .C0(n6060), .Y(n14313)
         );
  AOI211XL U2644 ( .A0(n1053), .A1(n1298), .B0(n15777), .C0(n5672), .Y(n15888)
         );
  AOI211XL U2645 ( .A0(n983), .A1(n1313), .B0(n17352), .C0(n5276), .Y(n17463)
         );
  AOI32XL U2646 ( .A0(n3448), .A1(n1279), .A2(n6117), .B0(n6107), .B1(n14098), 
        .Y(n14097) );
  AOI32XL U2647 ( .A0(n2847), .A1(n1309), .A2(n5334), .B0(n5325), .B1(n17248), 
        .Y(n17247) );
  AOI32XL U2648 ( .A0(n2605), .A1(n1321), .A2(n4980), .B0(n4971), .B1(n18508), 
        .Y(n18507) );
  AOI32XL U2649 ( .A0(n3207), .A1(n1291), .A2(n5806), .B0(n5797), .B1(n15358), 
        .Y(n15357) );
  AOI32XL U2650 ( .A0(n3146), .A1(n1294), .A2(n5722), .B0(n5713), .B1(n15673), 
        .Y(n15672) );
  AOI32XL U2651 ( .A0(n2544), .A1(n1324), .A2(n4864), .B0(n4855), .B1(n18823), 
        .Y(n18822) );
  AOI32XL U2652 ( .A0(n2908), .A1(n1306), .A2(n5418), .B0(n5409), .B1(n16933), 
        .Y(n16932) );
  AOI32XL U2653 ( .A0(n3268), .A1(n1288), .A2(n5882), .B0(n5873), .B1(n15043), 
        .Y(n15042) );
  AOI32XL U2654 ( .A0(n2969), .A1(n1303), .A2(n5494), .B0(n5485), .B1(n16618), 
        .Y(n16617) );
  AOI32XL U2655 ( .A0(n2666), .A1(n1318), .A2(n5064), .B0(n5055), .B1(n18193), 
        .Y(n18192) );
  AOI32XL U2656 ( .A0(n3329), .A1(n1285), .A2(n5958), .B0(n5949), .B1(n14728), 
        .Y(n14727) );
  AOI32XL U2657 ( .A0(n3027), .A1(n1300), .A2(n5570), .B0(n5561), .B1(n16303), 
        .Y(n16302) );
  AOI32XL U2658 ( .A0(n2726), .A1(n1315), .A2(n5172), .B0(n5163), .B1(n17878), 
        .Y(n17877) );
  AOI32XL U2659 ( .A0(n3387), .A1(n1282), .A2(n6034), .B0(n6025), .B1(n14413), 
        .Y(n14412) );
  AOI32XL U2660 ( .A0(n3088), .A1(n1297), .A2(n5646), .B0(n5637), .B1(n15988), 
        .Y(n15987) );
  AOI32XL U2661 ( .A0(n2787), .A1(n1312), .A2(n5250), .B0(n5241), .B1(n17563), 
        .Y(n17562) );
  AOI222XL U2662 ( .A0(n5380), .A1(n2886), .B0(n17060), .B1(n17061), .C0(n5378), .C1(n2880), .Y(n17054) );
  AOI222XL U2663 ( .A0(n5026), .A1(n2644), .B0(n18320), .B1(n18321), .C0(n5024), .C1(n2638), .Y(n18314) );
  AOI222XL U2664 ( .A0(n5852), .A1(n3246), .B0(n15170), .B1(n15171), .C0(n5850), .C1(n3240), .Y(n15164) );
  AOI222XL U2665 ( .A0(n5768), .A1(n3186), .B0(n15485), .B1(n15486), .C0(n5766), .C1(n3179), .Y(n15479) );
  AOI222XL U2666 ( .A0(n4910), .A1(n2584), .B0(n18635), .B1(n18636), .C0(n4908), .C1(n2577), .Y(n18629) );
  AOI222XL U2667 ( .A0(n5464), .A1(n2949), .B0(n16745), .B1(n16746), .C0(n5462), .C1(n2941), .Y(n16739) );
  AOI222XL U2668 ( .A0(n5928), .A1(n3307), .B0(n14855), .B1(n14856), .C0(n5926), .C1(n3301), .Y(n14849) );
  AOI222XL U2669 ( .A0(n5540), .A1(n3008), .B0(n16430), .B1(n16431), .C0(n5538), .C1(n3002), .Y(n16424) );
  AOI222XL U2670 ( .A0(n5110), .A1(n2706), .B0(n18005), .B1(n18006), .C0(n5108), .C1(n2699), .Y(n17999) );
  AOI222XL U2671 ( .A0(n6004), .A1(n3369), .B0(n14540), .B1(n14541), .C0(n6002), .C1(n3362), .Y(n14534) );
  AOI222XL U2672 ( .A0(n5616), .A1(n3066), .B0(n16115), .B1(n16116), .C0(n5614), .C1(n3060), .Y(n16109) );
  AOI222XL U2673 ( .A0(n5218), .A1(n2766), .B0(n17690), .B1(n17691), .C0(n5216), .C1(n2759), .Y(n17684) );
  AOI222XL U2674 ( .A0(n6080), .A1(n3426), .B0(n14225), .B1(n14226), .C0(n6078), .C1(n3420), .Y(n14219) );
  AOI222XL U2675 ( .A0(n5692), .A1(n3128), .B0(n15800), .B1(n15801), .C0(n5690), .C1(n3121), .Y(n15794) );
  AOI222XL U2676 ( .A0(n5296), .A1(n2826), .B0(n17375), .B1(n17376), .C0(n5294), .C1(n2820), .Y(n17369) );
  AOI222XL U2677 ( .A0(n6151), .A1(n3487), .B0(n13910), .B1(n13911), .C0(n6149), .C1(n3490), .Y(n13904) );
  AOI222XL U2678 ( .A0(n5388), .A1(n2895), .B0(n135), .B1(n2888), .C0(n5384), 
        .C1(n433), .Y(n9967) );
  AOI222XL U2679 ( .A0(n6175), .A1(n3501), .B0(n136), .B1(n3489), .C0(n6169), 
        .C1(n434), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n152) );
  AOI222XL U2680 ( .A0(n5034), .A1(n2652), .B0(n137), .B1(n2646), .C0(n5030), 
        .C1(n435), .Y(n11135) );
  AOI222XL U2681 ( .A0(n5860), .A1(n3255), .B0(n138), .B1(n3248), .C0(n5856), 
        .C1(n436), .Y(n8215) );
  AOI222XL U2682 ( .A0(n5118), .A1(n2719), .B0(n139), .B1(n2708), .C0(n5114), 
        .C1(n442), .Y(n10843) );
  AOI222XL U2683 ( .A0(n5624), .A1(n3074), .B0(n140), .B1(n3068), .C0(n5620), 
        .C1(n444), .Y(n9091) );
  AOI222XL U2684 ( .A0(n6088), .A1(n3441), .B0(n141), .B1(n3428), .C0(n6084), 
        .C1(n446), .Y(n7339) );
  AOI222XL U2685 ( .A0(n5304), .A1(n2842), .B0(n142), .B1(n2828), .C0(n5300), 
        .C1(n448), .Y(n10259) );
  AOI222XL U2686 ( .A0(n5548), .A1(n3021), .B0(n143), .B1(n3010), .C0(n5544), 
        .C1(n441), .Y(n9383) );
  AOI222XL U2687 ( .A0(n5776), .A1(n3194), .B0(n144), .B1(n3188), .C0(n5772), 
        .C1(n437), .Y(n8507) );
  AOI222XL U2688 ( .A0(n6012), .A1(n3381), .B0(n145), .B1(n3371), .C0(n6008), 
        .C1(n443), .Y(n7631) );
  AOI222XL U2689 ( .A0(n4918), .A1(n2591), .B0(n146), .B1(n2586), .C0(n4914), 
        .C1(n439), .Y(n11427) );
  AOI222XL U2690 ( .A0(n5226), .A1(n2776), .B0(n147), .B1(n2768), .C0(n5222), 
        .C1(n445), .Y(n10551) );
  AOI222XL U2691 ( .A0(n5472), .A1(n2956), .B0(n148), .B1(n2949), .C0(n5468), 
        .C1(n438), .Y(n9675) );
  AOI222XL U2692 ( .A0(n5700), .A1(n3140), .B0(n149), .B1(n3130), .C0(n5696), 
        .C1(n447), .Y(n8799) );
  AOI222XL U2693 ( .A0(n5936), .A1(n3323), .B0(n150), .B1(n3309), .C0(n5932), 
        .C1(n440), .Y(n7923) );
  OAI211XL U2694 ( .A0(n2881), .A1(n9960), .B0(n9955), .C0(n9896), .Y(n10020)
         );
  OAI211XL U2695 ( .A0(n3482), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n145), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n140), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n206) );
  OAI211XL U2696 ( .A0(n2639), .A1(n11128), .B0(n11123), .C0(n11064), .Y(
        n11188) );
  OAI211XL U2697 ( .A0(n3241), .A1(n8208), .B0(n8203), .C0(n8144), .Y(n8268)
         );
  OAI211XL U2698 ( .A0(n2700), .A1(n10836), .B0(n10831), .C0(n10772), .Y(
        n10896) );
  OAI211XL U2699 ( .A0(n3061), .A1(n9084), .B0(n9079), .C0(n9020), .Y(n9144)
         );
  OAI211XL U2700 ( .A0(n3421), .A1(n7332), .B0(n7327), .C0(n7268), .Y(n7392)
         );
  OAI211XL U2701 ( .A0(n2821), .A1(n10252), .B0(n10247), .C0(n10188), .Y(
        n10312) );
  OAI211XL U2702 ( .A0(n3003), .A1(n9376), .B0(n9371), .C0(n9312), .Y(n9436)
         );
  OAI211XL U2703 ( .A0(n3180), .A1(n8500), .B0(n8495), .C0(n8436), .Y(n8560)
         );
  OAI211XL U2704 ( .A0(n3363), .A1(n7624), .B0(n7619), .C0(n7560), .Y(n7684)
         );
  OAI211XL U2705 ( .A0(n2578), .A1(n11420), .B0(n11415), .C0(n11356), .Y(
        n11480) );
  OAI211XL U2706 ( .A0(n2760), .A1(n10544), .B0(n10539), .C0(n10480), .Y(
        n10604) );
  OAI211XL U2707 ( .A0(n2942), .A1(n9668), .B0(n9663), .C0(n9604), .Y(n9728)
         );
  OAI211XL U2708 ( .A0(n3122), .A1(n8792), .B0(n8787), .C0(n8728), .Y(n8852)
         );
  OAI211XL U2709 ( .A0(n3302), .A1(n7916), .B0(n7911), .C0(n7852), .Y(n7976)
         );
  AOI31XL U2710 ( .A0(n2867), .A1(n17047), .A2(n5335), .B0(n17137), .Y(n17131)
         );
  AOI31XL U2711 ( .A0(n3468), .A1(n13897), .A2(n6118), .B0(n13987), .Y(n13981)
         );
  AOI31XL U2712 ( .A0(n2625), .A1(n18307), .A2(n4981), .B0(n18397), .Y(n18391)
         );
  AOI31XL U2713 ( .A0(n3227), .A1(n15157), .A2(n5807), .B0(n15247), .Y(n15241)
         );
  AOI31XL U2714 ( .A0(n3166), .A1(n15472), .A2(n5723), .B0(n15562), .Y(n15556)
         );
  AOI31XL U2715 ( .A0(n2564), .A1(n18622), .A2(n4865), .B0(n18712), .Y(n18706)
         );
  AOI31XL U2716 ( .A0(n2928), .A1(n16732), .A2(n5419), .B0(n16822), .Y(n16816)
         );
  AOI31XL U2717 ( .A0(n3288), .A1(n14842), .A2(n5883), .B0(n14932), .Y(n14926)
         );
  AOI31XL U2718 ( .A0(n2989), .A1(n16417), .A2(n5495), .B0(n16507), .Y(n16501)
         );
  AOI31XL U2719 ( .A0(n2686), .A1(n17992), .A2(n5065), .B0(n18082), .Y(n18076)
         );
  AOI31XL U2720 ( .A0(n3349), .A1(n14527), .A2(n5959), .B0(n14617), .Y(n14611)
         );
  AOI31XL U2721 ( .A0(n3047), .A1(n16102), .A2(n5571), .B0(n16192), .Y(n16186)
         );
  AOI31XL U2722 ( .A0(n2746), .A1(n17677), .A2(n5173), .B0(n17767), .Y(n17761)
         );
  AOI31XL U2723 ( .A0(n3407), .A1(n14212), .A2(n6035), .B0(n14302), .Y(n14296)
         );
  AOI31XL U2724 ( .A0(n3108), .A1(n15787), .A2(n5647), .B0(n15877), .Y(n15871)
         );
  AOI31XL U2725 ( .A0(n2807), .A1(n17362), .A2(n5251), .B0(n17452), .Y(n17446)
         );
  AOI211XL U2726 ( .A0(n10723), .A1(n2732), .B0(n10724), .C0(n10584), .Y(
        n10703) );
  AOI211XL U2727 ( .A0(n9555), .A1(n2975), .B0(n9556), .C0(n9416), .Y(n9535)
         );
  AOI211XL U2728 ( .A0(n7803), .A1(n3335), .B0(n7804), .C0(n7664), .Y(n7783)
         );
  AOI211XL U2729 ( .A0(n8971), .A1(n3094), .B0(n8972), .C0(n8832), .Y(n8951)
         );
  AOI211XL U2730 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n325), .A1(n3454), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n326), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n186), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n305) );
  AOI211XL U2731 ( .A0(n10139), .A1(n2853), .B0(n10140), .C0(n10000), .Y(
        n10119) );
  AOI211XL U2732 ( .A0(n11307), .A1(n2611), .B0(n11308), .C0(n11168), .Y(
        n11287) );
  AOI211XL U2733 ( .A0(n8387), .A1(n3213), .B0(n8388), .C0(n8248), .Y(n8367)
         );
  AOI211XL U2734 ( .A0(n11015), .A1(n2672), .B0(n11016), .C0(n10876), .Y(
        n10995) );
  AOI211XL U2735 ( .A0(n9263), .A1(n3033), .B0(n9264), .C0(n9124), .Y(n9243)
         );
  AOI211XL U2736 ( .A0(n7511), .A1(n3393), .B0(n7512), .C0(n7372), .Y(n7491)
         );
  AOI211XL U2737 ( .A0(n10431), .A1(n2793), .B0(n10432), .C0(n10292), .Y(
        n10411) );
  AOI211XL U2738 ( .A0(n8679), .A1(n3152), .B0(n8680), .C0(n8540), .Y(n8659)
         );
  AOI211XL U2739 ( .A0(n11599), .A1(n2550), .B0(n11600), .C0(n11460), .Y(
        n11579) );
  AOI211XL U2740 ( .A0(n9847), .A1(n2914), .B0(n9848), .C0(n9708), .Y(n9827)
         );
  AOI211XL U2741 ( .A0(n8095), .A1(n3274), .B0(n8096), .C0(n7956), .Y(n8075)
         );
  AOI31XL U2742 ( .A0(n13246), .A1(n13247), .A2(n13248), .B0(n1667), .Y(n13245) );
  NAND4XL U2743 ( .A(n10065), .B(n15), .C(n9947), .D(n10066), .Y(n10059) );
  NAND4XL U2744 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n251), .B(n14), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n132), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n252), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n245) );
  NAND4XL U2745 ( .A(n11233), .B(n16), .C(n11115), .D(n11234), .Y(n11227) );
  NAND4XL U2746 ( .A(n8313), .B(n17), .C(n8195), .D(n8314), .Y(n8307) );
  NAND4XL U2747 ( .A(n10941), .B(n18), .C(n10823), .D(n10942), .Y(n10935) );
  NAND4XL U2748 ( .A(n7437), .B(n20), .C(n7319), .D(n7438), .Y(n7431) );
  NAND4XL U2749 ( .A(n9189), .B(n19), .C(n9071), .D(n9190), .Y(n9183) );
  NAND4XL U2750 ( .A(n10357), .B(n21), .C(n10239), .D(n10358), .Y(n10351) );
  NAND4XL U2751 ( .A(n9481), .B(n22), .C(n9363), .D(n9482), .Y(n9475) );
  NAND4XL U2752 ( .A(n8605), .B(n23), .C(n8487), .D(n8606), .Y(n8599) );
  NAND4XL U2753 ( .A(n7729), .B(n24), .C(n7611), .D(n7730), .Y(n7723) );
  NAND4XL U2754 ( .A(n11525), .B(n25), .C(n11407), .D(n11526), .Y(n11519) );
  NAND4XL U2755 ( .A(n10649), .B(n26), .C(n10531), .D(n10650), .Y(n10643) );
  NAND4XL U2756 ( .A(n9773), .B(n27), .C(n9655), .D(n9774), .Y(n9767) );
  NAND4XL U2757 ( .A(n8897), .B(n28), .C(n8779), .D(n8898), .Y(n8891) );
  NAND4XL U2758 ( .A(n8021), .B(n29), .C(n7903), .D(n8022), .Y(n8015) );
  AOI211XL U2759 ( .A0(n16998), .A1(n17047), .B0(n17037), .C0(n5359), .Y(
        n17194) );
  AOI211XL U2760 ( .A0(n13848), .A1(n13897), .B0(n13887), .C0(n6127), .Y(
        n14044) );
  AOI211XL U2761 ( .A0(n18258), .A1(n18307), .B0(n18297), .C0(n5005), .Y(
        n18454) );
  AOI211XL U2762 ( .A0(n15108), .A1(n15157), .B0(n15147), .C0(n5831), .Y(
        n15304) );
  AOI211XL U2763 ( .A0(n15423), .A1(n15472), .B0(n15462), .C0(n5747), .Y(
        n15619) );
  AOI211XL U2764 ( .A0(n16683), .A1(n16732), .B0(n16722), .C0(n5443), .Y(
        n16879) );
  AOI211XL U2765 ( .A0(n18573), .A1(n18622), .B0(n18612), .C0(n4889), .Y(
        n18769) );
  AOI211XL U2766 ( .A0(n14793), .A1(n14842), .B0(n14832), .C0(n5907), .Y(
        n14989) );
  AOI211XL U2767 ( .A0(n16368), .A1(n16417), .B0(n16407), .C0(n5519), .Y(
        n16564) );
  AOI211XL U2768 ( .A0(n17943), .A1(n17992), .B0(n17982), .C0(n5089), .Y(
        n18139) );
  AOI211XL U2769 ( .A0(n14478), .A1(n14527), .B0(n14517), .C0(n5983), .Y(
        n14674) );
  AOI211XL U2770 ( .A0(n16053), .A1(n16102), .B0(n16092), .C0(n5595), .Y(
        n16249) );
  AOI211XL U2771 ( .A0(n17628), .A1(n17677), .B0(n17667), .C0(n5197), .Y(
        n17824) );
  AOI211XL U2772 ( .A0(n14163), .A1(n14212), .B0(n14202), .C0(n6059), .Y(
        n14359) );
  AOI211XL U2773 ( .A0(n15738), .A1(n15787), .B0(n15777), .C0(n5671), .Y(
        n15934) );
  AOI211XL U2774 ( .A0(n17313), .A1(n17362), .B0(n17352), .C0(n5275), .Y(
        n17509) );
  OAI211XL U2775 ( .A0(n57), .A1(n1309), .B0(n17129), .C0(n17136), .Y(n17133)
         );
  AOI22XL U2776 ( .A0(n998), .A1(n17017), .B0(n995), .B1(n2880), .Y(n17136) );
  OAI211XL U2777 ( .A0(n58), .A1(n1279), .B0(n13979), .C0(n13986), .Y(n13983)
         );
  AOI22XL U2778 ( .A0(n1137), .A1(n13867), .B0(n1134), .B1(n3481), .Y(n13986)
         );
  OAI211XL U2779 ( .A0(n59), .A1(n1321), .B0(n18389), .C0(n18396), .Y(n18393)
         );
  AOI22XL U2780 ( .A0(n942), .A1(n18277), .B0(n939), .B1(n2638), .Y(n18396) );
  OAI211XL U2781 ( .A0(n60), .A1(n1291), .B0(n15239), .C0(n15246), .Y(n15243)
         );
  AOI22XL U2782 ( .A0(n1082), .A1(n15127), .B0(n1079), .B1(n3240), .Y(n15246)
         );
  OAI211XL U2783 ( .A0(n61), .A1(n1294), .B0(n15554), .C0(n15561), .Y(n15558)
         );
  AOI22XL U2784 ( .A0(n1068), .A1(n15442), .B0(n1065), .B1(n3179), .Y(n15561)
         );
  OAI211XL U2785 ( .A0(n63), .A1(n1324), .B0(n18704), .C0(n18711), .Y(n18708)
         );
  AOI22XL U2786 ( .A0(n928), .A1(n18592), .B0(n925), .B1(n2577), .Y(n18711) );
  OAI211XL U2787 ( .A0(n62), .A1(n1306), .B0(n16814), .C0(n16821), .Y(n16818)
         );
  AOI22XL U2788 ( .A0(n1012), .A1(n16702), .B0(n1009), .B1(n2941), .Y(n16821)
         );
  OAI211XL U2789 ( .A0(n64), .A1(n1288), .B0(n14924), .C0(n14931), .Y(n14928)
         );
  AOI22XL U2790 ( .A0(n1096), .A1(n14812), .B0(n1093), .B1(n3301), .Y(n14931)
         );
  OAI211XL U2791 ( .A0(n65), .A1(n1303), .B0(n16499), .C0(n16506), .Y(n16503)
         );
  AOI22XL U2792 ( .A0(n1026), .A1(n16387), .B0(n1023), .B1(n3002), .Y(n16506)
         );
  OAI211XL U2793 ( .A0(n66), .A1(n1318), .B0(n18074), .C0(n18081), .Y(n18078)
         );
  AOI22XL U2794 ( .A0(n956), .A1(n17962), .B0(n953), .B1(n2699), .Y(n18081) );
  OAI211XL U2795 ( .A0(n67), .A1(n1285), .B0(n14609), .C0(n14616), .Y(n14613)
         );
  AOI22XL U2796 ( .A0(n1110), .A1(n14497), .B0(n1107), .B1(n3362), .Y(n14616)
         );
  OAI211XL U2797 ( .A0(n68), .A1(n1300), .B0(n16184), .C0(n16191), .Y(n16188)
         );
  AOI22XL U2798 ( .A0(n1040), .A1(n16072), .B0(n1037), .B1(n3060), .Y(n16191)
         );
  OAI211XL U2799 ( .A0(n69), .A1(n1315), .B0(n17759), .C0(n17766), .Y(n17763)
         );
  AOI22XL U2800 ( .A0(n970), .A1(n17647), .B0(n967), .B1(n2759), .Y(n17766) );
  OAI211XL U2801 ( .A0(n70), .A1(n1282), .B0(n14294), .C0(n14301), .Y(n14298)
         );
  AOI22XL U2802 ( .A0(n1124), .A1(n14182), .B0(n1121), .B1(n3420), .Y(n14301)
         );
  OAI211XL U2803 ( .A0(n71), .A1(n1297), .B0(n15869), .C0(n15876), .Y(n15873)
         );
  AOI22XL U2804 ( .A0(n1054), .A1(n15757), .B0(n1051), .B1(n3121), .Y(n15876)
         );
  OAI211XL U2805 ( .A0(n72), .A1(n1312), .B0(n17444), .C0(n17451), .Y(n17448)
         );
  AOI22XL U2806 ( .A0(n984), .A1(n17332), .B0(n981), .B1(n2820), .Y(n17451) );
  AOI31XL U2807 ( .A0(n9930), .A1(n90), .A2(n10157), .B0(n2853), .Y(n10156) );
  AOI31XL U2808 ( .A0(n10011), .A1(n15), .A2(n10158), .B0(n2861), .Y(n10155)
         );
  AOI22XL U2809 ( .A0(n698), .A1(n433), .B0(n5348), .B1(n9913), .Y(n10157) );
  AOI31XL U2810 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n115), .A1(n91), .A2(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n343), .B0(n3454), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n342) );
  AOI31XL U2811 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n197), .A1(n14), .A2(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n344), .B0(n3463), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n341) );
  AOI22XL U2812 ( .A0(n699), .A1(n434), .B0(n6144), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n343) );
  AOI31XL U2813 ( .A0(n8178), .A1(n93), .A2(n8405), .B0(n3213), .Y(n8404) );
  AOI31XL U2814 ( .A0(n8259), .A1(n17), .A2(n8406), .B0(n3221), .Y(n8403) );
  AOI22XL U2815 ( .A0(n701), .A1(n436), .B0(n5820), .B1(n8161), .Y(n8405) );
  AOI31XL U2816 ( .A0(n11098), .A1(n92), .A2(n11325), .B0(n2611), .Y(n11324)
         );
  AOI31XL U2817 ( .A0(n11179), .A1(n16), .A2(n11326), .B0(n2614), .Y(n11323)
         );
  AOI22XL U2818 ( .A0(n700), .A1(n435), .B0(n4994), .B1(n11081), .Y(n11325) );
  AOI31XL U2819 ( .A0(n10806), .A1(n94), .A2(n11033), .B0(n2672), .Y(n11032)
         );
  AOI31XL U2820 ( .A0(n10887), .A1(n18), .A2(n11034), .B0(n2680), .Y(n11031)
         );
  AOI22XL U2821 ( .A0(n707), .A1(n442), .B0(n5078), .B1(n10789), .Y(n11033) );
  AOI31XL U2822 ( .A0(n7302), .A1(n95), .A2(n7529), .B0(n3393), .Y(n7528) );
  AOI31XL U2823 ( .A0(n7383), .A1(n20), .A2(n7530), .B0(n3396), .Y(n7527) );
  AOI22XL U2824 ( .A0(n711), .A1(n446), .B0(n6048), .B1(n7285), .Y(n7529) );
  AOI31XL U2825 ( .A0(n9054), .A1(n96), .A2(n9281), .B0(n3033), .Y(n9280) );
  AOI31XL U2826 ( .A0(n9135), .A1(n19), .A2(n9282), .B0(n3036), .Y(n9279) );
  AOI22XL U2827 ( .A0(n709), .A1(n444), .B0(n5584), .B1(n9037), .Y(n9281) );
  AOI31XL U2828 ( .A0(n10222), .A1(n97), .A2(n10449), .B0(n2793), .Y(n10448)
         );
  AOI31XL U2829 ( .A0(n10303), .A1(n21), .A2(n10450), .B0(n2796), .Y(n10447)
         );
  AOI22XL U2830 ( .A0(n713), .A1(n448), .B0(n5264), .B1(n10205), .Y(n10449) );
  AOI31XL U2831 ( .A0(n9346), .A1(n98), .A2(n9573), .B0(n2975), .Y(n9572) );
  AOI31XL U2832 ( .A0(n9427), .A1(n22), .A2(n9574), .B0(n2978), .Y(n9571) );
  AOI22XL U2833 ( .A0(n706), .A1(n441), .B0(n5508), .B1(n9329), .Y(n9573) );
  AOI31XL U2834 ( .A0(n8470), .A1(n99), .A2(n8697), .B0(n3152), .Y(n8696) );
  AOI31XL U2835 ( .A0(n8551), .A1(n23), .A2(n8698), .B0(n3155), .Y(n8695) );
  AOI22XL U2836 ( .A0(n702), .A1(n437), .B0(n5736), .B1(n8453), .Y(n8697) );
  AOI31XL U2837 ( .A0(n7594), .A1(n100), .A2(n7821), .B0(n3335), .Y(n7820) );
  AOI31XL U2838 ( .A0(n7675), .A1(n24), .A2(n7822), .B0(n3338), .Y(n7819) );
  AOI22XL U2839 ( .A0(n708), .A1(n443), .B0(n5972), .B1(n7577), .Y(n7821) );
  AOI31XL U2840 ( .A0(n11390), .A1(n101), .A2(n11617), .B0(n2550), .Y(n11616)
         );
  AOI31XL U2841 ( .A0(n11471), .A1(n25), .A2(n11618), .B0(n2558), .Y(n11615)
         );
  AOI22XL U2842 ( .A0(n704), .A1(n439), .B0(n4878), .B1(n11373), .Y(n11617) );
  AOI31XL U2843 ( .A0(n10514), .A1(n102), .A2(n10741), .B0(n2732), .Y(n10740)
         );
  AOI31XL U2844 ( .A0(n10595), .A1(n26), .A2(n10742), .B0(n2740), .Y(n10739)
         );
  AOI22XL U2845 ( .A0(n710), .A1(n445), .B0(n5186), .B1(n10497), .Y(n10741) );
  AOI31XL U2846 ( .A0(n9638), .A1(n103), .A2(n9865), .B0(n2914), .Y(n9864) );
  AOI31XL U2847 ( .A0(n9719), .A1(n27), .A2(n9866), .B0(n2917), .Y(n9863) );
  AOI22XL U2848 ( .A0(n703), .A1(n438), .B0(n5432), .B1(n9621), .Y(n9865) );
  AOI31XL U2849 ( .A0(n8762), .A1(n104), .A2(n8989), .B0(n3094), .Y(n8988) );
  AOI31XL U2850 ( .A0(n8843), .A1(n28), .A2(n8990), .B0(n3102), .Y(n8987) );
  AOI22XL U2851 ( .A0(n712), .A1(n447), .B0(n5660), .B1(n8745), .Y(n8989) );
  AOI31XL U2852 ( .A0(n7886), .A1(n105), .A2(n8113), .B0(n3274), .Y(n8112) );
  AOI31XL U2853 ( .A0(n7967), .A1(n29), .A2(n8114), .B0(n3277), .Y(n8111) );
  AOI22XL U2854 ( .A0(n705), .A1(n440), .B0(n5896), .B1(n7869), .Y(n8113) );
  AOI211XL U2855 ( .A0(n135), .A1(n433), .B0(n10020), .C0(n5349), .Y(n10017)
         );
  AOI211XL U2856 ( .A0(n137), .A1(n435), .B0(n11188), .C0(n4995), .Y(n11185)
         );
  AOI211XL U2857 ( .A0(n138), .A1(n436), .B0(n8268), .C0(n5821), .Y(n8265) );
  AOI211XL U2858 ( .A0(n139), .A1(n442), .B0(n10896), .C0(n5079), .Y(n10893)
         );
  AOI211XL U2859 ( .A0(n140), .A1(n444), .B0(n9144), .C0(n5585), .Y(n9141) );
  AOI211XL U2860 ( .A0(n141), .A1(n446), .B0(n7392), .C0(n6049), .Y(n7389) );
  AOI211XL U2861 ( .A0(n142), .A1(n448), .B0(n10312), .C0(n5265), .Y(n10309)
         );
  AOI211XL U2862 ( .A0(n143), .A1(n441), .B0(n9436), .C0(n5509), .Y(n9433) );
  AOI211XL U2863 ( .A0(n144), .A1(n437), .B0(n8560), .C0(n5737), .Y(n8557) );
  AOI211XL U2864 ( .A0(n145), .A1(n443), .B0(n7684), .C0(n5973), .Y(n7681) );
  AOI211XL U2865 ( .A0(n146), .A1(n439), .B0(n11480), .C0(n4879), .Y(n11477)
         );
  AOI211XL U2866 ( .A0(n147), .A1(n445), .B0(n10604), .C0(n5187), .Y(n10601)
         );
  AOI211XL U2867 ( .A0(n148), .A1(n438), .B0(n9728), .C0(n5433), .Y(n9725) );
  AOI211XL U2868 ( .A0(n149), .A1(n447), .B0(n8852), .C0(n5661), .Y(n8849) );
  AOI211XL U2869 ( .A0(n150), .A1(n440), .B0(n7976), .C0(n5897), .Y(n7973) );
  AOI211XL U2870 ( .A0(n136), .A1(n434), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n206), .C0(n6145), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n203) );
  NAND4XL U2871 ( .A(n9885), .B(n9956), .C(n10010), .D(n10039), .Y(n10025) );
  NAND4XL U2872 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n67), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n141), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n196), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n225), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n211) );
  NAND4XL U2873 ( .A(n11053), .B(n11124), .C(n11178), .D(n11207), .Y(n11193)
         );
  NAND4XL U2874 ( .A(n8133), .B(n8204), .C(n8258), .D(n8287), .Y(n8273) );
  NAND4XL U2875 ( .A(n10761), .B(n10832), .C(n10886), .D(n10915), .Y(n10901)
         );
  NAND4XL U2876 ( .A(n9009), .B(n9080), .C(n9134), .D(n9163), .Y(n9149) );
  NAND4XL U2877 ( .A(n7257), .B(n7328), .C(n7382), .D(n7411), .Y(n7397) );
  NAND4XL U2878 ( .A(n10177), .B(n10248), .C(n10302), .D(n10331), .Y(n10317)
         );
  NAND4XL U2879 ( .A(n9301), .B(n9372), .C(n9426), .D(n9455), .Y(n9441) );
  NAND4XL U2880 ( .A(n8425), .B(n8496), .C(n8550), .D(n8579), .Y(n8565) );
  NAND4XL U2881 ( .A(n7549), .B(n7620), .C(n7674), .D(n7703), .Y(n7689) );
  NAND4XL U2882 ( .A(n11345), .B(n11416), .C(n11470), .D(n11499), .Y(n11485)
         );
  NAND4XL U2883 ( .A(n10469), .B(n10540), .C(n10594), .D(n10623), .Y(n10609)
         );
  NAND4XL U2884 ( .A(n9593), .B(n9664), .C(n9718), .D(n9747), .Y(n9733) );
  NAND4XL U2885 ( .A(n8717), .B(n8788), .C(n8842), .D(n8871), .Y(n8857) );
  NAND4XL U2886 ( .A(n7841), .B(n7912), .C(n7966), .D(n7995), .Y(n7981) );
  AOI21XL U2887 ( .A0(n169), .A1(n18604), .B0(n2554), .Y(n18760) );
  AOI21XL U2888 ( .A0(n175), .A1(n16084), .B0(n3037), .Y(n16240) );
  AOI21XL U2889 ( .A0(n179), .A1(n17344), .B0(n2797), .Y(n17500) );
  AOI21XL U2890 ( .A0(n173), .A1(n17974), .B0(n2676), .Y(n18130) );
  AOI21XL U2891 ( .A0(n177), .A1(n14194), .B0(n3397), .Y(n14350) );
  AOI21XL U2892 ( .A0(n171), .A1(n14824), .B0(n3278), .Y(n14980) );
  AOI21XL U2893 ( .A0(n168), .A1(n15454), .B0(n3156), .Y(n15610) );
  AOI21XL U2894 ( .A0(n164), .A1(n17029), .B0(n2857), .Y(n17185) );
  AOI21XL U2895 ( .A0(n165), .A1(n13879), .B0(n3458), .Y(n14035) );
  AOI21XL U2896 ( .A0(n166), .A1(n18289), .B0(n2615), .Y(n18445) );
  AOI21XL U2897 ( .A0(n167), .A1(n15139), .B0(n3217), .Y(n15295) );
  AOI21XL U2898 ( .A0(n170), .A1(n16714), .B0(n2918), .Y(n16870) );
  AOI21XL U2899 ( .A0(n172), .A1(n16399), .B0(n2979), .Y(n16555) );
  AOI21XL U2900 ( .A0(n174), .A1(n14509), .B0(n3339), .Y(n14665) );
  AOI21XL U2901 ( .A0(n176), .A1(n17659), .B0(n2736), .Y(n17815) );
  AOI21XL U2902 ( .A0(n178), .A1(n15769), .B0(n3098), .Y(n15925) );
  AOI22XL U2903 ( .A0(n15433), .A1(n1295), .B0(n469), .B1(n5718), .Y(n15465)
         );
  AOI22XL U2904 ( .A0(n17953), .A1(n1319), .B0(n474), .B1(n5060), .Y(n17985)
         );
  AOI22XL U2905 ( .A0(n14173), .A1(n1283), .B0(n478), .B1(n6030), .Y(n14205)
         );
  AOI22XL U2906 ( .A0(n18583), .A1(n1325), .B0(n471), .B1(n4860), .Y(n18615)
         );
  AOI22XL U2907 ( .A0(n14803), .A1(n1289), .B0(n472), .B1(n5878), .Y(n14835)
         );
  AOI22XL U2908 ( .A0(n16063), .A1(n1301), .B0(n476), .B1(n5566), .Y(n16095)
         );
  AOI22XL U2909 ( .A0(n17323), .A1(n1313), .B0(n480), .B1(n5246), .Y(n17355)
         );
  AOI22XL U2910 ( .A0(n17008), .A1(n1310), .B0(n465), .B1(n5330), .Y(n17040)
         );
  AOI22XL U2911 ( .A0(n18268), .A1(n1322), .B0(n467), .B1(n4976), .Y(n18300)
         );
  AOI22XL U2912 ( .A0(n15118), .A1(n1292), .B0(n468), .B1(n5802), .Y(n15150)
         );
  AOI22XL U2913 ( .A0(n16693), .A1(n1307), .B0(n470), .B1(n5414), .Y(n16725)
         );
  AOI22XL U2914 ( .A0(n16378), .A1(n1304), .B0(n473), .B1(n5490), .Y(n16410)
         );
  AOI22XL U2915 ( .A0(n14488), .A1(n1286), .B0(n475), .B1(n5954), .Y(n14520)
         );
  AOI22XL U2916 ( .A0(n17638), .A1(n1316), .B0(n477), .B1(n5168), .Y(n17670)
         );
  AOI22XL U2917 ( .A0(n15748), .A1(n1298), .B0(n479), .B1(n5642), .Y(n15780)
         );
  AOI22XL U2918 ( .A0(n13858), .A1(n1280), .B0(n466), .B1(n6114), .Y(n13890)
         );
  AOI222XL U2919 ( .A0(n5388), .A1(n9970), .B0(n562), .B1(n2888), .C0(n546), 
        .C1(n1245), .Y(n9969) );
  AOI222XL U2920 ( .A0(n6175), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), 
        .B0(n561), .B1(n3484), .C0(n545), .C1(n1327), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n155) );
  AOI222XL U2921 ( .A0(n5034), .A1(n11138), .B0(n563), .B1(n2646), .C0(n547), 
        .C1(n1253), .Y(n11137) );
  AOI222XL U2922 ( .A0(n5860), .A1(n8218), .B0(n564), .B1(n3248), .C0(n548), 
        .C1(n1233), .Y(n8217) );
  AOI222XL U2923 ( .A0(n5118), .A1(n10846), .B0(n565), .B1(n2708), .C0(n549), 
        .C1(n1251), .Y(n10845) );
  AOI222XL U2924 ( .A0(n5624), .A1(n9094), .B0(n566), .B1(n3068), .C0(n550), 
        .C1(n1239), .Y(n9093) );
  AOI222XL U2925 ( .A0(n6088), .A1(n7342), .B0(n567), .B1(n3428), .C0(n551), 
        .C1(n1227), .Y(n7341) );
  AOI222XL U2926 ( .A0(n5304), .A1(n10262), .B0(n568), .B1(n2828), .C0(n552), 
        .C1(n1247), .Y(n10261) );
  AOI222XL U2927 ( .A0(n5548), .A1(n9386), .B0(n569), .B1(n3010), .C0(n553), 
        .C1(n1241), .Y(n9385) );
  AOI222XL U2928 ( .A0(n5776), .A1(n8510), .B0(n570), .B1(n3188), .C0(n554), 
        .C1(n1235), .Y(n8509) );
  AOI222XL U2929 ( .A0(n6012), .A1(n7634), .B0(n571), .B1(n3371), .C0(n555), 
        .C1(n1229), .Y(n7633) );
  AOI222XL U2930 ( .A0(n4918), .A1(n11430), .B0(n572), .B1(n2586), .C0(n556), 
        .C1(n1255), .Y(n11429) );
  AOI222XL U2931 ( .A0(n5226), .A1(n10554), .B0(n573), .B1(n2768), .C0(n557), 
        .C1(n1249), .Y(n10553) );
  AOI222XL U2932 ( .A0(n5472), .A1(n9678), .B0(n574), .B1(n2949), .C0(n558), 
        .C1(n1243), .Y(n9677) );
  AOI222XL U2933 ( .A0(n5700), .A1(n8802), .B0(n575), .B1(n3130), .C0(n559), 
        .C1(n1237), .Y(n8801) );
  AOI222XL U2934 ( .A0(n5936), .A1(n7926), .B0(n576), .B1(n3309), .C0(n560), 
        .C1(n1231), .Y(n7925) );
  AOI21XL U2935 ( .A0(n995), .A1(n17047), .B0(n17121), .Y(n17120) );
  AOI21XL U2936 ( .A0(n1134), .A1(n13897), .B0(n13971), .Y(n13970) );
  AOI21XL U2937 ( .A0(n939), .A1(n18307), .B0(n18381), .Y(n18380) );
  AOI21XL U2938 ( .A0(n1079), .A1(n15157), .B0(n15231), .Y(n15230) );
  AOI21XL U2939 ( .A0(n1065), .A1(n15472), .B0(n15546), .Y(n15545) );
  AOI21XL U2940 ( .A0(n925), .A1(n18622), .B0(n18696), .Y(n18695) );
  AOI21XL U2941 ( .A0(n1009), .A1(n16732), .B0(n16806), .Y(n16805) );
  AOI21XL U2942 ( .A0(n1093), .A1(n14842), .B0(n14916), .Y(n14915) );
  AOI21XL U2943 ( .A0(n1023), .A1(n16417), .B0(n16491), .Y(n16490) );
  AOI21XL U2944 ( .A0(n953), .A1(n17992), .B0(n18066), .Y(n18065) );
  AOI21XL U2945 ( .A0(n1107), .A1(n14527), .B0(n14601), .Y(n14600) );
  AOI21XL U2946 ( .A0(n1037), .A1(n16102), .B0(n16176), .Y(n16175) );
  AOI21XL U2947 ( .A0(n967), .A1(n17677), .B0(n17751), .Y(n17750) );
  AOI21XL U2948 ( .A0(n1121), .A1(n14212), .B0(n14286), .Y(n14285) );
  AOI21XL U2949 ( .A0(n1051), .A1(n15787), .B0(n15861), .Y(n15860) );
  AOI21XL U2950 ( .A0(n981), .A1(n17362), .B0(n17436), .Y(n17435) );
  AOI222XL U2951 ( .A0(n2558), .A1(n18853), .B0(n4857), .B1(n1325), .C0(n4858), 
        .C1(n18622), .Y(n18852) );
  AOI222XL U2952 ( .A0(n3283), .A1(n15073), .B0(n5875), .B1(n1289), .C0(n5876), 
        .C1(n14842), .Y(n15072) );
  AOI222XL U2953 ( .A0(n3042), .A1(n16333), .B0(n5563), .B1(n1301), .C0(n5564), 
        .C1(n16102), .Y(n16332) );
  AOI222XL U2954 ( .A0(n2802), .A1(n17593), .B0(n5243), .B1(n1313), .C0(n5244), 
        .C1(n17362), .Y(n17592) );
  AOI222XL U2955 ( .A0(n3161), .A1(n15703), .B0(n5715), .B1(n1295), .C0(n5716), 
        .C1(n15472), .Y(n15702) );
  AOI222XL U2956 ( .A0(n2681), .A1(n18223), .B0(n5057), .B1(n1319), .C0(n5058), 
        .C1(n17992), .Y(n18222) );
  AOI222XL U2957 ( .A0(n3402), .A1(n14443), .B0(n6027), .B1(n1283), .C0(n6028), 
        .C1(n14212), .Y(n14442) );
  AOI222XL U2958 ( .A0(n2862), .A1(n17278), .B0(n5327), .B1(n1310), .C0(n5328), 
        .C1(n17047), .Y(n17277) );
  AOI222XL U2959 ( .A0(n3463), .A1(n14128), .B0(n6111), .B1(n1280), .C0(n6112), 
        .C1(n13897), .Y(n14127) );
  AOI222XL U2960 ( .A0(n3222), .A1(n15388), .B0(n5799), .B1(n1292), .C0(n5800), 
        .C1(n15157), .Y(n15387) );
  AOI222XL U2961 ( .A0(n2620), .A1(n18538), .B0(n4973), .B1(n1322), .C0(n4974), 
        .C1(n18307), .Y(n18537) );
  AOI222XL U2962 ( .A0(n2923), .A1(n16963), .B0(n5411), .B1(n1307), .C0(n5412), 
        .C1(n16732), .Y(n16962) );
  AOI222XL U2963 ( .A0(n2984), .A1(n16648), .B0(n5487), .B1(n1304), .C0(n5488), 
        .C1(n16417), .Y(n16647) );
  AOI222XL U2964 ( .A0(n3344), .A1(n14758), .B0(n5951), .B1(n1286), .C0(n5952), 
        .C1(n14527), .Y(n14757) );
  AOI222XL U2965 ( .A0(n2741), .A1(n17908), .B0(n5165), .B1(n1316), .C0(n5166), 
        .C1(n17677), .Y(n17907) );
  AOI222XL U2966 ( .A0(n3103), .A1(n16018), .B0(n5639), .B1(n1298), .C0(n5640), 
        .C1(n15787), .Y(n16017) );
  AOI211XL U2967 ( .A0(n5357), .A1(n1311), .B0(n17117), .C0(n17118), .Y(n17116) );
  AOI211XL U2968 ( .A0(n6125), .A1(n1281), .B0(n13967), .C0(n13968), .Y(n13966) );
  AOI211XL U2969 ( .A0(n5003), .A1(n1323), .B0(n18377), .C0(n18378), .Y(n18376) );
  AOI211XL U2970 ( .A0(n5829), .A1(n1293), .B0(n15227), .C0(n15228), .Y(n15226) );
  AOI211XL U2971 ( .A0(n5745), .A1(n1296), .B0(n15542), .C0(n15543), .Y(n15541) );
  AOI211XL U2972 ( .A0(n4887), .A1(n1326), .B0(n18692), .C0(n18693), .Y(n18691) );
  AOI211XL U2973 ( .A0(n5441), .A1(n1308), .B0(n16802), .C0(n16803), .Y(n16801) );
  AOI211XL U2974 ( .A0(n5905), .A1(n1290), .B0(n14912), .C0(n14913), .Y(n14911) );
  AOI211XL U2975 ( .A0(n5517), .A1(n1305), .B0(n16487), .C0(n16488), .Y(n16486) );
  AOI211XL U2976 ( .A0(n5087), .A1(n1320), .B0(n18062), .C0(n18063), .Y(n18061) );
  AOI211XL U2977 ( .A0(n5981), .A1(n1287), .B0(n14597), .C0(n14598), .Y(n14596) );
  AOI211XL U2978 ( .A0(n5593), .A1(n1302), .B0(n16172), .C0(n16173), .Y(n16171) );
  AOI211XL U2979 ( .A0(n5195), .A1(n1317), .B0(n17747), .C0(n17748), .Y(n17746) );
  AOI211XL U2980 ( .A0(n6057), .A1(n1284), .B0(n14282), .C0(n14283), .Y(n14281) );
  AOI211XL U2981 ( .A0(n5669), .A1(n1299), .B0(n15857), .C0(n15858), .Y(n15856) );
  AOI211XL U2982 ( .A0(n5273), .A1(n1314), .B0(n17432), .C0(n17433), .Y(n17431) );
  NAND3XL U2983 ( .A(n9970), .B(n2868), .C(n17205), .Y(n17207) );
  NAND3XL U2984 ( .A(n11138), .B(n2626), .C(n18465), .Y(n18467) );
  NAND3XL U2985 ( .A(n8218), .B(n3228), .C(n15315), .Y(n15317) );
  NAND3XL U2986 ( .A(n8510), .B(n3167), .C(n15630), .Y(n15632) );
  NAND3XL U2987 ( .A(n9678), .B(n2929), .C(n16890), .Y(n16892) );
  NAND3XL U2988 ( .A(n11430), .B(n2565), .C(n18780), .Y(n18782) );
  NAND3XL U2989 ( .A(n7926), .B(n3289), .C(n15000), .Y(n15002) );
  NAND3XL U2990 ( .A(n9386), .B(n2990), .C(n16575), .Y(n16577) );
  NAND3XL U2991 ( .A(n10846), .B(n2688), .C(n18150), .Y(n18152) );
  NAND3XL U2992 ( .A(n7634), .B(n3350), .C(n14685), .Y(n14687) );
  NAND3XL U2993 ( .A(n9094), .B(n3048), .C(n16260), .Y(n16262) );
  NAND3XL U2994 ( .A(n10554), .B(n2748), .C(n17835), .Y(n17837) );
  NAND3XL U2995 ( .A(n7342), .B(n3408), .C(n14370), .Y(n14372) );
  NAND3XL U2996 ( .A(n8802), .B(n3109), .C(n15945), .Y(n15947) );
  NAND3XL U2997 ( .A(n10262), .B(n2808), .C(n17520), .Y(n17522) );
  NAND3XL U2998 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .B(n3470), .C(
        n14055), .Y(n14057) );
  AOI222XL U2999 ( .A0(n994), .A1(n1310), .B0(n17167), .B1(n2889), .C0(n5357), 
        .C1(n1615), .Y(n17166) );
  NAND3XL U3000 ( .A(n2877), .B(n1311), .C(n650), .Y(n17165) );
  AOI222XL U3001 ( .A0(n1133), .A1(n1280), .B0(n14017), .B1(
        top_core_EC_ss_in[1]), .C0(n6125), .C1(n1625), .Y(n14016) );
  NAND3XL U3002 ( .A(n3474), .B(n1281), .C(n649), .Y(n14015) );
  AOI222XL U3003 ( .A0(n938), .A1(n1322), .B0(n18427), .B1(
        top_core_EC_ss_in[113]), .C0(n5003), .C1(n1611), .Y(n18426) );
  NAND3XL U3004 ( .A(n2635), .B(n1323), .C(n651), .Y(n18425) );
  AOI222XL U3005 ( .A0(n1078), .A1(n1292), .B0(n15277), .B1(
        top_core_EC_ss_in[33]), .C0(n5829), .C1(n1621), .Y(n15276) );
  NAND3XL U3006 ( .A(n3233), .B(n1293), .C(n652), .Y(n15275) );
  AOI222XL U3007 ( .A0(n1064), .A1(n1295), .B0(n15592), .B1(n3189), .C0(n5745), 
        .C1(n1620), .Y(n15591) );
  NAND3XL U3008 ( .A(n3172), .B(n1296), .C(n653), .Y(n15590) );
  AOI222XL U3009 ( .A0(n924), .A1(n1325), .B0(n18742), .B1(n2587), .C0(n4887), 
        .C1(n1610), .Y(n18741) );
  NAND3XL U3010 ( .A(n2574), .B(n1326), .C(n654), .Y(n18740) );
  AOI222XL U3011 ( .A0(n1008), .A1(n1307), .B0(n16852), .B1(
        top_core_EC_ss_in[73]), .C0(n5441), .C1(n1616), .Y(n16851) );
  NAND3XL U3012 ( .A(n2938), .B(n1308), .C(n655), .Y(n16850) );
  AOI222XL U3013 ( .A0(n1092), .A1(n1289), .B0(n14962), .B1(n3310), .C0(n5905), 
        .C1(n1622), .Y(n14961) );
  NAND3XL U3014 ( .A(n3296), .B(n1290), .C(n656), .Y(n14960) );
  AOI222XL U3015 ( .A0(n1022), .A1(n1304), .B0(n16537), .B1(n3011), .C0(n5517), 
        .C1(n1617), .Y(n16536) );
  NAND3XL U3016 ( .A(n2999), .B(n1305), .C(n657), .Y(n16535) );
  AOI222XL U3017 ( .A0(n952), .A1(n1319), .B0(n18112), .B1(
        top_core_EC_ss_in[105]), .C0(n5087), .C1(n1612), .Y(n18111) );
  NAND3XL U3018 ( .A(n2696), .B(n1320), .C(n658), .Y(n18110) );
  AOI222XL U3019 ( .A0(n1106), .A1(n1286), .B0(n14647), .B1(n3372), .C0(n5981), 
        .C1(n1623), .Y(n14646) );
  NAND3XL U3020 ( .A(n3355), .B(n1287), .C(n659), .Y(n14645) );
  AOI222XL U3021 ( .A0(n1036), .A1(n1301), .B0(n16222), .B1(
        top_core_EC_ss_in[57]), .C0(n5593), .C1(n1618), .Y(n16221) );
  NAND3XL U3022 ( .A(n3057), .B(n1302), .C(n660), .Y(n16220) );
  AOI222XL U3023 ( .A0(n966), .A1(n1316), .B0(n17797), .B1(n2769), .C0(n5195), 
        .C1(n1613), .Y(n17796) );
  NAND3XL U3024 ( .A(n2752), .B(n1317), .C(n661), .Y(n17795) );
  AOI222XL U3025 ( .A0(n1120), .A1(n1283), .B0(n14332), .B1(
        top_core_EC_ss_in[9]), .C0(n6057), .C1(n1624), .Y(n14331) );
  NAND3XL U3026 ( .A(n3417), .B(n1284), .C(n662), .Y(n14330) );
  AOI222XL U3027 ( .A0(n1050), .A1(n1298), .B0(n15907), .B1(n3131), .C0(n5669), 
        .C1(n1619), .Y(n15906) );
  NAND3XL U3028 ( .A(n3118), .B(n1299), .C(n663), .Y(n15905) );
  AOI222XL U3029 ( .A0(n980), .A1(n1313), .B0(n17482), .B1(
        top_core_EC_ss_in[89]), .C0(n5273), .C1(n1614), .Y(n17481) );
  NAND3XL U3030 ( .A(n2815), .B(n1314), .C(n664), .Y(n17480) );
  AOI222XL U3031 ( .A0(n5357), .A1(n1310), .B0(n17057), .B1(n465), .C0(n5380), 
        .C1(n1002), .Y(n17145) );
  AOI222XL U3032 ( .A0(n6125), .A1(n1280), .B0(n13907), .B1(n466), .C0(n6151), 
        .C1(n1141), .Y(n13995) );
  AOI222XL U3033 ( .A0(n5003), .A1(n1322), .B0(n18317), .B1(n467), .C0(n5026), 
        .C1(n946), .Y(n18405) );
  AOI222XL U3034 ( .A0(n5829), .A1(n1292), .B0(n15167), .B1(n468), .C0(n5852), 
        .C1(n1086), .Y(n15255) );
  AOI222XL U3035 ( .A0(n5745), .A1(n1295), .B0(n15482), .B1(n469), .C0(n5768), 
        .C1(n1072), .Y(n15570) );
  AOI222XL U3036 ( .A0(n4887), .A1(n1325), .B0(n18632), .B1(n471), .C0(n4910), 
        .C1(n932), .Y(n18720) );
  AOI222XL U3037 ( .A0(n5441), .A1(n1307), .B0(n16742), .B1(n470), .C0(n5464), 
        .C1(n1016), .Y(n16830) );
  AOI222XL U3038 ( .A0(n5905), .A1(n1289), .B0(n14852), .B1(n472), .C0(n5928), 
        .C1(n1100), .Y(n14940) );
  AOI222XL U3039 ( .A0(n5517), .A1(n1304), .B0(n16427), .B1(n473), .C0(n5540), 
        .C1(n1030), .Y(n16515) );
  AOI222XL U3040 ( .A0(n5087), .A1(n1319), .B0(n18002), .B1(n474), .C0(n5110), 
        .C1(n960), .Y(n18090) );
  AOI222XL U3041 ( .A0(n5981), .A1(n1286), .B0(n14537), .B1(n475), .C0(n6004), 
        .C1(n1114), .Y(n14625) );
  AOI222XL U3042 ( .A0(n5593), .A1(n1301), .B0(n16112), .B1(n476), .C0(n5616), 
        .C1(n1044), .Y(n16200) );
  AOI222XL U3043 ( .A0(n5195), .A1(n1316), .B0(n17687), .B1(n477), .C0(n5218), 
        .C1(n974), .Y(n17775) );
  AOI222XL U3044 ( .A0(n6057), .A1(n1283), .B0(n14222), .B1(n478), .C0(n6080), 
        .C1(n1128), .Y(n14310) );
  AOI222XL U3045 ( .A0(n5669), .A1(n1298), .B0(n15797), .B1(n479), .C0(n5692), 
        .C1(n1058), .Y(n15885) );
  AOI222XL U3046 ( .A0(n5273), .A1(n1313), .B0(n17372), .B1(n480), .C0(n5296), 
        .C1(n988), .Y(n17460) );
  AOI32XL U3047 ( .A0(n2758), .A1(n2749), .A2(n2772), .B0(n17797), .B1(n17647), 
        .Y(n17892) );
  AOI32XL U3048 ( .A0(n2993), .A1(n2992), .A2(n3015), .B0(n16537), .B1(n16387), 
        .Y(n16632) );
  AOI32XL U3049 ( .A0(n3361), .A1(n3352), .A2(n3375), .B0(n14647), .B1(n14497), 
        .Y(n14742) );
  AOI32XL U3050 ( .A0(n3120), .A1(n3111), .A2(n3134), .B0(n15907), .B1(n15757), 
        .Y(n16002) );
  AOI32XL U3051 ( .A0(n3473), .A1(n3471), .A2(n3494), .B0(n14017), .B1(n13867), 
        .Y(n14112) );
  AOI32XL U3052 ( .A0(n2879), .A1(n2870), .A2(n2893), .B0(n17167), .B1(n17017), 
        .Y(n17262) );
  AOI32XL U3053 ( .A0(n2637), .A1(n2628), .A2(n2650), .B0(n18427), .B1(n18277), 
        .Y(n18522) );
  AOI32XL U3054 ( .A0(n3239), .A1(n3230), .A2(n3253), .B0(n15277), .B1(n15127), 
        .Y(n15372) );
  AOI32XL U3055 ( .A0(n3178), .A1(n3169), .A2(n3192), .B0(n15592), .B1(n15442), 
        .Y(n15687) );
  AOI32XL U3056 ( .A0(n2576), .A1(n2567), .A2(n2590), .B0(n18742), .B1(n18592), 
        .Y(n18837) );
  AOI32XL U3057 ( .A0(n2932), .A1(n2931), .A2(n2954), .B0(n16852), .B1(n16702), 
        .Y(n16947) );
  AOI32XL U3058 ( .A0(n3293), .A1(n3291), .A2(n3314), .B0(n14962), .B1(n14812), 
        .Y(n15057) );
  AOI32XL U3059 ( .A0(n2690), .A1(n2689), .A2(n2711), .B0(n18112), .B1(n17962), 
        .Y(n18207) );
  AOI32XL U3060 ( .A0(n3059), .A1(n3050), .A2(n3072), .B0(n16222), .B1(n16072), 
        .Y(n16317) );
  AOI32XL U3061 ( .A0(n3411), .A1(n3410), .A2(n3433), .B0(n14332), .B1(n14182), 
        .Y(n14427) );
  AOI32XL U3062 ( .A0(n2812), .A1(n2810), .A2(n2833), .B0(n17482), .B1(n17332), 
        .Y(n17577) );
  AOI22XL U3063 ( .A0(n722), .A1(n2899), .B0(n5375), .B1(n9900), .Y(n10162) );
  AOI22XL U3064 ( .A0(n723), .A1(n3495), .B0(n6165), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n348) );
  AOI22XL U3065 ( .A0(n725), .A1(n3259), .B0(n5847), .B1(n8148), .Y(n8410) );
  AOI22XL U3066 ( .A0(n724), .A1(n2662), .B0(n5021), .B1(n11068), .Y(n11330)
         );
  AOI22XL U3067 ( .A0(n731), .A1(n2712), .B0(n5105), .B1(n10776), .Y(n11038)
         );
  AOI22XL U3068 ( .A0(n735), .A1(n3434), .B0(n6075), .B1(n7272), .Y(n7534) );
  AOI22XL U3069 ( .A0(n733), .A1(n3084), .B0(n5611), .B1(n9024), .Y(n9286) );
  AOI22XL U3070 ( .A0(n737), .A1(n2836), .B0(n5291), .B1(n10192), .Y(n10454)
         );
  AOI22XL U3071 ( .A0(n730), .A1(n3017), .B0(n5535), .B1(n9316), .Y(n9578) );
  AOI22XL U3072 ( .A0(n726), .A1(n3198), .B0(n5763), .B1(n8440), .Y(n8702) );
  AOI22XL U3073 ( .A0(n732), .A1(n3377), .B0(n5999), .B1(n7564), .Y(n7826) );
  AOI22XL U3074 ( .A0(n728), .A1(n2601), .B0(n4905), .B1(n11360), .Y(n11622)
         );
  AOI22XL U3075 ( .A0(n734), .A1(n2775), .B0(n5213), .B1(n10484), .Y(n10746)
         );
  AOI22XL U3076 ( .A0(n727), .A1(n2960), .B0(n5459), .B1(n9608), .Y(n9870) );
  AOI22XL U3077 ( .A0(n736), .A1(n3136), .B0(n5687), .B1(n8732), .Y(n8994) );
  AOI22XL U3078 ( .A0(n729), .A1(n3316), .B0(n5923), .B1(n7856), .Y(n8118) );
  AOI22XL U3079 ( .A0(n13918), .A1(n1281), .B0(n14033), .B1(n514), .Y(n14117)
         );
  AOI22XL U3080 ( .A0(n17068), .A1(n1311), .B0(n17183), .B1(n513), .Y(n17267)
         );
  AOI22XL U3081 ( .A0(n18328), .A1(n1323), .B0(n18443), .B1(n515), .Y(n18527)
         );
  AOI22XL U3082 ( .A0(n15178), .A1(n1293), .B0(n15293), .B1(n516), .Y(n15377)
         );
  AOI22XL U3083 ( .A0(n15493), .A1(n1296), .B0(n15608), .B1(n517), .Y(n15692)
         );
  AOI22XL U3084 ( .A0(n18643), .A1(n1326), .B0(n18758), .B1(n518), .Y(n18842)
         );
  AOI22XL U3085 ( .A0(n16753), .A1(n1308), .B0(n16868), .B1(n519), .Y(n16952)
         );
  AOI22XL U3086 ( .A0(n14863), .A1(n1290), .B0(n14978), .B1(n520), .Y(n15062)
         );
  AOI22XL U3087 ( .A0(n16438), .A1(n1305), .B0(n16553), .B1(n521), .Y(n16637)
         );
  AOI22XL U3088 ( .A0(n18013), .A1(n1320), .B0(n18128), .B1(n522), .Y(n18212)
         );
  AOI22XL U3089 ( .A0(n14548), .A1(n1287), .B0(n14663), .B1(n523), .Y(n14747)
         );
  AOI22XL U3090 ( .A0(n16123), .A1(n1302), .B0(n16238), .B1(n524), .Y(n16322)
         );
  AOI22XL U3091 ( .A0(n17698), .A1(n1317), .B0(n17813), .B1(n525), .Y(n17897)
         );
  AOI22XL U3092 ( .A0(n14233), .A1(n1284), .B0(n14348), .B1(n526), .Y(n14432)
         );
  AOI22XL U3093 ( .A0(n15808), .A1(n1299), .B0(n15923), .B1(n527), .Y(n16007)
         );
  AOI22XL U3094 ( .A0(n17383), .A1(n1314), .B0(n17498), .B1(n528), .Y(n17582)
         );
  OAI211XL U3095 ( .A0(n17073), .A1(n1309), .B0(n17077), .C0(n17160), .Y(
        n17159) );
  OAI211XL U3096 ( .A0(n13923), .A1(n1279), .B0(n13927), .C0(n14010), .Y(
        n14009) );
  OAI211XL U3097 ( .A0(n18333), .A1(n1321), .B0(n18337), .C0(n18420), .Y(
        n18419) );
  OAI211XL U3098 ( .A0(n15183), .A1(n1291), .B0(n15187), .C0(n15270), .Y(
        n15269) );
  OAI211XL U3099 ( .A0(n15498), .A1(n1294), .B0(n15502), .C0(n15585), .Y(
        n15584) );
  OAI211XL U3100 ( .A0(n18648), .A1(n1324), .B0(n18652), .C0(n18735), .Y(
        n18734) );
  OAI211XL U3101 ( .A0(n16758), .A1(n1306), .B0(n16762), .C0(n16845), .Y(
        n16844) );
  OAI211XL U3102 ( .A0(n14868), .A1(n1288), .B0(n14872), .C0(n14955), .Y(
        n14954) );
  OAI211XL U3103 ( .A0(n16443), .A1(n1303), .B0(n16447), .C0(n16530), .Y(
        n16529) );
  OAI211XL U3104 ( .A0(n18018), .A1(n1318), .B0(n18022), .C0(n18105), .Y(
        n18104) );
  OAI211XL U3105 ( .A0(n14553), .A1(n1285), .B0(n14557), .C0(n14640), .Y(
        n14639) );
  OAI211XL U3106 ( .A0(n16128), .A1(n1300), .B0(n16132), .C0(n16215), .Y(
        n16214) );
  OAI211XL U3107 ( .A0(n17703), .A1(n1315), .B0(n17707), .C0(n17790), .Y(
        n17789) );
  OAI211XL U3108 ( .A0(n14238), .A1(n1282), .B0(n14242), .C0(n14325), .Y(
        n14324) );
  OAI211XL U3109 ( .A0(n15813), .A1(n1297), .B0(n15817), .C0(n15900), .Y(
        n15899) );
  OAI211XL U3110 ( .A0(n17388), .A1(n1312), .B0(n17392), .C0(n17475), .Y(
        n17474) );
  AOI22XL U3111 ( .A0(n1805), .A1(n745), .B0(n11651), .B1(n1202), .Y(n11690)
         );
  AOI22XL U3112 ( .A0(n1826), .A1(n746), .B0(top_core_KE_sb1_n76), .B1(n1193), 
        .Y(top_core_KE_sb1_n115) );
  AOI22XL U3113 ( .A0(n1766), .A1(n744), .B0(n12283), .B1(n1162), .Y(n12321)
         );
  AOI22XL U3114 ( .A0(n1784), .A1(n747), .B0(n11967), .B1(n1153), .Y(n12006)
         );
  AOI22XL U3115 ( .A0(n1683), .A1(n1151), .B0(n13228), .B1(n1148), .Y(n13267)
         );
  AOI22XL U3116 ( .A0(n1712), .A1(n1200), .B0(n12913), .B1(n1197), .Y(n12952)
         );
  AOI22XL U3117 ( .A0(n1741), .A1(n1191), .B0(n12598), .B1(n1188), .Y(n12637)
         );
  AOI22XL U3118 ( .A0(n1653), .A1(n1160), .B0(n13543), .B1(n1157), .Y(n13582)
         );
  AOI222XL U3119 ( .A0(n1625), .A1(n1140), .B0(n3504), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n174), .C0(n6166), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n311) );
  AOI222XL U3120 ( .A0(n1615), .A1(n1000), .B0(top_core_EC_ss_in[80]), .B1(
        n9988), .C0(n5376), .C1(n9970), .Y(n10125) );
  AOI222XL U3121 ( .A0(n1611), .A1(n944), .B0(n2651), .B1(n11156), .C0(n5022), 
        .C1(n11138), .Y(n11293) );
  AOI222XL U3122 ( .A0(n1621), .A1(n1084), .B0(top_core_EC_ss_in[32]), .B1(
        n8236), .C0(n5848), .C1(n8218), .Y(n8373) );
  AOI222XL U3123 ( .A0(n1612), .A1(n958), .B0(n2721), .B1(n10864), .C0(n5106), 
        .C1(n10846), .Y(n11001) );
  AOI222XL U3124 ( .A0(n1618), .A1(n1042), .B0(n3073), .B1(n9112), .C0(n5612), 
        .C1(n9094), .Y(n9249) );
  AOI222XL U3125 ( .A0(n1624), .A1(n1126), .B0(n3443), .B1(n7360), .C0(n6076), 
        .C1(n7342), .Y(n7497) );
  AOI222XL U3126 ( .A0(n1614), .A1(n986), .B0(n2834), .B1(n10280), .C0(n5292), 
        .C1(n10262), .Y(n10417) );
  AOI222XL U3127 ( .A0(n1617), .A1(n1028), .B0(n3016), .B1(n9404), .C0(n5536), 
        .C1(n9386), .Y(n9541) );
  AOI222XL U3128 ( .A0(n1620), .A1(n1070), .B0(top_core_EC_ss_in[40]), .B1(
        n8528), .C0(n5764), .C1(n8510), .Y(n8665) );
  AOI222XL U3129 ( .A0(n1623), .A1(n1112), .B0(n3376), .B1(n7652), .C0(n6000), 
        .C1(n7634), .Y(n7789) );
  AOI222XL U3130 ( .A0(n1610), .A1(n930), .B0(n2590), .B1(n11448), .C0(n4906), 
        .C1(n11430), .Y(n11585) );
  AOI222XL U3131 ( .A0(n1613), .A1(n972), .B0(n2773), .B1(n10572), .C0(n5214), 
        .C1(n10554), .Y(n10709) );
  AOI222XL U3132 ( .A0(n1616), .A1(n1014), .B0(top_core_EC_ss_in[72]), .B1(
        n9696), .C0(n5460), .C1(n9678), .Y(n9833) );
  AOI222XL U3133 ( .A0(n1619), .A1(n1056), .B0(n3135), .B1(n8820), .C0(n5688), 
        .C1(n8802), .Y(n8957) );
  AOI222XL U3134 ( .A0(n1622), .A1(n1098), .B0(n3324), .B1(n7944), .C0(n5924), 
        .C1(n7926), .Y(n8081) );
  AOI211XL U3135 ( .A0(n562), .A1(n9900), .B0(n10030), .C0(n10031), .Y(n10029)
         );
  AOI211XL U3136 ( .A0(n561), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n216), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n217), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n215) );
  AOI211XL U3137 ( .A0(n563), .A1(n11068), .B0(n11198), .C0(n11199), .Y(n11197) );
  AOI211XL U3138 ( .A0(n564), .A1(n8148), .B0(n8278), .C0(n8279), .Y(n8277) );
  AOI211XL U3139 ( .A0(n565), .A1(n10776), .B0(n10906), .C0(n10907), .Y(n10905) );
  AOI211XL U3140 ( .A0(n566), .A1(n9024), .B0(n9154), .C0(n9155), .Y(n9153) );
  AOI211XL U3141 ( .A0(n567), .A1(n7272), .B0(n7402), .C0(n7403), .Y(n7401) );
  AOI211XL U3142 ( .A0(n568), .A1(n10192), .B0(n10322), .C0(n10323), .Y(n10321) );
  AOI211XL U3143 ( .A0(n569), .A1(n9316), .B0(n9446), .C0(n9447), .Y(n9445) );
  AOI211XL U3144 ( .A0(n570), .A1(n8440), .B0(n8570), .C0(n8571), .Y(n8569) );
  AOI211XL U3145 ( .A0(n571), .A1(n7564), .B0(n7694), .C0(n7695), .Y(n7693) );
  AOI211XL U3146 ( .A0(n572), .A1(n11360), .B0(n11490), .C0(n11491), .Y(n11489) );
  AOI211XL U3147 ( .A0(n573), .A1(n10484), .B0(n10614), .C0(n10615), .Y(n10613) );
  AOI211XL U3148 ( .A0(n574), .A1(n9608), .B0(n9738), .C0(n9739), .Y(n9737) );
  AOI211XL U3149 ( .A0(n575), .A1(n8732), .B0(n8862), .C0(n8863), .Y(n8861) );
  AOI211XL U3150 ( .A0(n576), .A1(n7856), .B0(n7986), .C0(n7987), .Y(n7985) );
  AOI211XL U3151 ( .A0(n5371), .A1(n9970), .B0(n9986), .C0(n9987), .Y(n9984)
         );
  AOI211XL U3152 ( .A0(n6161), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n172), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n173), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n170) );
  AOI211XL U3153 ( .A0(n5017), .A1(n11138), .B0(n11154), .C0(n11155), .Y(
        n11152) );
  AOI211XL U3154 ( .A0(n5843), .A1(n8218), .B0(n8234), .C0(n8235), .Y(n8232)
         );
  AOI211XL U3155 ( .A0(n5101), .A1(n10846), .B0(n10862), .C0(n10863), .Y(
        n10860) );
  AOI211XL U3156 ( .A0(n5607), .A1(n9094), .B0(n9110), .C0(n9111), .Y(n9108)
         );
  AOI211XL U3157 ( .A0(n6071), .A1(n7342), .B0(n7358), .C0(n7359), .Y(n7356)
         );
  AOI211XL U3158 ( .A0(n5287), .A1(n10262), .B0(n10278), .C0(n10279), .Y(
        n10276) );
  AOI211XL U3159 ( .A0(n5531), .A1(n9386), .B0(n9402), .C0(n9403), .Y(n9400)
         );
  AOI211XL U3160 ( .A0(n5759), .A1(n8510), .B0(n8526), .C0(n8527), .Y(n8524)
         );
  AOI211XL U3161 ( .A0(n5995), .A1(n7634), .B0(n7650), .C0(n7651), .Y(n7648)
         );
  AOI211XL U3162 ( .A0(n4901), .A1(n11430), .B0(n11446), .C0(n11447), .Y(
        n11444) );
  AOI211XL U3163 ( .A0(n5209), .A1(n10554), .B0(n10570), .C0(n10571), .Y(
        n10568) );
  AOI211XL U3164 ( .A0(n5455), .A1(n9678), .B0(n9694), .C0(n9695), .Y(n9692)
         );
  AOI211XL U3165 ( .A0(n5683), .A1(n8802), .B0(n8818), .C0(n8819), .Y(n8816)
         );
  AOI211XL U3166 ( .A0(n5919), .A1(n7926), .B0(n7942), .C0(n7943), .Y(n7940)
         );
  AOI31XL U3167 ( .A0(n15432), .A1(n1070), .A2(n15433), .B0(n15434), .Y(n15426) );
  AOI31XL U3168 ( .A0(n17952), .A1(n958), .A2(n17953), .B0(n17954), .Y(n17946)
         );
  AOI31XL U3169 ( .A0(n14172), .A1(n1126), .A2(n14173), .B0(n14174), .Y(n14166) );
  AOI31XL U3170 ( .A0(n18582), .A1(n930), .A2(n18583), .B0(n18584), .Y(n18576)
         );
  AOI31XL U3171 ( .A0(n14802), .A1(n1098), .A2(n14803), .B0(n14804), .Y(n14796) );
  AOI31XL U3172 ( .A0(n16062), .A1(n1042), .A2(n16063), .B0(n16064), .Y(n16056) );
  AOI31XL U3173 ( .A0(n17322), .A1(n986), .A2(n17323), .B0(n17324), .Y(n17316)
         );
  AOI31XL U3174 ( .A0(n13857), .A1(n1140), .A2(n13858), .B0(n13859), .Y(n13851) );
  AOI31XL U3175 ( .A0(n17007), .A1(n1000), .A2(n17008), .B0(n17009), .Y(n17001) );
  AOI31XL U3176 ( .A0(n18267), .A1(n944), .A2(n18268), .B0(n18269), .Y(n18261)
         );
  AOI31XL U3177 ( .A0(n15117), .A1(n1084), .A2(n15118), .B0(n15119), .Y(n15111) );
  AOI31XL U3178 ( .A0(n16692), .A1(n1014), .A2(n16693), .B0(n16694), .Y(n16686) );
  AOI31XL U3179 ( .A0(n16377), .A1(n1028), .A2(n16378), .B0(n16379), .Y(n16371) );
  AOI31XL U3180 ( .A0(n14487), .A1(n1112), .A2(n14488), .B0(n14489), .Y(n14481) );
  AOI31XL U3181 ( .A0(n17637), .A1(n972), .A2(n17638), .B0(n17639), .Y(n17631)
         );
  AOI31XL U3182 ( .A0(n15747), .A1(n1056), .A2(n15748), .B0(n15749), .Y(n15741) );
  AOI22XL U3183 ( .A0(n634), .A1(n3498), .B0(n1134), .B1(n13911), .Y(n14105)
         );
  AOI22XL U3184 ( .A0(n633), .A1(n2900), .B0(n995), .B1(n17061), .Y(n17255) );
  AOI22XL U3185 ( .A0(n635), .A1(n2663), .B0(n939), .B1(n18321), .Y(n18515) );
  AOI22XL U3186 ( .A0(n636), .A1(n3260), .B0(n1079), .B1(n15171), .Y(n15365)
         );
  AOI22XL U3187 ( .A0(n637), .A1(n3199), .B0(n1065), .B1(n15486), .Y(n15680)
         );
  AOI22XL U3188 ( .A0(n638), .A1(n2602), .B0(n925), .B1(n18636), .Y(n18830) );
  AOI22XL U3189 ( .A0(n639), .A1(n2961), .B0(n1009), .B1(n16746), .Y(n16940)
         );
  AOI22XL U3190 ( .A0(n640), .A1(n3315), .B0(n1093), .B1(n14856), .Y(n15050)
         );
  AOI22XL U3191 ( .A0(n641), .A1(n3025), .B0(n1023), .B1(n16431), .Y(n16625)
         );
  AOI22XL U3192 ( .A0(n642), .A1(n2716), .B0(n953), .B1(n18006), .Y(n18200) );
  AOI22XL U3193 ( .A0(n643), .A1(n3385), .B0(n1107), .B1(n14541), .Y(n14735)
         );
  AOI22XL U3194 ( .A0(n644), .A1(n3085), .B0(n1037), .B1(n16116), .Y(n16310)
         );
  AOI22XL U3195 ( .A0(n645), .A1(n2774), .B0(n967), .B1(n17691), .Y(n17885) );
  AOI22XL U3196 ( .A0(n646), .A1(n3438), .B0(n1121), .B1(n14226), .Y(n14420)
         );
  AOI22XL U3197 ( .A0(n647), .A1(n3144), .B0(n1051), .B1(n15801), .Y(n15995)
         );
  AOI22XL U3198 ( .A0(n648), .A1(n2835), .B0(n981), .B1(n17376), .Y(n17570) );
  AOI211XL U3199 ( .A0(n1625), .A1(n3473), .B0(n6135), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n106), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n105) );
  AOI211XL U3200 ( .A0(n1203), .A1(n1257), .B0(n11681), .C0(n11664), .Y(n11678) );
  AOI211XL U3201 ( .A0(n1194), .A1(n1329), .B0(top_core_KE_sb1_n106), .C0(
        top_core_KE_sb1_n89), .Y(top_core_KE_sb1_n103) );
  AOI211XL U3202 ( .A0(n1154), .A1(n1260), .B0(n11997), .C0(n11980), .Y(n11994) );
  AOI211XL U3203 ( .A0(n1133), .A1(n13857), .B0(n14023), .C0(n6126), .Y(n14099) );
  AOI211XL U3204 ( .A0(n994), .A1(n17007), .B0(n17173), .C0(n5358), .Y(n17249)
         );
  AOI211XL U3205 ( .A0(n938), .A1(n18267), .B0(n18433), .C0(n5004), .Y(n18509)
         );
  AOI211XL U3206 ( .A0(n1078), .A1(n15117), .B0(n15283), .C0(n5830), .Y(n15359) );
  AOI211XL U3207 ( .A0(n1064), .A1(n15432), .B0(n15598), .C0(n5746), .Y(n15674) );
  AOI211XL U3208 ( .A0(n924), .A1(n18582), .B0(n18748), .C0(n4888), .Y(n18824)
         );
  AOI211XL U3209 ( .A0(n1008), .A1(n16692), .B0(n16858), .C0(n5442), .Y(n16934) );
  AOI211XL U3210 ( .A0(n1092), .A1(n14802), .B0(n14968), .C0(n5906), .Y(n15044) );
  AOI211XL U3211 ( .A0(n1022), .A1(n16377), .B0(n16543), .C0(n5518), .Y(n16619) );
  AOI211XL U3212 ( .A0(n952), .A1(n17952), .B0(n18118), .C0(n5088), .Y(n18194)
         );
  AOI211XL U3213 ( .A0(n1106), .A1(n14487), .B0(n14653), .C0(n5982), .Y(n14729) );
  AOI211XL U3214 ( .A0(n1036), .A1(n16062), .B0(n16228), .C0(n5594), .Y(n16304) );
  AOI211XL U3215 ( .A0(n966), .A1(n17637), .B0(n17803), .C0(n5196), .Y(n17879)
         );
  AOI211XL U3216 ( .A0(n1120), .A1(n14172), .B0(n14338), .C0(n6058), .Y(n14414) );
  AOI211XL U3217 ( .A0(n1050), .A1(n15747), .B0(n15913), .C0(n5670), .Y(n15989) );
  AOI211XL U3218 ( .A0(n980), .A1(n17322), .B0(n17488), .C0(n5274), .Y(n17564)
         );
  AOI211XL U3219 ( .A0(n1163), .A1(n1263), .B0(n12312), .C0(n12295), .Y(n12309) );
  AOI211XL U3220 ( .A0(n5378), .A1(n17007), .B0(n17069), .C0(n17070), .Y(
        n17066) );
  OAI31XL U3221 ( .A0(n17047), .A1(n2867), .A2(n2873), .B0(n17071), .Y(n17070)
         );
  AOI211XL U3222 ( .A0(n6149), .A1(n13857), .B0(n13919), .C0(n13920), .Y(
        n13916) );
  OAI31XL U3223 ( .A0(n13897), .A1(n3468), .A2(n3475), .B0(n13921), .Y(n13920)
         );
  AOI211XL U3224 ( .A0(n5024), .A1(n18267), .B0(n18329), .C0(n18330), .Y(
        n18326) );
  OAI31XL U3225 ( .A0(n18307), .A1(n2625), .A2(n2631), .B0(n18331), .Y(n18330)
         );
  AOI211XL U3226 ( .A0(n5850), .A1(n15117), .B0(n15179), .C0(n15180), .Y(
        n15176) );
  OAI31XL U3227 ( .A0(n15157), .A1(n3227), .A2(n3234), .B0(n15181), .Y(n15180)
         );
  AOI211XL U3228 ( .A0(n5766), .A1(n15432), .B0(n15494), .C0(n15495), .Y(
        n15491) );
  OAI31XL U3229 ( .A0(n15472), .A1(n3166), .A2(n3173), .B0(n15496), .Y(n15495)
         );
  AOI211XL U3230 ( .A0(n4908), .A1(n18582), .B0(n18644), .C0(n18645), .Y(
        n18641) );
  OAI31XL U3231 ( .A0(n18622), .A1(n2564), .A2(n2570), .B0(n18646), .Y(n18645)
         );
  AOI211XL U3232 ( .A0(n5462), .A1(n16692), .B0(n16754), .C0(n16755), .Y(
        n16751) );
  OAI31XL U3233 ( .A0(n16732), .A1(n2928), .A2(n2934), .B0(n16756), .Y(n16755)
         );
  AOI211XL U3234 ( .A0(n5926), .A1(n14802), .B0(n14864), .C0(n14865), .Y(
        n14861) );
  OAI31XL U3235 ( .A0(n14842), .A1(n3288), .A2(n3294), .B0(n14866), .Y(n14865)
         );
  AOI211XL U3236 ( .A0(n5538), .A1(n16377), .B0(n16439), .C0(n16440), .Y(
        n16436) );
  OAI31XL U3237 ( .A0(n16417), .A1(n2989), .A2(n2995), .B0(n16441), .Y(n16440)
         );
  AOI211XL U3238 ( .A0(n5108), .A1(n17952), .B0(n18014), .C0(n18015), .Y(
        n18011) );
  OAI31XL U3239 ( .A0(n17992), .A1(n2686), .A2(n2692), .B0(n18016), .Y(n18015)
         );
  AOI211XL U3240 ( .A0(n6002), .A1(n14487), .B0(n14549), .C0(n14550), .Y(
        n14546) );
  OAI31XL U3241 ( .A0(n14527), .A1(n3349), .A2(n3356), .B0(n14551), .Y(n14550)
         );
  AOI211XL U3242 ( .A0(n5614), .A1(n16062), .B0(n16124), .C0(n16125), .Y(
        n16121) );
  OAI31XL U3243 ( .A0(n16102), .A1(n3047), .A2(n3053), .B0(n16126), .Y(n16125)
         );
  AOI211XL U3244 ( .A0(n5216), .A1(n17637), .B0(n17699), .C0(n17700), .Y(
        n17696) );
  OAI31XL U3245 ( .A0(n17677), .A1(n2746), .A2(n2753), .B0(n17701), .Y(n17700)
         );
  AOI211XL U3246 ( .A0(n6078), .A1(n14172), .B0(n14234), .C0(n14235), .Y(
        n14231) );
  OAI31XL U3247 ( .A0(n14212), .A1(n3407), .A2(n3413), .B0(n14236), .Y(n14235)
         );
  AOI211XL U3248 ( .A0(n5690), .A1(n15747), .B0(n15809), .C0(n15810), .Y(
        n15806) );
  OAI31XL U3249 ( .A0(n15787), .A1(n3108), .A2(n3114), .B0(n15811), .Y(n15810)
         );
  AOI211XL U3250 ( .A0(n5294), .A1(n17322), .B0(n17384), .C0(n17385), .Y(
        n17381) );
  OAI31XL U3251 ( .A0(n17362), .A1(n2807), .A2(n2813), .B0(n17386), .Y(n17385)
         );
  AOI22XL U3252 ( .A0(n1152), .A1(n13238), .B0(n1149), .B1(n1680), .Y(n13356)
         );
  AOI211XL U3253 ( .A0(n1158), .A1(n1276), .B0(n13573), .C0(n13556), .Y(n13570) );
  AOI211XL U3254 ( .A0(n6132), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n317), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n318), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n313) );
  AOI211XL U3255 ( .A0(n5336), .A1(n9891), .B0(n10131), .C0(n10132), .Y(n10127) );
  AOI211XL U3256 ( .A0(n4982), .A1(n11059), .B0(n11299), .C0(n11300), .Y(
        n11295) );
  AOI211XL U3257 ( .A0(n5808), .A1(n8139), .B0(n8379), .C0(n8380), .Y(n8375)
         );
  AOI211XL U3258 ( .A0(n5066), .A1(n10767), .B0(n11007), .C0(n11008), .Y(
        n11003) );
  AOI211XL U3259 ( .A0(n5572), .A1(n9015), .B0(n9255), .C0(n9256), .Y(n9251)
         );
  AOI211XL U3260 ( .A0(n6036), .A1(n7263), .B0(n7503), .C0(n7504), .Y(n7499)
         );
  AOI211XL U3261 ( .A0(n5252), .A1(n10183), .B0(n10423), .C0(n10424), .Y(
        n10419) );
  AOI211XL U3262 ( .A0(n5496), .A1(n9307), .B0(n9547), .C0(n9548), .Y(n9543)
         );
  AOI211XL U3263 ( .A0(n5724), .A1(n8431), .B0(n8671), .C0(n8672), .Y(n8667)
         );
  AOI211XL U3264 ( .A0(n5960), .A1(n7555), .B0(n7795), .C0(n7796), .Y(n7791)
         );
  AOI211XL U3265 ( .A0(n4866), .A1(n11351), .B0(n11591), .C0(n11592), .Y(
        n11587) );
  AOI211XL U3266 ( .A0(n5174), .A1(n10475), .B0(n10715), .C0(n10716), .Y(
        n10711) );
  AOI211XL U3267 ( .A0(n5420), .A1(n9599), .B0(n9839), .C0(n9840), .Y(n9835)
         );
  AOI211XL U3268 ( .A0(n5648), .A1(n8723), .B0(n8963), .C0(n8964), .Y(n8959)
         );
  AOI211XL U3269 ( .A0(n5884), .A1(n7847), .B0(n8087), .C0(n8088), .Y(n8083)
         );
  AOI211XL U3270 ( .A0(n11641), .A1(n11691), .B0(n11681), .C0(n6911), .Y(
        n11838) );
  AOI211XL U3271 ( .A0(top_core_KE_sb1_n66), .A1(top_core_KE_sb1_n116), .B0(
        top_core_KE_sb1_n106), .C0(n6865), .Y(top_core_KE_sb1_n267) );
  AOI211XL U3272 ( .A0(n12273), .A1(n12322), .B0(n12312), .C0(n6618), .Y(
        n12469) );
  AOI211XL U3273 ( .A0(n11957), .A1(n12007), .B0(n11997), .C0(n6571), .Y(
        n12154) );
  AOI211XL U3274 ( .A0(n1149), .A1(n1273), .B0(n13258), .C0(n13241), .Y(n13255) );
  AOI211XL U3275 ( .A0(n1198), .A1(n1270), .B0(n12943), .C0(n12926), .Y(n12940) );
  AOI211XL U3276 ( .A0(n1189), .A1(n1267), .B0(n12628), .C0(n12611), .Y(n12625) );
  NAND2XL U3277 ( .A(n10795), .B(n10765), .Y(n10830) );
  NAND2XL U3278 ( .A(n9919), .B(n9889), .Y(n9954) );
  NAND2XL U3279 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n104), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n71), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n139) );
  NAND2XL U3280 ( .A(n9043), .B(n9013), .Y(n9078) );
  NAND2XL U3281 ( .A(n7291), .B(n7261), .Y(n7326) );
  NAND2XL U3282 ( .A(n8167), .B(n8137), .Y(n8202) );
  NAND2XL U3283 ( .A(n11087), .B(n11057), .Y(n11122) );
  NAND2XL U3284 ( .A(n10211), .B(n10181), .Y(n10246) );
  NAND2XL U3285 ( .A(n9335), .B(n9305), .Y(n9370) );
  NAND2XL U3286 ( .A(n8459), .B(n8429), .Y(n8494) );
  NAND2XL U3287 ( .A(n7583), .B(n7553), .Y(n7618) );
  NAND2XL U3288 ( .A(n11379), .B(n11349), .Y(n11414) );
  NAND2XL U3289 ( .A(n10503), .B(n10473), .Y(n10538) );
  NAND2XL U3290 ( .A(n9627), .B(n9597), .Y(n9662) );
  NAND2XL U3291 ( .A(n8751), .B(n8721), .Y(n8786) );
  NAND2XL U3292 ( .A(n7875), .B(n7845), .Y(n7910) );
  NOR4BBXL U3293 ( .AN(n9208), .BN(n9085), .C(n9209), .D(n9159), .Y(n9207) );
  NOR4BBXL U3294 ( .AN(n11544), .BN(n11421), .C(n11545), .D(n11495), .Y(n11543) );
  NOR4BBXL U3295 ( .AN(n8040), .BN(n7917), .C(n8041), .D(n7991), .Y(n8039) );
  NOR4BBXL U3296 ( .AN(n8624), .BN(n8501), .C(n8625), .D(n8575), .Y(n8623) );
  NOR4BBXL U3297 ( .AN(n9792), .BN(n9669), .C(n9793), .D(n9743), .Y(n9791) );
  NOR4BBXL U3298 ( .AN(n10376), .BN(n10253), .C(n10377), .D(n10327), .Y(n10375) );
  NOR4BBXL U3299 ( .AN(n10960), .BN(n10837), .C(n10961), .D(n10911), .Y(n10959) );
  NOR4BBXL U3300 ( .AN(n10084), .BN(n9961), .C(n10085), .D(n10035), .Y(n10083)
         );
  NOR4BBXL U3301 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n270), .BN(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n146), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n271), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n221), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n269) );
  NOR4BBXL U3302 ( .AN(n11252), .BN(n11129), .C(n11253), .D(n11203), .Y(n11251) );
  NOR4BBXL U3303 ( .AN(n8332), .BN(n8209), .C(n8333), .D(n8283), .Y(n8331) );
  NOR4BBXL U3304 ( .AN(n7456), .BN(n7333), .C(n7457), .D(n7407), .Y(n7455) );
  NOR4BBXL U3305 ( .AN(n9500), .BN(n9377), .C(n9501), .D(n9451), .Y(n9499) );
  NOR4BBXL U3306 ( .AN(n7748), .BN(n7625), .C(n7749), .D(n7699), .Y(n7747) );
  NOR4BBXL U3307 ( .AN(n10668), .BN(n10545), .C(n10669), .D(n10619), .Y(n10667) );
  NOR4BBXL U3308 ( .AN(n8916), .BN(n8793), .C(n8917), .D(n8867), .Y(n8915) );
  AOI211XL U3309 ( .A0(n140), .A1(n3062), .B0(n9210), .C0(n9211), .Y(n9206) );
  OR2XL U3310 ( .A(n9188), .B(n9179), .Y(n9211) );
  AOI211XL U3311 ( .A0(n146), .A1(n2579), .B0(n11546), .C0(n11547), .Y(n11542)
         );
  OR2XL U3312 ( .A(n11524), .B(n11515), .Y(n11547) );
  AOI211XL U3313 ( .A0(n150), .A1(n3303), .B0(n8042), .C0(n8043), .Y(n8038) );
  OR2XL U3314 ( .A(n8020), .B(n8011), .Y(n8043) );
  AOI211XL U3315 ( .A0(n144), .A1(n3181), .B0(n8626), .C0(n8627), .Y(n8622) );
  OR2XL U3316 ( .A(n8604), .B(n8595), .Y(n8627) );
  AOI211XL U3317 ( .A0(n148), .A1(n2943), .B0(n9794), .C0(n9795), .Y(n9790) );
  OR2XL U3318 ( .A(n9772), .B(n9763), .Y(n9795) );
  AOI211XL U3319 ( .A0(n142), .A1(n2822), .B0(n10378), .C0(n10379), .Y(n10374)
         );
  OR2XL U3320 ( .A(n10356), .B(n10347), .Y(n10379) );
  AOI211XL U3321 ( .A0(n139), .A1(n2701), .B0(n10962), .C0(n10963), .Y(n10958)
         );
  OR2XL U3322 ( .A(n10940), .B(n10931), .Y(n10963) );
  AOI211XL U3323 ( .A0(n135), .A1(n2882), .B0(n10086), .C0(n10087), .Y(n10082)
         );
  OR2XL U3324 ( .A(n10064), .B(n10055), .Y(n10087) );
  AOI211XL U3325 ( .A0(n136), .A1(n3483), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n272), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n273), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n268) );
  OR2XL U3326 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n250), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n241), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n273) );
  AOI211XL U3327 ( .A0(n137), .A1(n2640), .B0(n11254), .C0(n11255), .Y(n11250)
         );
  OR2XL U3328 ( .A(n11232), .B(n11223), .Y(n11255) );
  AOI211XL U3329 ( .A0(n138), .A1(n3242), .B0(n8334), .C0(n8335), .Y(n8330) );
  OR2XL U3330 ( .A(n8312), .B(n8303), .Y(n8335) );
  AOI211XL U3331 ( .A0(n141), .A1(n3422), .B0(n7458), .C0(n7459), .Y(n7454) );
  OR2XL U3332 ( .A(n7436), .B(n7427), .Y(n7459) );
  AOI211XL U3333 ( .A0(n143), .A1(n3004), .B0(n9502), .C0(n9503), .Y(n9498) );
  OR2XL U3334 ( .A(n9480), .B(n9471), .Y(n9503) );
  AOI211XL U3335 ( .A0(n145), .A1(n3364), .B0(n7750), .C0(n7751), .Y(n7746) );
  OR2XL U3336 ( .A(n7728), .B(n7719), .Y(n7751) );
  AOI211XL U3337 ( .A0(n147), .A1(n2761), .B0(n10670), .C0(n10671), .Y(n10666)
         );
  OR2XL U3338 ( .A(n10648), .B(n10639), .Y(n10671) );
  AOI211XL U3339 ( .A0(n149), .A1(n3123), .B0(n8918), .C0(n8919), .Y(n8914) );
  OR2XL U3340 ( .A(n8896), .B(n8887), .Y(n8919) );
  AOI211XL U3341 ( .A0(n135), .A1(n2882), .B0(n10105), .C0(n10106), .Y(n10102)
         );
  AOI211XL U3342 ( .A0(n136), .A1(n3483), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n291), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n292), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n288) );
  AOI211XL U3343 ( .A0(n138), .A1(n3242), .B0(n8353), .C0(n8354), .Y(n8350) );
  AOI211XL U3344 ( .A0(n137), .A1(n2640), .B0(n11273), .C0(n11274), .Y(n11270)
         );
  AOI211XL U3345 ( .A0(n139), .A1(n2701), .B0(n10981), .C0(n10982), .Y(n10978)
         );
  AOI211XL U3346 ( .A0(n141), .A1(n3422), .B0(n7477), .C0(n7478), .Y(n7474) );
  AOI211XL U3347 ( .A0(n140), .A1(n3062), .B0(n9229), .C0(n9230), .Y(n9226) );
  AOI211XL U3348 ( .A0(n142), .A1(n2822), .B0(n10397), .C0(n10398), .Y(n10394)
         );
  AOI211XL U3349 ( .A0(n143), .A1(n3004), .B0(n9521), .C0(n9522), .Y(n9518) );
  AOI211XL U3350 ( .A0(n144), .A1(n3181), .B0(n8645), .C0(n8646), .Y(n8642) );
  AOI211XL U3351 ( .A0(n145), .A1(n3364), .B0(n7769), .C0(n7770), .Y(n7766) );
  AOI211XL U3352 ( .A0(n146), .A1(n2579), .B0(n11565), .C0(n11566), .Y(n11562)
         );
  AOI211XL U3353 ( .A0(n147), .A1(n2761), .B0(n10689), .C0(n10690), .Y(n10686)
         );
  AOI211XL U3354 ( .A0(n148), .A1(n2943), .B0(n9813), .C0(n9814), .Y(n9810) );
  AOI211XL U3355 ( .A0(n149), .A1(n3123), .B0(n8937), .C0(n8938), .Y(n8934) );
  AOI211XL U3356 ( .A0(n150), .A1(n3303), .B0(n8061), .C0(n8062), .Y(n8058) );
  NAND4XL U3357 ( .A(n9949), .B(n9956), .C(n9957), .D(n9958), .Y(n9951) );
  NAND4XL U3358 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n134), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n141), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n142), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n143), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n136) );
  NAND4XL U3359 ( .A(n11117), .B(n11124), .C(n11125), .D(n11126), .Y(n11119)
         );
  NAND4XL U3360 ( .A(n8197), .B(n8204), .C(n8205), .D(n8206), .Y(n8199) );
  NAND4XL U3361 ( .A(n10825), .B(n10832), .C(n10833), .D(n10834), .Y(n10827)
         );
  NAND4XL U3362 ( .A(n9073), .B(n9080), .C(n9081), .D(n9082), .Y(n9075) );
  NAND4XL U3363 ( .A(n7321), .B(n7328), .C(n7329), .D(n7330), .Y(n7323) );
  NAND4XL U3364 ( .A(n10241), .B(n10248), .C(n10249), .D(n10250), .Y(n10243)
         );
  NAND4XL U3365 ( .A(n9365), .B(n9372), .C(n9373), .D(n9374), .Y(n9367) );
  NAND4XL U3366 ( .A(n8489), .B(n8496), .C(n8497), .D(n8498), .Y(n8491) );
  NAND4XL U3367 ( .A(n7613), .B(n7620), .C(n7621), .D(n7622), .Y(n7615) );
  NAND4XL U3368 ( .A(n11409), .B(n11416), .C(n11417), .D(n11418), .Y(n11411)
         );
  NAND4XL U3369 ( .A(n10533), .B(n10540), .C(n10541), .D(n10542), .Y(n10535)
         );
  NAND4XL U3370 ( .A(n9657), .B(n9664), .C(n9665), .D(n9666), .Y(n9659) );
  NAND4XL U3371 ( .A(n8781), .B(n8788), .C(n8789), .D(n8790), .Y(n8783) );
  NAND4XL U3372 ( .A(n7905), .B(n7912), .C(n7913), .D(n7914), .Y(n7907) );
  NAND4XL U3373 ( .A(n9961), .B(n9958), .C(n9962), .D(n9963), .Y(n9936) );
  NAND4XL U3374 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n146), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n143), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n147), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n148), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n121) );
  NAND4XL U3375 ( .A(n11129), .B(n11126), .C(n11130), .D(n11131), .Y(n11104)
         );
  NAND4XL U3376 ( .A(n8209), .B(n8206), .C(n8210), .D(n8211), .Y(n8184) );
  NAND4XL U3377 ( .A(n10837), .B(n10834), .C(n10838), .D(n10839), .Y(n10812)
         );
  NAND4XL U3378 ( .A(n9085), .B(n9082), .C(n9086), .D(n9087), .Y(n9060) );
  NAND4XL U3379 ( .A(n7333), .B(n7330), .C(n7334), .D(n7335), .Y(n7308) );
  NAND4XL U3380 ( .A(n10253), .B(n10250), .C(n10254), .D(n10255), .Y(n10228)
         );
  NAND4XL U3381 ( .A(n9377), .B(n9374), .C(n9378), .D(n9379), .Y(n9352) );
  NAND4XL U3382 ( .A(n8501), .B(n8498), .C(n8502), .D(n8503), .Y(n8476) );
  NAND4XL U3383 ( .A(n7625), .B(n7622), .C(n7626), .D(n7627), .Y(n7600) );
  NAND4XL U3384 ( .A(n11421), .B(n11418), .C(n11422), .D(n11423), .Y(n11396)
         );
  NAND4XL U3385 ( .A(n10545), .B(n10542), .C(n10546), .D(n10547), .Y(n10520)
         );
  NAND4XL U3386 ( .A(n9669), .B(n9666), .C(n9670), .D(n9671), .Y(n9644) );
  NAND4XL U3387 ( .A(n8793), .B(n8790), .C(n8794), .D(n8795), .Y(n8768) );
  NAND4XL U3388 ( .A(n7917), .B(n7914), .C(n7918), .D(n7919), .Y(n7892) );
  NAND4XL U3389 ( .A(n10010), .B(n9904), .C(n10109), .D(n10110), .Y(n10108) );
  NAND4XL U3390 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n196), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n87), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n295), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n296), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n294) );
  NAND4XL U3391 ( .A(n8258), .B(n8152), .C(n8357), .D(n8358), .Y(n8356) );
  NAND4XL U3392 ( .A(n11178), .B(n11072), .C(n11277), .D(n11278), .Y(n11276)
         );
  NAND4XL U3393 ( .A(n10886), .B(n10780), .C(n10985), .D(n10986), .Y(n10984)
         );
  NAND4XL U3394 ( .A(n7382), .B(n7276), .C(n7481), .D(n7482), .Y(n7480) );
  NAND4XL U3395 ( .A(n9134), .B(n9028), .C(n9233), .D(n9234), .Y(n9232) );
  NAND4XL U3396 ( .A(n10302), .B(n10196), .C(n10401), .D(n10402), .Y(n10400)
         );
  NAND4XL U3397 ( .A(n9426), .B(n9320), .C(n9525), .D(n9526), .Y(n9524) );
  NAND4XL U3398 ( .A(n8550), .B(n8444), .C(n8649), .D(n8650), .Y(n8648) );
  NAND4XL U3399 ( .A(n7674), .B(n7568), .C(n7773), .D(n7774), .Y(n7772) );
  NAND4XL U3400 ( .A(n11470), .B(n11364), .C(n11569), .D(n11570), .Y(n11568)
         );
  NAND4XL U3401 ( .A(n10594), .B(n10488), .C(n10693), .D(n10694), .Y(n10692)
         );
  NAND4XL U3402 ( .A(n9718), .B(n9612), .C(n9817), .D(n9818), .Y(n9816) );
  NAND4XL U3403 ( .A(n8842), .B(n8736), .C(n8941), .D(n8942), .Y(n8940) );
  NAND4XL U3404 ( .A(n7966), .B(n7860), .C(n8065), .D(n8066), .Y(n8064) );
  AOI21XL U3405 ( .A0(n6556), .A1(n13228), .B0(n6548), .Y(n13419) );
  AOI21XL U3406 ( .A0(n6851), .A1(n12598), .B0(n6843), .Y(n12789) );
  AOI21XL U3407 ( .A0(n6897), .A1(n12913), .B0(n6889), .Y(n13104) );
  AOI22XL U3408 ( .A0(n6121), .A1(n1142), .B0(n6130), .B1(n1281), .Y(n14103)
         );
  AOI22XL U3409 ( .A0(n5353), .A1(n1003), .B0(n5362), .B1(n1311), .Y(n17253)
         );
  AOI22XL U3410 ( .A0(n4999), .A1(n947), .B0(n5008), .B1(n1323), .Y(n18513) );
  AOI22XL U3411 ( .A0(n5825), .A1(n1087), .B0(n5834), .B1(n1293), .Y(n15363)
         );
  AOI22XL U3412 ( .A0(n5741), .A1(n1073), .B0(n5750), .B1(n1296), .Y(n15678)
         );
  AOI22XL U3413 ( .A0(n4883), .A1(n933), .B0(n4892), .B1(n1326), .Y(n18828) );
  AOI22XL U3414 ( .A0(n5437), .A1(n1017), .B0(n5446), .B1(n1308), .Y(n16938)
         );
  AOI22XL U3415 ( .A0(n5901), .A1(n1101), .B0(n5910), .B1(n1290), .Y(n15048)
         );
  AOI22XL U3416 ( .A0(n5513), .A1(n1031), .B0(n5522), .B1(n1305), .Y(n16623)
         );
  AOI22XL U3417 ( .A0(n5083), .A1(n961), .B0(n5092), .B1(n1320), .Y(n18198) );
  AOI22XL U3418 ( .A0(n5977), .A1(n1115), .B0(n5986), .B1(n1287), .Y(n14733)
         );
  AOI22XL U3419 ( .A0(n5589), .A1(n1045), .B0(n5598), .B1(n1302), .Y(n16308)
         );
  AOI22XL U3420 ( .A0(n5191), .A1(n975), .B0(n5200), .B1(n1317), .Y(n17883) );
  AOI22XL U3421 ( .A0(n6053), .A1(n1129), .B0(n6062), .B1(n1284), .Y(n14418)
         );
  AOI22XL U3422 ( .A0(n5665), .A1(n1059), .B0(n5674), .B1(n1299), .Y(n15993)
         );
  AOI22XL U3423 ( .A0(n5269), .A1(n989), .B0(n5278), .B1(n1314), .Y(n17568) );
  OAI211XL U3424 ( .A0(n2881), .A1(n90), .B0(n10099), .C0(n10154), .Y(n10146)
         );
  OAI211XL U3425 ( .A0(n3482), .A1(n91), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n285), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n340), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n332) );
  OAI211XL U3426 ( .A0(n3241), .A1(n93), .B0(n8347), .C0(n8402), .Y(n8394) );
  OAI211XL U3427 ( .A0(n2639), .A1(n92), .B0(n11267), .C0(n11322), .Y(n11314)
         );
  OAI211XL U3428 ( .A0(n2700), .A1(n94), .B0(n10975), .C0(n11030), .Y(n11022)
         );
  OAI211XL U3429 ( .A0(n3421), .A1(n95), .B0(n7471), .C0(n7526), .Y(n7518) );
  OAI211XL U3430 ( .A0(n3061), .A1(n96), .B0(n9223), .C0(n9278), .Y(n9270) );
  OAI211XL U3431 ( .A0(n2821), .A1(n97), .B0(n10391), .C0(n10446), .Y(n10438)
         );
  OAI211XL U3432 ( .A0(n3003), .A1(n98), .B0(n9515), .C0(n9570), .Y(n9562) );
  OAI211XL U3433 ( .A0(n3180), .A1(n99), .B0(n8639), .C0(n8694), .Y(n8686) );
  OAI211XL U3434 ( .A0(n3363), .A1(n100), .B0(n7763), .C0(n7818), .Y(n7810) );
  OAI211XL U3435 ( .A0(n2578), .A1(n101), .B0(n11559), .C0(n11614), .Y(n11606)
         );
  OAI211XL U3436 ( .A0(n2760), .A1(n102), .B0(n10683), .C0(n10738), .Y(n10730)
         );
  OAI211XL U3437 ( .A0(n2942), .A1(n103), .B0(n9807), .C0(n9862), .Y(n9854) );
  OAI211XL U3438 ( .A0(n3122), .A1(n104), .B0(n8931), .C0(n8986), .Y(n8978) );
  OAI211XL U3439 ( .A0(n3302), .A1(n105), .B0(n8055), .C0(n8110), .Y(n8102) );
  AOI222XL U3440 ( .A0(n759), .A1(n1655), .B0(n1160), .B1(n1178), .C0(n6597), 
        .C1(n13543), .Y(n13600) );
  AOI222XL U3441 ( .A0(n757), .A1(n1742), .B0(n1191), .B1(n1213), .C0(n6844), 
        .C1(n12598), .Y(n12655) );
  AOI222XL U3442 ( .A0(n758), .A1(n1713), .B0(n1200), .B1(n1219), .C0(n6890), 
        .C1(n12913), .Y(n12970) );
  AOI222XL U3443 ( .A0(n756), .A1(n1684), .B0(n1151), .B1(n1173), .C0(n6549), 
        .C1(n13228), .Y(n13285) );
  AND2X1 U3444 ( .A(n18647), .B(n18710), .Y(n654) );
  AND2X1 U3445 ( .A(n15497), .B(n15560), .Y(n653) );
  AND2X1 U3446 ( .A(n14867), .B(n14930), .Y(n656) );
  AND2X1 U3447 ( .A(n18017), .B(n18080), .Y(n658) );
  AND2X1 U3448 ( .A(n14237), .B(n14300), .Y(n662) );
  AND2X1 U3449 ( .A(n16127), .B(n16190), .Y(n660) );
  AND2X1 U3450 ( .A(n17387), .B(n17450), .Y(n664) );
  AND2X1 U3451 ( .A(n13922), .B(n13985), .Y(n649) );
  AND2X1 U3452 ( .A(n17072), .B(n17135), .Y(n650) );
  AND2X1 U3453 ( .A(n18332), .B(n18395), .Y(n651) );
  AND2X1 U3454 ( .A(n15182), .B(n15245), .Y(n652) );
  AND2X1 U3455 ( .A(n16757), .B(n16820), .Y(n655) );
  AND2X1 U3456 ( .A(n16442), .B(n16505), .Y(n657) );
  AND2X1 U3457 ( .A(n14552), .B(n14615), .Y(n659) );
  AND2X1 U3458 ( .A(n17702), .B(n17765), .Y(n661) );
  AND2X1 U3459 ( .A(n15812), .B(n15875), .Y(n663) );
  AOI222XL U3460 ( .A0(n1072), .A1(n5768), .B0(n15442), .B1(n15444), .C0(
        n15472), .C1(n5741), .Y(n15469) );
  AOI222XL U3461 ( .A0(n960), .A1(n5110), .B0(n17962), .B1(n17964), .C0(n17992), .C1(n5083), .Y(n17989) );
  AOI222XL U3462 ( .A0(n1128), .A1(n6080), .B0(n14182), .B1(n14184), .C0(
        n14212), .C1(n6053), .Y(n14209) );
  AOI222XL U3463 ( .A0(n932), .A1(n4910), .B0(n18592), .B1(n18594), .C0(n18622), .C1(n4883), .Y(n18619) );
  AOI222XL U3464 ( .A0(n1100), .A1(n5928), .B0(n14812), .B1(n14814), .C0(
        n14842), .C1(n5901), .Y(n14839) );
  AOI222XL U3465 ( .A0(n1044), .A1(n5616), .B0(n16072), .B1(n16074), .C0(
        n16102), .C1(n5589), .Y(n16099) );
  AOI222XL U3466 ( .A0(n988), .A1(n5296), .B0(n17332), .B1(n17334), .C0(n17362), .C1(n5269), .Y(n17359) );
  AOI222XL U3467 ( .A0(n1141), .A1(n6151), .B0(n13867), .B1(n13869), .C0(
        n13897), .C1(n6121), .Y(n13894) );
  AOI222XL U3468 ( .A0(n1002), .A1(n5380), .B0(n17017), .B1(n17019), .C0(
        n17047), .C1(n5353), .Y(n17044) );
  AOI222XL U3469 ( .A0(n946), .A1(n5026), .B0(n18277), .B1(n18279), .C0(n18307), .C1(n4999), .Y(n18304) );
  AOI222XL U3470 ( .A0(n1086), .A1(n5852), .B0(n15127), .B1(n15129), .C0(
        n15157), .C1(n5825), .Y(n15154) );
  AOI222XL U3471 ( .A0(n1016), .A1(n5464), .B0(n16702), .B1(n16704), .C0(
        n16732), .C1(n5437), .Y(n16729) );
  AOI222XL U3472 ( .A0(n1030), .A1(n5540), .B0(n16387), .B1(n16389), .C0(
        n16417), .C1(n5513), .Y(n16414) );
  AOI222XL U3473 ( .A0(n1114), .A1(n6004), .B0(n14497), .B1(n14499), .C0(
        n14527), .C1(n5977), .Y(n14524) );
  AOI222XL U3474 ( .A0(n974), .A1(n5218), .B0(n17647), .B1(n17649), .C0(n17677), .C1(n5191), .Y(n17674) );
  AOI222XL U3475 ( .A0(n1058), .A1(n5692), .B0(n15757), .B1(n15759), .C0(
        n15787), .C1(n5665), .Y(n15784) );
  OAI211XL U3476 ( .A0(n12663), .A1(n1267), .B0(n12667), .C0(n12750), .Y(
        n12749) );
  OAI211XL U3477 ( .A0(n12978), .A1(n1270), .B0(n12982), .C0(n13065), .Y(
        n13064) );
  OAI211XL U3478 ( .A0(n13293), .A1(n1273), .B0(n13297), .C0(n13380), .Y(
        n13379) );
  NOR2X4 U3479 ( .A(n4140), .B(n4142), .Y(n302) );
  NOR2X2 U3480 ( .A(n4143), .B(n4138), .Y(n303) );
  AOI211XL U3481 ( .A0(n6919), .A1(n11691), .B0(n11741), .C0(n11878), .Y(
        n11877) );
  AOI211XL U3482 ( .A0(n6873), .A1(top_core_KE_sb1_n116), .B0(
        top_core_KE_sb1_n168), .C0(top_core_KE_sb1_n307), .Y(
        top_core_KE_sb1_n306) );
  AOI211XL U3483 ( .A0(n6626), .A1(n12322), .B0(n12372), .C0(n12509), .Y(
        n12508) );
  AOI211XL U3484 ( .A0(n6579), .A1(n12007), .B0(n12057), .C0(n12194), .Y(
        n12193) );
  AOI211XL U3485 ( .A0(n6602), .A1(n13583), .B0(n13633), .C0(n13769), .Y(
        n13768) );
  NOR2XL U3486 ( .A(n13538), .B(n1647), .Y(n13595) );
  AOI222XL U3487 ( .A0(n1172), .A1(n6633), .B0(n13395), .B1(n1693), .C0(n6544), 
        .C1(n13268), .Y(n13424) );
  AOI21XL U3488 ( .A0(n6598), .A1(n1277), .B0(n6586), .Y(n13704) );
  AOI31XL U3489 ( .A0(n1172), .A1(n1150), .A2(n13425), .B0(n263), .Y(n13429)
         );
  AOI31XL U3490 ( .A0(n1212), .A1(n1190), .A2(n12795), .B0(n262), .Y(n12799)
         );
  AOI31XL U3491 ( .A0(n1180), .A1(n1159), .A2(n13740), .B0(n261), .Y(n13744)
         );
  AOI31XL U3492 ( .A0(n1218), .A1(n1199), .A2(n13110), .B0(n260), .Y(n13114)
         );
  AOI31XL U3493 ( .A0(n1215), .A1(n1195), .A2(top_core_KE_sb1_n278), .B0(n242), 
        .Y(top_core_KE_sb1_n282) );
  AOI31XL U3494 ( .A0(n1183), .A1(n1164), .A2(n12480), .B0(n241), .Y(n12484)
         );
  AOI31XL U3495 ( .A0(n1221), .A1(n1204), .A2(n11849), .B0(n243), .Y(n11853)
         );
  AOI31XL U3496 ( .A0(n1175), .A1(n1155), .A2(n12165), .B0(n240), .Y(n12169)
         );
  AOI21XL U3497 ( .A0(n6915), .A1(n1258), .B0(n6903), .Y(n11813) );
  AOI21XL U3498 ( .A0(n6869), .A1(n1330), .B0(n6857), .Y(top_core_KE_sb1_n241)
         );
  AOI21XL U3499 ( .A0(n6575), .A1(n1261), .B0(n6563), .Y(n12129) );
  AOI211XL U3500 ( .A0(n6849), .A1(n12598), .B0(n12660), .C0(n12661), .Y(
        n12657) );
  AOI211XL U3501 ( .A0(n6895), .A1(n12913), .B0(n12975), .C0(n12976), .Y(
        n12972) );
  AOI211XL U3502 ( .A0(n6554), .A1(n13228), .B0(n13290), .C0(n13291), .Y(
        n13287) );
  AOI21XL U3503 ( .A0(n6622), .A1(n1265), .B0(n6610), .Y(n12444) );
  AOI211XL U3504 ( .A0(n6849), .A1(n12638), .B0(n12688), .C0(n12824), .Y(
        n12823) );
  AOI211XL U3505 ( .A0(n6895), .A1(n12953), .B0(n13003), .C0(n13139), .Y(
        n13138) );
  AOI211XL U3506 ( .A0(n6554), .A1(n13268), .B0(n13318), .C0(n13454), .Y(
        n13453) );
  AOI222XL U3507 ( .A0(n1221), .A1(n6920), .B0(n11661), .B1(n11663), .C0(
        n11691), .C1(n6904), .Y(n11688) );
  AOI222XL U3508 ( .A0(n1215), .A1(n6874), .B0(top_core_KE_sb1_n86), .B1(
        top_core_KE_sb1_n88), .C0(top_core_KE_sb1_n116), .C1(n6858), .Y(
        top_core_KE_sb1_n113) );
  AOI222XL U3509 ( .A0(n1175), .A1(n6580), .B0(n11977), .B1(n11979), .C0(
        n12007), .C1(n6564), .Y(n12004) );
  AOI222XL U3510 ( .A0(n1183), .A1(n6627), .B0(n1263), .B1(n12294), .C0(n12322), .C1(n6611), .Y(n12319) );
  AOI21XL U3511 ( .A0(n11646), .A1(n6919), .B0(n11702), .Y(n11937) );
  AOI21XL U3512 ( .A0(top_core_KE_sb1_n71), .A1(n6873), .B0(
        top_core_KE_sb1_n127), .Y(top_core_KE_sb1_n366) );
  AOI21XL U3513 ( .A0(n12278), .A1(n6626), .B0(n12333), .Y(n12568) );
  AOI21XL U3514 ( .A0(n11962), .A1(n6579), .B0(n12018), .Y(n12253) );
  AOI211XL U3515 ( .A0(n6919), .A1(n11651), .B0(n11713), .C0(n11714), .Y(
        n11710) );
  AOI211XL U3516 ( .A0(n6873), .A1(top_core_KE_sb1_n76), .B0(
        top_core_KE_sb1_n139), .C0(top_core_KE_sb1_n140), .Y(
        top_core_KE_sb1_n136) );
  AOI211XL U3517 ( .A0(n6579), .A1(n11967), .B0(n12029), .C0(n12030), .Y(
        n12026) );
  AOI211XL U3518 ( .A0(n6626), .A1(n12283), .B0(n12344), .C0(n12345), .Y(
        n12341) );
  AOI211XL U3519 ( .A0(n6602), .A1(n13543), .B0(n13605), .C0(n13606), .Y(
        n13602) );
  AOI222XL U3520 ( .A0(n1162), .A1(n12278), .B0(n12442), .B1(n1761), .C0(n6616), .C1(n667), .Y(n12441) );
  AOI222XL U3521 ( .A0(n1202), .A1(n11646), .B0(n11811), .B1(n1803), .C0(n6909), .C1(n665), .Y(n11810) );
  AOI222XL U3522 ( .A0(n1193), .A1(top_core_KE_sb1_n71), .B0(
        top_core_KE_sb1_n239), .B1(n1824), .C0(n6863), .C1(n666), .Y(
        top_core_KE_sb1_n238) );
  AOI222XL U3523 ( .A0(n1153), .A1(n11962), .B0(n12127), .B1(n1782), .C0(n6569), .C1(n668), .Y(n12126) );
  OAI211XL U3524 ( .A0(n4), .A1(n12608), .B0(n12719), .C0(n12726), .Y(n12723)
         );
  AOI22XL U3525 ( .A0(n1192), .A1(n12608), .B0(n1189), .B1(n1738), .Y(n12726)
         );
  OAI211XL U3526 ( .A0(n5), .A1(n12923), .B0(n13034), .C0(n13041), .Y(n13038)
         );
  AOI22XL U3527 ( .A0(n1201), .A1(n12923), .B0(n1198), .B1(n1709), .Y(n13041)
         );
  AOI22XL U3528 ( .A0(n1205), .A1(n11661), .B0(n1203), .B1(n1802), .Y(n11780)
         );
  AOI22XL U3529 ( .A0(n1196), .A1(top_core_KE_sb1_n86), .B0(n1194), .B1(n1823), 
        .Y(top_core_KE_sb1_n208) );
  AOI22XL U3530 ( .A0(n1156), .A1(n11977), .B0(n1154), .B1(n1781), .Y(n12096)
         );
  AOI22XL U3531 ( .A0(n1165), .A1(n1263), .B0(n1163), .B1(n1760), .Y(n12411)
         );
  OAI211XL U3532 ( .A0(n6), .A1(n1276), .B0(n13664), .C0(n13671), .Y(n13668)
         );
  AOI22XL U3533 ( .A0(n1161), .A1(n13553), .B0(n1158), .B1(n1651), .Y(n13671)
         );
  AOI21XL U3534 ( .A0(n13223), .A1(n6554), .B0(n13279), .Y(n13513) );
  OAI211XL U3535 ( .A0(n17093), .A1(n106), .B0(n17094), .C0(n17095), .Y(n17078) );
  OAI211XL U3536 ( .A0(n13943), .A1(n107), .B0(n13944), .C0(n13945), .Y(n13928) );
  OAI211XL U3537 ( .A0(n18353), .A1(n108), .B0(n18354), .C0(n18355), .Y(n18338) );
  OAI211XL U3538 ( .A0(n15203), .A1(n109), .B0(n15204), .C0(n15205), .Y(n15188) );
  OAI211XL U3539 ( .A0(n15518), .A1(n110), .B0(n15519), .C0(n15520), .Y(n15503) );
  OAI211XL U3540 ( .A0(n18668), .A1(n111), .B0(n18669), .C0(n18670), .Y(n18653) );
  OAI211XL U3541 ( .A0(n16778), .A1(n112), .B0(n16779), .C0(n16780), .Y(n16763) );
  OAI211XL U3542 ( .A0(n14888), .A1(n113), .B0(n14889), .C0(n14890), .Y(n14873) );
  OAI211XL U3543 ( .A0(n16463), .A1(n114), .B0(n16464), .C0(n16465), .Y(n16448) );
  OAI211XL U3544 ( .A0(n18038), .A1(n115), .B0(n18039), .C0(n18040), .Y(n18023) );
  OAI211XL U3545 ( .A0(n14573), .A1(n116), .B0(n14574), .C0(n14575), .Y(n14558) );
  OAI211XL U3546 ( .A0(n16148), .A1(n117), .B0(n16149), .C0(n16150), .Y(n16133) );
  OAI211XL U3547 ( .A0(n17723), .A1(n118), .B0(n17724), .C0(n17725), .Y(n17708) );
  OAI211XL U3548 ( .A0(n14258), .A1(n119), .B0(n14259), .C0(n14260), .Y(n14243) );
  OAI211XL U3549 ( .A0(n15833), .A1(n120), .B0(n15834), .C0(n15835), .Y(n15818) );
  OAI211XL U3550 ( .A0(n17408), .A1(n121), .B0(n17409), .C0(n17410), .Y(n17393) );
  AOI222XL U3551 ( .A0(n11717), .A1(n753), .B0(n1202), .B1(n1223), .C0(n1205), 
        .C1(n1258), .Y(n11830) );
  AOI222XL U3552 ( .A0(top_core_KE_sb1_n144), .A1(n754), .B0(n1193), .B1(n1217), .C0(n1196), .C1(n1330), .Y(top_core_KE_sb1_n259) );
  AOI222XL U3553 ( .A0(n12033), .A1(n755), .B0(n1153), .B1(n1177), .C0(n1156), 
        .C1(n1261), .Y(n12146) );
  AOI222XL U3554 ( .A0(n12348), .A1(n752), .B0(n1162), .B1(n1182), .C0(n1165), 
        .C1(n1265), .Y(n12461) );
  NAND3XL U3555 ( .A(n1274), .B(n1150), .C(n13425), .Y(n13427) );
  AOI222XL U3556 ( .A0(n6839), .A1(n1268), .B0(n12648), .B1(n678), .C0(n6851), 
        .C1(n1212), .Y(n12735) );
  AOI222XL U3557 ( .A0(n6592), .A1(n1277), .B0(n13593), .B1(n679), .C0(n6604), 
        .C1(n1180), .Y(n13680) );
  AOI222XL U3558 ( .A0(n6885), .A1(n1271), .B0(n12963), .B1(n680), .C0(n6897), 
        .C1(n1218), .Y(n13050) );
  AOI222XL U3559 ( .A0(n6544), .A1(n1274), .B0(n13278), .B1(n692), .C0(n6556), 
        .C1(n1172), .Y(n13365) );
  NAND3XL U3560 ( .A(top_core_KE_prev_key1_reg_90_), .B(n1278), .C(n720), .Y(
        n13700) );
  OAI2BB1XL U3561 ( .A0N(n1688), .A1N(n13395), .B0(n180), .Y(n13394) );
  OAI2BB1XL U3562 ( .A0N(n1746), .A1N(n12765), .B0(n181), .Y(n12764) );
  OAI2BB1XL U3563 ( .A0N(n1659), .A1N(n13710), .B0(n183), .Y(n13709) );
  OAI2BB1XL U3564 ( .A0N(n1717), .A1N(n13080), .B0(n182), .Y(n13079) );
  AOI222XL U3565 ( .A0(top_core_KE_prev_key1_reg_29_), .A1(n12553), .B0(n6527), 
        .B1(n1265), .C0(n6528), .C1(n12322), .Y(n12552) );
  AOI222XL U3566 ( .A0(n1639), .A1(n13813), .B0(n6516), .B1(n1277), .C0(n6517), 
        .C1(n13583), .Y(n13812) );
  AOI222XL U3567 ( .A0(n1797), .A1(n11922), .B0(n6823), .B1(n1258), .C0(n6824), 
        .C1(n11691), .Y(n11921) );
  AOI222XL U3568 ( .A0(n1818), .A1(top_core_KE_sb1_n351), .B0(n6799), .B1(
        n1330), .C0(n6802), .C1(top_core_KE_sb1_n116), .Y(top_core_KE_sb1_n350) );
  AOI222XL U3569 ( .A0(n1776), .A1(n12238), .B0(n6502), .B1(n1261), .C0(n6505), 
        .C1(n12007), .Y(n12237) );
  AOI21XL U3570 ( .A0(n6604), .A1(n13543), .B0(n6596), .Y(n13734) );
  AOI21XL U3571 ( .A0(n6920), .A1(n11651), .B0(n6913), .Y(n11843) );
  AOI21XL U3572 ( .A0(n6874), .A1(top_core_KE_sb1_n76), .B0(n6867), .Y(
        top_core_KE_sb1_n272) );
  AOI21XL U3573 ( .A0(n6580), .A1(n11967), .B0(n6573), .Y(n12159) );
  AOI21XL U3574 ( .A0(n6627), .A1(n12283), .B0(n6620), .Y(n12474) );
  AOI222XL U3575 ( .A0(n6604), .A1(n1653), .B0(n13596), .B1(n13597), .C0(n6602), .C1(n1652), .Y(n13590) );
  AOI222XL U3576 ( .A0(n1215), .A1(n6933), .B0(top_core_KE_sb1_n247), .B1(
        n1836), .C0(n6863), .C1(top_core_KE_sb1_n116), .Y(top_core_KE_sb1_n277) );
  AOI222XL U3577 ( .A0(n1183), .A1(n6658), .B0(n12450), .B1(n1771), .C0(n6616), 
        .C1(n12322), .Y(n12479) );
  AOI222XL U3578 ( .A0(n1221), .A1(n6948), .B0(n11819), .B1(n1815), .C0(n6909), 
        .C1(n11691), .Y(n11848) );
  AOI222XL U3579 ( .A0(n1175), .A1(n6642), .B0(n12135), .B1(n1794), .C0(n6569), 
        .C1(n12007), .Y(n12164) );
  AOI222XL U3580 ( .A0(n1212), .A1(n6925), .B0(n12765), .B1(n1751), .C0(n6839), 
        .C1(n12638), .Y(n12794) );
  AOI222XL U3581 ( .A0(n1180), .A1(n6650), .B0(n13710), .B1(n1661), .C0(n6592), 
        .C1(n13583), .Y(n13739) );
  AOI222XL U3582 ( .A0(n1218), .A1(n6940), .B0(n13080), .B1(n1722), .C0(n6885), 
        .C1(n12953), .Y(n13109) );
  NAND4XL U3583 ( .A(n13333), .B(n13246), .C(n13482), .D(n13483), .Y(n13481)
         );
  AOI32XL U3584 ( .A0(n1677), .A1(n1150), .A2(n1688), .B0(n13387), .B1(n1273), 
        .Y(n13482) );
  NAND4XL U3585 ( .A(n12703), .B(n12616), .C(n12852), .D(n12853), .Y(n12851)
         );
  AOI32XL U3586 ( .A0(n1736), .A1(n1190), .A2(n1746), .B0(n12757), .B1(n1267), 
        .Y(n12852) );
  NAND4XL U3587 ( .A(n13018), .B(n12931), .C(n13167), .D(n13168), .Y(n13166)
         );
  AOI32XL U3588 ( .A0(n1707), .A1(n1199), .A2(n1717), .B0(n13072), .B1(n1270), 
        .Y(n13167) );
  NAND4XL U3589 ( .A(n13648), .B(n13561), .C(n13797), .D(n13798), .Y(n13796)
         );
  AOI32XL U3590 ( .A0(n1644), .A1(n1159), .A2(n1659), .B0(n13702), .B1(n1276), 
        .Y(n13797) );
  AOI222XL U3591 ( .A0(n6920), .A1(n1807), .B0(n11704), .B1(n11705), .C0(n6919), .C1(n1803), .Y(n11698) );
  AOI222XL U3592 ( .A0(n6874), .A1(n1828), .B0(top_core_KE_sb1_n129), .B1(
        top_core_KE_sb1_n130), .C0(n6873), .C1(n1824), .Y(top_core_KE_sb1_n123) );
  AOI222XL U3593 ( .A0(n6580), .A1(n1786), .B0(n12020), .B1(n12021), .C0(n6579), .C1(n1782), .Y(n12014) );
  AOI222XL U3594 ( .A0(n6627), .A1(n1763), .B0(n12335), .B1(n12336), .C0(n6626), .C1(n1761), .Y(n12329) );
  AOI222XL U3595 ( .A0(n6851), .A1(n1742), .B0(n12651), .B1(n12652), .C0(n6849), .C1(n1739), .Y(n12645) );
  AOI222XL U3596 ( .A0(n6897), .A1(n1713), .B0(n12966), .B1(n12967), .C0(n6895), .C1(n1710), .Y(n12960) );
  AOI222XL U3597 ( .A0(n6556), .A1(n1684), .B0(n13281), .B1(n13282), .C0(n6554), .C1(n1681), .Y(n13275) );
  AOI222XL U3598 ( .A0(n761), .A1(n1807), .B0(n745), .B1(n1222), .C0(n6914), 
        .C1(n11651), .Y(n11708) );
  AOI222XL U3599 ( .A0(n762), .A1(n1828), .B0(n746), .B1(n1216), .C0(n6868), 
        .C1(top_core_KE_sb1_n76), .Y(top_core_KE_sb1_n133) );
  AOI222XL U3600 ( .A0(n760), .A1(n1765), .B0(n744), .B1(n1181), .C0(n6621), 
        .C1(n12283), .Y(n12339) );
  AOI222XL U3601 ( .A0(n763), .A1(n1786), .B0(n747), .B1(n1176), .C0(n6574), 
        .C1(n11967), .Y(n12024) );
  AOI222XL U3602 ( .A0(n1148), .A1(n13223), .B0(n13387), .B1(n1681), .C0(n6544), .C1(n670), .Y(n13386) );
  NAND3XL U3603 ( .A(n1674), .B(n13282), .C(n717), .Y(n13385) );
  AOI32XL U3604 ( .A0(n1211), .A1(n1204), .A2(n1810), .B0(n11811), .B1(n1257), 
        .Y(n11906) );
  AOI32XL U3605 ( .A0(n1210), .A1(n1195), .A2(n1831), .B0(top_core_KE_sb1_n239), .B1(n1329), .Y(top_core_KE_sb1_n335) );
  AOI32XL U3606 ( .A0(n1171), .A1(n1164), .A2(n1768), .B0(n12442), .B1(n1263), 
        .Y(n12537) );
  AOI32XL U3607 ( .A0(n1170), .A1(n1155), .A2(n1789), .B0(n12127), .B1(n1260), 
        .Y(n12222) );
  AOI211XL U3608 ( .A0(n6616), .A1(n1266), .B0(n12391), .C0(n12392), .Y(n12390) );
  AOI211XL U3609 ( .A0(n6839), .A1(n1269), .B0(n12707), .C0(n12708), .Y(n12706) );
  AOI211XL U3610 ( .A0(n6592), .A1(n1278), .B0(n13652), .C0(n13653), .Y(n13651) );
  AOI211XL U3611 ( .A0(n6885), .A1(n1272), .B0(n13022), .C0(n13023), .Y(n13021) );
  AOI211XL U3612 ( .A0(n6544), .A1(n1275), .B0(n13337), .C0(n13338), .Y(n13336) );
  AND2X1 U3613 ( .A(n189), .B(n12725), .Y(n719) );
  AND2X1 U3614 ( .A(n191), .B(n13040), .Y(n721) );
  AND2X1 U3615 ( .A(n187), .B(n13355), .Y(n717) );
  AND2X1 U3616 ( .A(n190), .B(n13670), .Y(n720) );
  AND2X1 U3617 ( .A(n185), .B(n11778), .Y(n714) );
  AND2X1 U3618 ( .A(n186), .B(top_core_KE_sb1_n206), .Y(n715) );
  AND2X1 U3619 ( .A(n46), .B(n12409), .Y(n716) );
  AND2X1 U3620 ( .A(n188), .B(n12094), .Y(n718) );
  OAI211XL U3621 ( .A0(n13608), .A1(n13553), .B0(n13612), .C0(n13695), .Y(
        n13694) );
  AOI22XL U3622 ( .A0(n11661), .A1(n1344), .B0(n1211), .B1(n11691), .Y(n11662)
         );
  AOI22XL U3623 ( .A0(top_core_KE_sb1_n86), .A1(n1345), .B0(n1210), .B1(
        top_core_KE_sb1_n116), .Y(top_core_KE_sb1_n87) );
  AOI22XL U3624 ( .A0(n1264), .A1(n1358), .B0(n1171), .B1(n12322), .Y(n12293)
         );
  AOI22XL U3625 ( .A0(n11977), .A1(n1359), .B0(n1170), .B1(n12007), .Y(n11978)
         );
  AOI22XL U3626 ( .A0(n13553), .A1(n1647), .B0(n1643), .B1(n13583), .Y(n13554)
         );
  NOR2XL U3627 ( .A(n12278), .B(n1358), .Y(n12334) );
  NOR2XL U3628 ( .A(n11646), .B(n1344), .Y(n11703) );
  NOR2XL U3629 ( .A(top_core_KE_sb1_n71), .B(n1345), .Y(top_core_KE_sb1_n128)
         );
  NOR2XL U3630 ( .A(n11962), .B(n1359), .Y(n12019) );
  OAI31XL U3631 ( .A0(n11691), .A1(n1350), .A2(n1344), .B0(n11715), .Y(n11714)
         );
  OAI31XL U3632 ( .A0(top_core_KE_sb1_n116), .A1(n1352), .A2(n1345), .B0(
        top_core_KE_sb1_n141), .Y(top_core_KE_sb1_n140) );
  OAI31XL U3633 ( .A0(n12322), .A1(n1364), .A2(n1358), .B0(n12346), .Y(n12345)
         );
  OAI31XL U3634 ( .A0(n12007), .A1(n1366), .A2(n1359), .B0(n12031), .Y(n12030)
         );
  OAI31XL U3635 ( .A0(n13583), .A1(n1365), .A2(n1645), .B0(n13607), .Y(n13606)
         );
  OAI31XL U3636 ( .A0(n13268), .A1(n1367), .A2(n1674), .B0(n13292), .Y(n13291)
         );
  OAI31XL U3637 ( .A0(n12638), .A1(n1353), .A2(n1732), .B0(n12662), .Y(n12661)
         );
  OAI31XL U3638 ( .A0(n12953), .A1(n1351), .A2(n1703), .B0(n12977), .Y(n12976)
         );
  AOI31XL U3639 ( .A0(n1350), .A1(n11691), .A2(n6830), .B0(n11781), .Y(n11774)
         );
  AOI31XL U3640 ( .A0(n1352), .A1(top_core_KE_sb1_n116), .A2(n6809), .B0(
        top_core_KE_sb1_n209), .Y(top_core_KE_sb1_n202) );
  AOI31XL U3641 ( .A0(n1364), .A1(n12322), .A2(n6534), .B0(n12412), .Y(n12405)
         );
  AOI31XL U3642 ( .A0(n1366), .A1(n12007), .A2(n6512), .B0(n12097), .Y(n12090)
         );
  AOI31XL U3643 ( .A0(n1365), .A1(n13583), .A2(n6523), .B0(n13672), .Y(n13666)
         );
  AOI31XL U3644 ( .A0(n1353), .A1(n12638), .A2(n6780), .B0(n12727), .Y(n12721)
         );
  AOI31XL U3645 ( .A0(n1351), .A1(n12953), .A2(n6819), .B0(n13042), .Y(n13036)
         );
  AOI31XL U3646 ( .A0(n1367), .A1(n13268), .A2(n6477), .B0(n13357), .Y(n13351)
         );
  AOI22XL U3647 ( .A0(n13229), .A1(n13223), .B0(n692), .B1(n6472), .Y(n13261)
         );
  AOI22XL U3648 ( .A0(n12914), .A1(n12908), .B0(n696), .B1(n6815), .Y(n12946)
         );
  AOI22XL U3649 ( .A0(n12599), .A1(n12593), .B0(n694), .B1(n6775), .Y(n12631)
         );
  AOI22XL U3650 ( .A0(n13544), .A1(n13538), .B0(n695), .B1(n6519), .Y(n13576)
         );
  AOI22XL U3651 ( .A0(n12284), .A1(n12278), .B0(n691), .B1(n6530), .Y(n12315)
         );
  AOI22XL U3652 ( .A0(n11652), .A1(n11646), .B0(n689), .B1(n6826), .Y(n11684)
         );
  AOI22XL U3653 ( .A0(top_core_KE_sb1_n77), .A1(top_core_KE_sb1_n71), .B0(n690), .B1(n6804), .Y(top_core_KE_sb1_n109) );
  AOI22XL U3654 ( .A0(n11968), .A1(n11962), .B0(n693), .B1(n6507), .Y(n12000)
         );
  OAI211XL U3655 ( .A0(n11736), .A1(n50), .B0(n11737), .C0(n11738), .Y(n11721)
         );
  OAI211XL U3656 ( .A0(top_core_KE_sb1_n163), .A1(n51), .B0(
        top_core_KE_sb1_n164), .C0(top_core_KE_sb1_n165), .Y(
        top_core_KE_sb1_n148) );
  OAI211XL U3657 ( .A0(n12367), .A1(n89), .B0(n12368), .C0(n12369), .Y(n12352)
         );
  OAI211XL U3658 ( .A0(n12052), .A1(n53), .B0(n12053), .C0(n12054), .Y(n12037)
         );
  OAI211XL U3659 ( .A0(n12683), .A1(n54), .B0(n12684), .C0(n12685), .Y(n12668)
         );
  OAI211XL U3660 ( .A0(n12998), .A1(n56), .B0(n12999), .C0(n13000), .Y(n12983)
         );
  OAI211XL U3661 ( .A0(n13628), .A1(n55), .B0(n13629), .C0(n13630), .Y(n13613)
         );
  OAI211XL U3662 ( .A0(n13313), .A1(n52), .B0(n13314), .C0(n13315), .Y(n13298)
         );
  OAI211XL U3663 ( .A0(n11716), .A1(n1257), .B0(n11720), .C0(n11804), .Y(
        n11803) );
  OAI211XL U3664 ( .A0(top_core_KE_sb1_n143), .A1(n1329), .B0(
        top_core_KE_sb1_n147), .C0(top_core_KE_sb1_n232), .Y(
        top_core_KE_sb1_n231) );
  OAI211XL U3665 ( .A0(n12347), .A1(n1264), .B0(n12351), .C0(n12435), .Y(
        n12434) );
  OAI211XL U3666 ( .A0(n12032), .A1(n1260), .B0(n12036), .C0(n12120), .Y(
        n12119) );
  AOI32XL U3667 ( .A0(n1342), .A1(n1267), .A2(n6779), .B0(n6778), .B1(n12838), 
        .Y(n12837) );
  AOI211XL U3668 ( .A0(n1188), .A1(n12598), .B0(n12763), .C0(n6840), .Y(n12839) );
  AOI32XL U3669 ( .A0(n1369), .A1(n1276), .A2(n6522), .B0(n6433), .B1(n13783), 
        .Y(n13782) );
  AOI211XL U3670 ( .A0(n1157), .A1(n13543), .B0(n13708), .C0(n6593), .Y(n13784) );
  AOI32XL U3671 ( .A0(n1355), .A1(n1270), .A2(n6818), .B0(n6714), .B1(n13153), 
        .Y(n13152) );
  AOI211XL U3672 ( .A0(n1197), .A1(n12913), .B0(n13078), .C0(n6886), .Y(n13154) );
  AOI32XL U3673 ( .A0(n1354), .A1(n11661), .A2(n6829), .B0(n6745), .B1(n11892), 
        .Y(n11891) );
  AOI211XL U3674 ( .A0(n1202), .A1(n11651), .B0(n11817), .C0(n6910), .Y(n11893) );
  AOI32XL U3675 ( .A0(n1343), .A1(top_core_KE_sb1_n86), .A2(n6808), .B0(n6807), 
        .B1(top_core_KE_sb1_n321), .Y(top_core_KE_sb1_n320) );
  AOI211XL U3676 ( .A0(n1193), .A1(top_core_KE_sb1_n76), .B0(
        top_core_KE_sb1_n245), .C0(n6864), .Y(top_core_KE_sb1_n322) );
  AOI32XL U3677 ( .A0(n1368), .A1(n1264), .A2(n6533), .B0(n6442), .B1(n12523), 
        .Y(n12522) );
  AOI211XL U3678 ( .A0(n1162), .A1(n12283), .B0(n12448), .C0(n6617), .Y(n12524) );
  AOI32XL U3679 ( .A0(n1357), .A1(n11977), .A2(n6511), .B0(n6510), .B1(n12208), 
        .Y(n12207) );
  AOI211XL U3680 ( .A0(n1153), .A1(n11967), .B0(n12133), .C0(n6570), .Y(n12209) );
  AOI32XL U3681 ( .A0(n1356), .A1(n1273), .A2(n6476), .B0(n6475), .B1(n13468), 
        .Y(n13467) );
  AOI211XL U3682 ( .A0(n1148), .A1(n13228), .B0(n13393), .C0(n6545), .Y(n13469) );
  NAND3XL U3683 ( .A(n1739), .B(n12716), .C(n6775), .Y(n12771) );
  NAND3XL U3684 ( .A(n1710), .B(n13031), .C(n6815), .Y(n13086) );
  NAND3XL U3685 ( .A(n1681), .B(n13346), .C(n6472), .Y(n13401) );
  AOI222XL U3686 ( .A0(n6909), .A1(n1258), .B0(n11701), .B1(n689), .C0(n6920), 
        .C1(n1221), .Y(n11789) );
  NAND3XL U3687 ( .A(n11769), .B(n11705), .C(n1344), .Y(n11788) );
  AOI222XL U3688 ( .A0(n6863), .A1(n1330), .B0(top_core_KE_sb1_n126), .B1(n690), .C0(n6874), .C1(n1215), .Y(top_core_KE_sb1_n217) );
  NAND3XL U3689 ( .A(top_core_KE_sb1_n197), .B(top_core_KE_sb1_n130), .C(n1345), .Y(top_core_KE_sb1_n216) );
  AOI222XL U3690 ( .A0(n6616), .A1(n1265), .B0(n12332), .B1(n691), .C0(n6627), 
        .C1(n1183), .Y(n12420) );
  NAND3XL U3691 ( .A(n12400), .B(n12336), .C(n1358), .Y(n12419) );
  AOI222XL U3692 ( .A0(n6569), .A1(n1261), .B0(n12017), .B1(n693), .C0(n6580), 
        .C1(n1175), .Y(n12105) );
  NAND3XL U3693 ( .A(n12085), .B(n12021), .C(n1359), .Y(n12104) );
  NAND3XL U3694 ( .A(n1652), .B(n13661), .C(n6519), .Y(n13716) );
  AOI221XL U3695 ( .A0(n6627), .A1(n1761), .B0(n6533), .B1(n12278), .C0(n12279), .Y(n12277) );
  AOI31XL U3696 ( .A0(n12283), .A1(n1169), .A2(n12284), .B0(n12285), .Y(n12276) );
  NAND3XL U3697 ( .A(n1344), .B(n11705), .C(n714), .Y(n11809) );
  NAND3XL U3698 ( .A(n1345), .B(top_core_KE_sb1_n130), .C(n715), .Y(
        top_core_KE_sb1_n237) );
  NAND3XL U3699 ( .A(n1358), .B(n12336), .C(n716), .Y(n12440) );
  NAND3XL U3700 ( .A(n1359), .B(n12021), .C(n718), .Y(n12125) );
  NAND3XL U3701 ( .A(n1761), .B(n12400), .C(n6530), .Y(n12456) );
  NAND3XL U3702 ( .A(n1803), .B(n11769), .C(n6826), .Y(n11825) );
  NAND3XL U3703 ( .A(n1824), .B(top_core_KE_sb1_n197), .C(n6804), .Y(
        top_core_KE_sb1_n254) );
  NAND3XL U3704 ( .A(n1782), .B(n12085), .C(n6507), .Y(n12141) );
  AOI221XL U3705 ( .A0(n6920), .A1(n1803), .B0(n6829), .B1(n11646), .C0(n11647), .Y(n11645) );
  AOI31XL U3706 ( .A0(n11651), .A1(n1209), .A2(n11652), .B0(n11653), .Y(n11644) );
  AOI221XL U3707 ( .A0(n6874), .A1(n1824), .B0(n6808), .B1(top_core_KE_sb1_n71), .C0(top_core_KE_sb1_n72), .Y(top_core_KE_sb1_n70) );
  AOI31XL U3708 ( .A0(top_core_KE_sb1_n76), .A1(n1207), .A2(
        top_core_KE_sb1_n77), .B0(top_core_KE_sb1_n78), .Y(top_core_KE_sb1_n69) );
  AOI221XL U3709 ( .A0(n6580), .A1(n1782), .B0(n6511), .B1(n11962), .C0(n11963), .Y(n11961) );
  AOI31XL U3710 ( .A0(n11967), .A1(n1167), .A2(n11968), .B0(n11969), .Y(n11960) );
  AOI221XL U3711 ( .A0(n6556), .A1(n1681), .B0(n6476), .B1(n13223), .C0(n13224), .Y(n13222) );
  AOI31XL U3712 ( .A0(n13228), .A1(n1166), .A2(n13229), .B0(n13230), .Y(n13221) );
  AOI221XL U3713 ( .A0(n6897), .A1(n1710), .B0(n6818), .B1(n12908), .C0(n12909), .Y(n12907) );
  AOI31XL U3714 ( .A0(n12913), .A1(n1208), .A2(n12914), .B0(n12915), .Y(n12906) );
  AOI221XL U3715 ( .A0(n6851), .A1(n1739), .B0(n6779), .B1(n12593), .C0(n12594), .Y(n12592) );
  AOI31XL U3716 ( .A0(n12598), .A1(n1206), .A2(n12599), .B0(n12600), .Y(n12591) );
  AOI221XL U3717 ( .A0(n6604), .A1(n1652), .B0(n6522), .B1(n13538), .C0(n13539), .Y(n13537) );
  AOI31XL U3718 ( .A0(n13543), .A1(n1168), .A2(n13544), .B0(n13545), .Y(n13536) );
  AOI211XL U3719 ( .A0(n6909), .A1(n1259), .B0(n11760), .C0(n11761), .Y(n11759) );
  AOI211XL U3720 ( .A0(n6863), .A1(n1331), .B0(top_core_KE_sb1_n188), .C0(
        top_core_KE_sb1_n189), .Y(top_core_KE_sb1_n187) );
  AOI211XL U3721 ( .A0(n6569), .A1(n1262), .B0(n12076), .C0(n12077), .Y(n12075) );
  AOI222XL U3722 ( .A0(top_core_io_CORE_FULL), .A1(n4132), .B0(
        top_core_io_n188), .B1(top_core_io_operation), .C0(top_core_io_n177), 
        .C1(top_core_io_NK_0_), .Y(top_core_io_n661) );
  OAI22XL U3723 ( .A0(n6308), .A1(top_core_EC_n1026), .B0(top_core_EC_n25), 
        .B1(n1), .Y(top_core_EC_n1294) );
  OAI22XL U3724 ( .A0(n7004), .A1(n151), .B0(n1500), .B1(top_core_KE_n2711), 
        .Y(top_core_KE_n4926) );
  OAI22XL U3725 ( .A0(n7001), .A1(n151), .B0(n1500), .B1(top_core_KE_n2708), 
        .Y(top_core_KE_n4923) );
  CLKINVX3 U3726 ( .A(n2887), .Y(n2881) );
  CLKINVX3 U3727 ( .A(n3485), .Y(n3482) );
  CLKINVX3 U3728 ( .A(n2642), .Y(n2639) );
  CLKINVX3 U3729 ( .A(n3243), .Y(n3241) );
  CLKINVX3 U3730 ( .A(n3005), .Y(n3003) );
  CLKINVX3 U3731 ( .A(n2704), .Y(n2700) );
  CLKINVX3 U3732 ( .A(n3184), .Y(n3180) );
  CLKINVX3 U3733 ( .A(n3367), .Y(n3363) );
  CLKINVX3 U3734 ( .A(n3065), .Y(n3061) );
  CLKINVX3 U3735 ( .A(n2582), .Y(n2578) );
  CLKINVX3 U3736 ( .A(n2764), .Y(n2760) );
  CLKINVX3 U3737 ( .A(n3424), .Y(n3421) );
  CLKINVX3 U3738 ( .A(n2946), .Y(n2942) );
  CLKINVX3 U3739 ( .A(n3126), .Y(n3122) );
  CLKINVX3 U3740 ( .A(n2825), .Y(n2821) );
  CLKINVX3 U3741 ( .A(n3304), .Y(n3302) );
  XOR2X1 U3742 ( .A(n1548), .B(top_core_EC_mix_in[11]), .Y(
        top_core_EC_mc_mix_in_8[14]) );
  XOR2X1 U3743 ( .A(n1548), .B(top_core_EC_mix_in[8]), .Y(
        top_core_EC_mc_mix_in_4_10_) );
  XOR2X1 U3744 ( .A(n1545), .B(top_core_EC_mix_in[24]), .Y(
        top_core_EC_mc_mix_in_4_26_) );
  XOR2X1 U3745 ( .A(n1545), .B(top_core_EC_mix_in[27]), .Y(
        top_core_EC_mc_mix_in_8[30]) );
  CLKINVX3 U3746 ( .A(n1764), .Y(n1760) );
  CLKINVX3 U3747 ( .A(n1656), .Y(n1651) );
  CLKINVX3 U3748 ( .A(n1806), .Y(n1802) );
  CLKINVX3 U3749 ( .A(n1827), .Y(n1823) );
  CLKINVX3 U3750 ( .A(n1785), .Y(n1781) );
  CLKINVX3 U3751 ( .A(n1690), .Y(n1687) );
  CLKINVX3 U3752 ( .A(n1719), .Y(n1716) );
  CLKINVX3 U3753 ( .A(n1748), .Y(n1745) );
  CLKINVX3 U3754 ( .A(n1769), .Y(n1767) );
  CLKINVX3 U3755 ( .A(n1662), .Y(n1658) );
  CLKINVX3 U3756 ( .A(n1743), .Y(n1738) );
  CLKINVX3 U3757 ( .A(n1714), .Y(n1709) );
  CLKINVX3 U3758 ( .A(n1685), .Y(n1680) );
  CLKINVX3 U3759 ( .A(n1814), .Y(n1809) );
  CLKINVX3 U3760 ( .A(n1835), .Y(n1830) );
  CLKINVX3 U3761 ( .A(n1793), .Y(n1788) );
  OAI22X1 U3762 ( .A0(n2421), .A1(top_core_EC_ss_n213), .B0(n2369), .B1(n4841), 
        .Y(top_core_EC_mix_in[24]) );
  OAI22X1 U3763 ( .A0(n2481), .A1(top_core_EC_ss_n210), .B0(n2369), .B1(n4847), 
        .Y(top_core_EC_mix_in[27]) );
  OAI22X1 U3764 ( .A0(n2437), .A1(top_core_EC_ss_n178), .B0(n2371), .B1(n5233), 
        .Y(top_core_EC_mix_in[56]) );
  OAI22X1 U3765 ( .A0(n2434), .A1(top_core_EC_ss_n186), .B0(n2371), .B1(n4963), 
        .Y(top_core_EC_mc_mix_in_2_50_) );
  OAI22X1 U3766 ( .A0(n2453), .A1(top_core_EC_ss_n203), .B0(n2369), .B1(n5789), 
        .Y(top_core_EC_mc_mix_in_2_34_) );
  OAI22X1 U3767 ( .A0(n2422), .A1(top_core_EC_ss_n211), .B0(n2369), .B1(n4848), 
        .Y(top_core_EC_mix_in[26]) );
  OAI22X1 U3768 ( .A0(n2459), .A1(top_core_EC_ss_n218), .B0(n2368), .B1(n6102), 
        .Y(top_core_EC_mc_mix_in_2_2_) );
  OAI22X1 U3769 ( .A0(n2403), .A1(top_core_EC_ss_n221), .B0(n2368), .B1(n5317), 
        .Y(top_core_EC_mc_mix_in_2_18_) );
  XOR2X1 U3770 ( .A(n1536), .B(top_core_EC_mix_in[72]), .Y(
        top_core_EC_mc_mix_in_4_74_) );
  XOR2X1 U3771 ( .A(n1554), .B(top_core_EC_mix_in[104]), .Y(
        top_core_EC_mc_mix_in_4_106_) );
  XOR2X1 U3772 ( .A(n1536), .B(top_core_EC_mix_in[75]), .Y(
        top_core_EC_mc_mix_in_8[78]) );
  XOR2X1 U3773 ( .A(n1554), .B(top_core_EC_mix_in[107]), .Y(
        top_core_EC_mc_mix_in_8[110]) );
  XOR2X1 U3774 ( .A(n1539), .B(top_core_EC_mix_in[56]), .Y(
        top_core_EC_mc_mix_in_4_58_) );
  XOR2X1 U3775 ( .A(n1533), .B(top_core_EC_mix_in[88]), .Y(
        top_core_EC_mc_mix_in_4_90_) );
  XOR2X1 U3776 ( .A(n1551), .B(top_core_EC_mix_in[120]), .Y(
        top_core_EC_mc_mix_in_4_122_) );
  XOR2X1 U3777 ( .A(n1539), .B(top_core_EC_mix_in[59]), .Y(
        top_core_EC_mc_mix_in_8[62]) );
  XOR2X1 U3778 ( .A(n1533), .B(top_core_EC_mix_in[91]), .Y(
        top_core_EC_mc_mix_in_8[94]) );
  XOR2X1 U3779 ( .A(n1551), .B(top_core_EC_mix_in[123]), .Y(
        top_core_EC_mc_mix_in_8[126]) );
  BUFX3 U3780 ( .A(n5386), .Y(n1000) );
  BUFX3 U3781 ( .A(n5032), .Y(n944) );
  BUFX3 U3782 ( .A(n5858), .Y(n1084) );
  BUFX3 U3783 ( .A(n6170), .Y(n1140) );
  BUFX3 U3784 ( .A(n5116), .Y(n958) );
  BUFX3 U3785 ( .A(n6086), .Y(n1126) );
  BUFX3 U3786 ( .A(n5622), .Y(n1042) );
  BUFX3 U3787 ( .A(n5302), .Y(n986) );
  BUFX3 U3788 ( .A(n5546), .Y(n1028) );
  BUFX3 U3789 ( .A(n5774), .Y(n1070) );
  BUFX3 U3790 ( .A(n6010), .Y(n1112) );
  BUFX3 U3791 ( .A(n4916), .Y(n930) );
  BUFX3 U3792 ( .A(n5224), .Y(n972) );
  BUFX3 U3793 ( .A(n5470), .Y(n1014) );
  BUFX3 U3794 ( .A(n5698), .Y(n1056) );
  BUFX3 U3795 ( .A(n5934), .Y(n1098) );
  OAI22X1 U3796 ( .A0(n2454), .A1(top_core_EC_ss_n175), .B0(n2372), .B1(n193), 
        .Y(top_core_EC_mix_in[59]) );
  OAI22X1 U3797 ( .A0(n2534), .A1(top_core_EC_ss_n143), .B0(n2374), .B1(n211), 
        .Y(top_core_EC_mix_in[88]) );
  OAI22X1 U3798 ( .A0(n2533), .A1(top_core_EC_ss_n139), .B0(n2374), .B1(n213), 
        .Y(top_core_EC_mix_in[91]) );
  OAI22X1 U3799 ( .A0(n2541), .A1(top_core_EC_ss_n234), .B0(n2389), .B1(n231), 
        .Y(top_core_EC_mix_in[120]) );
  OAI22X1 U3800 ( .A0(n2540), .A1(top_core_EC_ss_n231), .B0(n2511), .B1(n233), 
        .Y(top_core_EC_mix_in[123]) );
  OAI22X1 U3801 ( .A0(n2469), .A1(top_core_EC_ss_n168), .B0(n2372), .B1(n198), 
        .Y(top_core_EC_mc_mix_in_2_66_) );
  OAI22X1 U3802 ( .A0(n2405), .A1(top_core_EC_ss_n140), .B0(n2374), .B1(n212), 
        .Y(top_core_EC_mix_in[90]) );
  OAI22X1 U3803 ( .A0(n2427), .A1(top_core_EC_ss_n242), .B0(n2381), .B1(n228), 
        .Y(top_core_EC_mc_mix_in_2_114_) );
  OAI22X1 U3804 ( .A0(n2437), .A1(top_core_EC_ss_n176), .B0(n2371), .B1(n192), 
        .Y(top_core_EC_mix_in[58]) );
  OAI22X1 U3805 ( .A0(n2530), .A1(top_core_EC_ss_n232), .B0(n2520), .B1(n232), 
        .Y(top_core_EC_mix_in[122]) );
  OAI22X1 U3806 ( .A0(n2488), .A1(top_core_EC_ss_n150), .B0(n2373), .B1(n208), 
        .Y(top_core_EC_mc_mix_in_2_82_) );
  OAI22X1 U3807 ( .A0(n2402), .A1(top_core_EC_ss_n133), .B0(n2375), .B1(n218), 
        .Y(top_core_EC_mc_mix_in_2_98_) );
  NAND2X1 U3808 ( .A(n1517), .B(n3473), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n218) );
  NAND2X1 U3809 ( .A(n1505), .B(n2872), .Y(n10032) );
  NAND2X1 U3810 ( .A(n1529), .B(n2630), .Y(n11200) );
  NAND2X1 U3811 ( .A(n1519), .B(n3232), .Y(n8280) );
  NAND2X1 U3812 ( .A(n1531), .B(n2691), .Y(n10908) );
  NAND2X1 U3813 ( .A(n1512), .B(n3052), .Y(n9156) );
  NAND2X1 U3814 ( .A(n1527), .B(n3412), .Y(n7404) );
  NAND2X1 U3815 ( .A(n1503), .B(n2812), .Y(n10324) );
  NAND2X1 U3816 ( .A(n1510), .B(n2994), .Y(n9448) );
  NAND2X1 U3817 ( .A(n1516), .B(n3171), .Y(n8572) );
  NAND2X1 U3818 ( .A(n1523), .B(n3354), .Y(n7696) );
  NAND2X1 U3819 ( .A(n1526), .B(n2569), .Y(n11492) );
  NAND2X1 U3820 ( .A(n1501), .B(n2751), .Y(n10616) );
  NAND2X1 U3821 ( .A(n1508), .B(n2933), .Y(n9740) );
  NAND2X1 U3822 ( .A(n1514), .B(n3113), .Y(n8864) );
  NAND2X1 U3823 ( .A(n1521), .B(n3293), .Y(n7988) );
  INVX1 U3824 ( .A(n13310), .Y(n6552) );
  INVX1 U3825 ( .A(n12680), .Y(n6847) );
  INVX1 U3826 ( .A(n12995), .Y(n6893) );
  INVX1 U3827 ( .A(n12364), .Y(n6624) );
  INVX1 U3828 ( .A(n11733), .Y(n6917) );
  INVX1 U3829 ( .A(top_core_KE_sb1_n160), .Y(n6871) );
  INVX1 U3830 ( .A(n12049), .Y(n6577) );
  INVX1 U3831 ( .A(n13625), .Y(n6600) );
  INVX1 U3832 ( .A(top_core_KE_prev_key1_reg_89_), .Y(n1654) );
  BUFX4 U3833 ( .A(n6677), .Y(n1171) );
  INVX1 U3834 ( .A(n1370), .Y(n6358) );
  NAND3X1 U3835 ( .A(n_WR), .B(n_ADDR[6]), .C(n4124), .Y(top_core_io_n5) );
  BUFX3 U3836 ( .A(top_core_KE_prev_key1_reg_71_), .Y(n1336) );
  BUFX3 U3837 ( .A(top_core_KE_prev_key1_reg_79_), .Y(n1337) );
  BUFX3 U3838 ( .A(top_core_KE_prev_key1_reg_30_), .Y(n1368) );
  BUFX3 U3839 ( .A(top_core_KE_prev_key1_reg_87_), .Y(n1340) );
  BUFX3 U3840 ( .A(top_core_KE_prev_key1_reg_95_), .Y(n1341) );
  BUFX3 U3841 ( .A(top_core_KE_prev_key1_reg_14_), .Y(n1354) );
  BUFX3 U3842 ( .A(top_core_KE_prev_key1_reg_6_), .Y(n1343) );
  BUFX3 U3843 ( .A(top_core_KE_prev_key1_reg_22_), .Y(n1357) );
  NOR3X1 U3844 ( .A(n7013), .B(n1334), .C(top_core_KE_n728), .Y(
        top_core_KE_n1866) );
  BUFX4 U3845 ( .A(top_core_KE_prev_key1_reg_26_), .Y(n1358) );
  BUFX4 U3846 ( .A(top_core_KE_prev_key1_reg_76_), .Y(n1351) );
  BUFX4 U3847 ( .A(top_core_KE_prev_key1_reg_68_), .Y(n1353) );
  BUFX4 U3848 ( .A(top_core_KE_prev_key1_reg_84_), .Y(n1367) );
  BUFX4 U3849 ( .A(top_core_KE_prev_key1_reg_10_), .Y(n1344) );
  BUFX4 U3850 ( .A(top_core_KE_prev_key1_reg_2_), .Y(n1345) );
  BUFX4 U3851 ( .A(top_core_KE_prev_key1_reg_18_), .Y(n1359) );
  BUFX4 U3852 ( .A(top_core_KE_prev_key1_reg_92_), .Y(n1365) );
  XNOR2X1 U3853 ( .A(top_core_KE_n635), .B(top_core_KE_prev_key0_reg_119_), 
        .Y(top_core_KE_n1925) );
  XNOR2X1 U3854 ( .A(top_core_KE_n636), .B(top_core_KE_prev_key0_reg_118_), 
        .Y(top_core_KE_n1927) );
  XNOR2X1 U3855 ( .A(top_core_KE_n637), .B(top_core_KE_prev_key0_reg_117_), 
        .Y(top_core_KE_n1929) );
  XNOR2X1 U3856 ( .A(top_core_KE_n638), .B(top_core_KE_prev_key0_reg_116_), 
        .Y(top_core_KE_n1931) );
  XNOR2X1 U3857 ( .A(top_core_KE_n639), .B(top_core_KE_prev_key0_reg_115_), 
        .Y(top_core_KE_n1933) );
  XNOR2X1 U3858 ( .A(top_core_KE_n640), .B(top_core_KE_prev_key0_reg_114_), 
        .Y(top_core_KE_n1935) );
  XNOR2X1 U3859 ( .A(top_core_KE_n641), .B(top_core_KE_prev_key0_reg_113_), 
        .Y(top_core_KE_n1937) );
  XNOR2X1 U3860 ( .A(top_core_KE_n642), .B(top_core_KE_prev_key0_reg_112_), 
        .Y(top_core_KE_n1939) );
  XNOR2X1 U3861 ( .A(top_core_KE_n643), .B(top_core_KE_prev_key0_reg_111_), 
        .Y(top_core_KE_n1941) );
  XNOR2X1 U3862 ( .A(top_core_KE_n644), .B(top_core_KE_prev_key0_reg_110_), 
        .Y(top_core_KE_n1943) );
  XNOR2X1 U3863 ( .A(top_core_KE_n645), .B(top_core_KE_prev_key0_reg_109_), 
        .Y(top_core_KE_n1945) );
  XNOR2X1 U3864 ( .A(top_core_KE_n646), .B(top_core_KE_prev_key0_reg_108_), 
        .Y(top_core_KE_n1947) );
  XNOR2X1 U3865 ( .A(top_core_KE_n647), .B(top_core_KE_prev_key0_reg_107_), 
        .Y(top_core_KE_n1949) );
  XNOR2X1 U3866 ( .A(top_core_KE_n648), .B(top_core_KE_prev_key0_reg_106_), 
        .Y(top_core_KE_n1951) );
  XNOR2X1 U3867 ( .A(top_core_KE_n649), .B(top_core_KE_prev_key0_reg_105_), 
        .Y(top_core_KE_n1953) );
  XNOR2X1 U3868 ( .A(top_core_KE_n650), .B(top_core_KE_prev_key0_reg_104_), 
        .Y(top_core_KE_n1955) );
  XNOR2X1 U3869 ( .A(top_core_KE_n651), .B(top_core_KE_prev_key0_reg_103_), 
        .Y(top_core_KE_n1957) );
  XNOR2X1 U3870 ( .A(top_core_KE_n652), .B(top_core_KE_prev_key0_reg_102_), 
        .Y(top_core_KE_n1959) );
  XNOR2X1 U3871 ( .A(top_core_KE_n653), .B(top_core_KE_prev_key0_reg_101_), 
        .Y(top_core_KE_n1961) );
  XNOR2X1 U3872 ( .A(top_core_KE_n654), .B(top_core_KE_prev_key0_reg_100_), 
        .Y(top_core_KE_n1963) );
  XNOR2X1 U3873 ( .A(top_core_KE_n655), .B(top_core_KE_prev_key0_reg_99_), .Y(
        top_core_KE_n1965) );
  XNOR2X1 U3874 ( .A(top_core_KE_n656), .B(top_core_KE_prev_key0_reg_98_), .Y(
        top_core_KE_n1967) );
  XNOR2X1 U3875 ( .A(top_core_KE_n657), .B(top_core_KE_prev_key0_reg_97_), .Y(
        top_core_KE_n1969) );
  XNOR2X1 U3876 ( .A(top_core_KE_n658), .B(top_core_KE_prev_key0_reg_96_), .Y(
        top_core_KE_n1971) );
  XNOR2X1 U3877 ( .A(top_core_KE_prev_key0_reg_95_), .B(n6341), .Y(
        top_core_KE_n1909) );
  XNOR2X1 U3878 ( .A(top_core_KE_prev_key0_reg_89_), .B(n6314), .Y(
        top_core_KE_n1921) );
  XNOR2X1 U3879 ( .A(top_core_KE_prev_key0_reg_88_), .B(n6695), .Y(
        top_core_KE_n1923) );
  XNOR2X1 U3880 ( .A(top_core_KE_prev_key0_reg_90_), .B(n6674), .Y(
        top_core_KE_n1919) );
  XNOR2X1 U3881 ( .A(top_core_KE_prev_key0_reg_91_), .B(n6655), .Y(
        top_core_KE_n1917) );
  XNOR2X1 U3882 ( .A(top_core_KE_prev_key0_reg_92_), .B(n6607), .Y(
        top_core_KE_n1915) );
  XNOR2X1 U3883 ( .A(top_core_KE_prev_key0_reg_93_), .B(n6524), .Y(
        top_core_KE_n1913) );
  XNOR2X1 U3884 ( .A(top_core_KE_prev_key0_reg_94_), .B(n6435), .Y(
        top_core_KE_n1911) );
  INVX1 U3885 ( .A(top_core_KE_prev_key0_reg_112_), .Y(n6689) );
  INVX1 U3886 ( .A(top_core_KE_prev_key0_reg_113_), .Y(n6682) );
  INVX1 U3887 ( .A(top_core_KE_prev_key0_reg_114_), .Y(n6667) );
  INVX1 U3888 ( .A(top_core_KE_prev_key0_reg_115_), .Y(n6639) );
  INVX1 U3889 ( .A(top_core_KE_prev_key0_reg_116_), .Y(n6560) );
  INVX1 U3890 ( .A(top_core_KE_prev_key0_reg_117_), .Y(n6480) );
  INVX1 U3891 ( .A(top_core_KE_prev_key0_reg_118_), .Y(n6402) );
  INVX1 U3892 ( .A(top_core_KE_prev_key0_reg_119_), .Y(n6394) );
  NOR2X2 U3893 ( .A(n4143), .B(n4138), .Y(n304) );
  BUFX3 U3894 ( .A(n385), .Y(n1144) );
  BUFX3 U3895 ( .A(n386), .Y(n1005) );
  BUFX3 U3896 ( .A(n387), .Y(n949) );
  BUFX3 U3897 ( .A(n388), .Y(n1089) );
  BUFX3 U3898 ( .A(n389), .Y(n1075) );
  BUFX3 U3899 ( .A(n391), .Y(n1019) );
  BUFX3 U3900 ( .A(n390), .Y(n935) );
  BUFX3 U3901 ( .A(n392), .Y(n1103) );
  BUFX3 U3902 ( .A(n393), .Y(n1033) );
  BUFX3 U3903 ( .A(n394), .Y(n963) );
  BUFX3 U3904 ( .A(n395), .Y(n1117) );
  BUFX3 U3905 ( .A(n396), .Y(n1047) );
  BUFX3 U3906 ( .A(n397), .Y(n977) );
  BUFX3 U3907 ( .A(n398), .Y(n1131) );
  BUFX3 U3908 ( .A(n399), .Y(n1061) );
  BUFX3 U3909 ( .A(n400), .Y(n991) );
  BUFX3 U3910 ( .A(n353), .Y(n1004) );
  BUFX3 U3911 ( .A(n354), .Y(n1145) );
  BUFX3 U3912 ( .A(n356), .Y(n948) );
  BUFX3 U3913 ( .A(n355), .Y(n1088) );
  BUFX3 U3914 ( .A(n357), .Y(n962) );
  BUFX3 U3915 ( .A(n359), .Y(n1046) );
  BUFX3 U3916 ( .A(n358), .Y(n1130) );
  BUFX3 U3917 ( .A(n360), .Y(n990) );
  BUFX3 U3918 ( .A(n361), .Y(n1032) );
  BUFX3 U3919 ( .A(n362), .Y(n1074) );
  BUFX3 U3920 ( .A(n363), .Y(n1116) );
  BUFX3 U3921 ( .A(n364), .Y(n934) );
  BUFX3 U3922 ( .A(n365), .Y(n976) );
  BUFX3 U3923 ( .A(n366), .Y(n1018) );
  BUFX3 U3924 ( .A(n367), .Y(n1060) );
  BUFX3 U3925 ( .A(n368), .Y(n1102) );
  NAND2X1 U3926 ( .A(n5371), .B(n353), .Y(n9905) );
  NAND2X1 U3927 ( .A(n6161), .B(n354), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n88) );
  NAND2X1 U3928 ( .A(n5843), .B(n355), .Y(n8153) );
  NAND2X1 U3929 ( .A(n5017), .B(n356), .Y(n11073) );
  NAND2X1 U3930 ( .A(n5101), .B(n357), .Y(n10781) );
  NAND2X1 U3931 ( .A(n6071), .B(n358), .Y(n7277) );
  NAND2X1 U3932 ( .A(n5607), .B(n359), .Y(n9029) );
  NAND2X1 U3933 ( .A(n5287), .B(n360), .Y(n10197) );
  NAND2X1 U3934 ( .A(n5531), .B(n361), .Y(n9321) );
  NAND2X1 U3935 ( .A(n5759), .B(n362), .Y(n8445) );
  NAND2X1 U3936 ( .A(n5995), .B(n363), .Y(n7569) );
  NAND2X1 U3937 ( .A(n4901), .B(n364), .Y(n11365) );
  NAND2X1 U3938 ( .A(n5209), .B(n365), .Y(n10489) );
  NAND2X1 U3939 ( .A(n5455), .B(n366), .Y(n9613) );
  NAND2X1 U3940 ( .A(n5683), .B(n367), .Y(n8737) );
  NAND2X1 U3941 ( .A(n5919), .B(n368), .Y(n7861) );
  CLKINVX3 U3942 ( .A(n17030), .Y(n5330) );
  CLKINVX3 U3943 ( .A(n13880), .Y(n6114) );
  CLKINVX3 U3944 ( .A(n18290), .Y(n4976) );
  CLKINVX3 U3945 ( .A(n15140), .Y(n5802) );
  CLKINVX3 U3946 ( .A(n15455), .Y(n5718) );
  CLKINVX3 U3947 ( .A(n18605), .Y(n4860) );
  CLKINVX3 U3948 ( .A(n16715), .Y(n5414) );
  CLKINVX3 U3949 ( .A(n14825), .Y(n5878) );
  CLKINVX3 U3950 ( .A(n16400), .Y(n5490) );
  CLKINVX3 U3951 ( .A(n17975), .Y(n5060) );
  CLKINVX3 U3952 ( .A(n14510), .Y(n5954) );
  CLKINVX3 U3953 ( .A(n16085), .Y(n5566) );
  CLKINVX3 U3954 ( .A(n17660), .Y(n5168) );
  CLKINVX3 U3955 ( .A(n14195), .Y(n6030) );
  CLKINVX3 U3956 ( .A(n15770), .Y(n5642) );
  CLKINVX3 U3957 ( .A(n17345), .Y(n5246) );
  CLKINVX3 U3958 ( .A(n3609), .Y(n3584) );
  CLKINVX3 U3959 ( .A(n3611), .Y(n3582) );
  CLKINVX3 U3960 ( .A(n3591), .Y(n3583) );
  CLKINVX3 U3961 ( .A(n3600), .Y(n3585) );
  CLKINVX3 U3962 ( .A(n3606), .Y(n3586) );
  CLKINVX3 U3963 ( .A(n1281), .Y(n1625) );
  CLKINVX3 U3964 ( .A(n1311), .Y(n1615) );
  CLKINVX3 U3965 ( .A(n1323), .Y(n1611) );
  CLKINVX3 U3966 ( .A(n1293), .Y(n1621) );
  CLKINVX3 U3967 ( .A(n1320), .Y(n1612) );
  CLKINVX3 U3968 ( .A(n1302), .Y(n1618) );
  CLKINVX3 U3969 ( .A(n1284), .Y(n1624) );
  CLKINVX3 U3970 ( .A(n1314), .Y(n1614) );
  CLKINVX3 U3971 ( .A(n1305), .Y(n1617) );
  CLKINVX3 U3972 ( .A(n1296), .Y(n1620) );
  CLKINVX3 U3973 ( .A(n1287), .Y(n1623) );
  CLKINVX3 U3974 ( .A(n1326), .Y(n1610) );
  CLKINVX3 U3975 ( .A(n1317), .Y(n1613) );
  CLKINVX3 U3976 ( .A(n1308), .Y(n1616) );
  CLKINVX3 U3977 ( .A(n1299), .Y(n1619) );
  CLKINVX3 U3978 ( .A(n1290), .Y(n1622) );
  INVX1 U3979 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n199), .Y(n6162) );
  INVX1 U3980 ( .A(n10013), .Y(n5372) );
  INVX1 U3981 ( .A(n11181), .Y(n5018) );
  INVX1 U3982 ( .A(n8261), .Y(n5844) );
  INVX1 U3983 ( .A(n10889), .Y(n5102) );
  INVX1 U3984 ( .A(n7385), .Y(n6072) );
  INVX1 U3985 ( .A(n9137), .Y(n5608) );
  INVX1 U3986 ( .A(n10305), .Y(n5288) );
  INVX1 U3987 ( .A(n9429), .Y(n5532) );
  INVX1 U3988 ( .A(n8553), .Y(n5760) );
  INVX1 U3989 ( .A(n7677), .Y(n5996) );
  INVX1 U3990 ( .A(n11473), .Y(n4902) );
  INVX1 U3991 ( .A(n10597), .Y(n5210) );
  INVX1 U3992 ( .A(n9721), .Y(n5456) );
  INVX1 U3993 ( .A(n8845), .Y(n5684) );
  INVX1 U3994 ( .A(n7969), .Y(n5920) );
  BUFX3 U3995 ( .A(n482), .Y(n1141) );
  BUFX3 U3996 ( .A(n481), .Y(n1002) );
  BUFX3 U3997 ( .A(n483), .Y(n946) );
  BUFX3 U3998 ( .A(n484), .Y(n1086) );
  BUFX3 U3999 ( .A(n490), .Y(n1072) );
  BUFX3 U4000 ( .A(n492), .Y(n932) );
  BUFX3 U4001 ( .A(n494), .Y(n1016) );
  BUFX3 U4002 ( .A(n496), .Y(n1100) );
  BUFX3 U4003 ( .A(n489), .Y(n1030) );
  BUFX3 U4004 ( .A(n485), .Y(n960) );
  BUFX3 U4005 ( .A(n491), .Y(n1114) );
  BUFX3 U4006 ( .A(n486), .Y(n1044) );
  BUFX3 U4007 ( .A(n493), .Y(n974) );
  BUFX3 U4008 ( .A(n487), .Y(n1128) );
  BUFX3 U4009 ( .A(n495), .Y(n1058) );
  BUFX3 U4010 ( .A(n488), .Y(n988) );
  INVX1 U4011 ( .A(n9957), .Y(n5346) );
  INVX1 U4012 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n142), .Y(n6142) );
  INVX1 U4013 ( .A(n8205), .Y(n5818) );
  INVX1 U4014 ( .A(n11125), .Y(n4992) );
  INVX1 U4015 ( .A(n10833), .Y(n5076) );
  INVX1 U4016 ( .A(n7329), .Y(n6046) );
  INVX1 U4017 ( .A(n9081), .Y(n5582) );
  INVX1 U4018 ( .A(n10249), .Y(n5262) );
  INVX1 U4019 ( .A(n9373), .Y(n5506) );
  INVX1 U4020 ( .A(n8497), .Y(n5734) );
  INVX1 U4021 ( .A(n7621), .Y(n5970) );
  INVX1 U4022 ( .A(n11417), .Y(n4876) );
  INVX1 U4023 ( .A(n10541), .Y(n5184) );
  INVX1 U4024 ( .A(n9665), .Y(n5430) );
  INVX1 U4025 ( .A(n8789), .Y(n5658) );
  INVX1 U4026 ( .A(n7913), .Y(n5894) );
  BUFX3 U4027 ( .A(n321), .Y(n1001) );
  BUFX3 U4028 ( .A(n322), .Y(n1143) );
  BUFX3 U4029 ( .A(n323), .Y(n945) );
  BUFX3 U4030 ( .A(n324), .Y(n1085) );
  BUFX3 U4031 ( .A(n325), .Y(n959) );
  BUFX3 U4032 ( .A(n326), .Y(n1127) );
  BUFX3 U4033 ( .A(n327), .Y(n1043) );
  BUFX3 U4034 ( .A(n328), .Y(n987) );
  BUFX3 U4035 ( .A(n329), .Y(n1029) );
  BUFX3 U4036 ( .A(n330), .Y(n1071) );
  BUFX3 U4037 ( .A(n331), .Y(n1113) );
  BUFX3 U4038 ( .A(n332), .Y(n931) );
  BUFX3 U4039 ( .A(n333), .Y(n973) );
  BUFX3 U4040 ( .A(n334), .Y(n1015) );
  BUFX3 U4041 ( .A(n335), .Y(n1057) );
  BUFX3 U4042 ( .A(n336), .Y(n1099) );
  INVX1 U4043 ( .A(n17082), .Y(n5361) );
  INVX1 U4044 ( .A(n13932), .Y(n6129) );
  INVX1 U4045 ( .A(n18342), .Y(n5007) );
  INVX1 U4046 ( .A(n15192), .Y(n5833) );
  INVX1 U4047 ( .A(n15507), .Y(n5749) );
  INVX1 U4048 ( .A(n16767), .Y(n5445) );
  INVX1 U4049 ( .A(n18657), .Y(n4891) );
  INVX1 U4050 ( .A(n14877), .Y(n5909) );
  INVX1 U4051 ( .A(n16452), .Y(n5521) );
  INVX1 U4052 ( .A(n18027), .Y(n5091) );
  INVX1 U4053 ( .A(n14562), .Y(n5985) );
  INVX1 U4054 ( .A(n16137), .Y(n5597) );
  INVX1 U4055 ( .A(n17712), .Y(n5199) );
  INVX1 U4056 ( .A(n14247), .Y(n6061) );
  INVX1 U4057 ( .A(n15822), .Y(n5673) );
  INVX1 U4058 ( .A(n17397), .Y(n5277) );
  INVX1 U4059 ( .A(n17113), .Y(n5359) );
  INVX1 U4060 ( .A(n13963), .Y(n6127) );
  INVX1 U4061 ( .A(n18373), .Y(n5005) );
  INVX1 U4062 ( .A(n15223), .Y(n5831) );
  INVX1 U4063 ( .A(n15538), .Y(n5747) );
  INVX1 U4064 ( .A(n16798), .Y(n5443) );
  INVX1 U4065 ( .A(n18688), .Y(n4889) );
  INVX1 U4066 ( .A(n14908), .Y(n5907) );
  INVX1 U4067 ( .A(n16483), .Y(n5519) );
  INVX1 U4068 ( .A(n18058), .Y(n5089) );
  INVX1 U4069 ( .A(n14593), .Y(n5983) );
  INVX1 U4070 ( .A(n16168), .Y(n5595) );
  INVX1 U4071 ( .A(n17743), .Y(n5197) );
  INVX1 U4072 ( .A(n14278), .Y(n6059) );
  INVX1 U4073 ( .A(n15853), .Y(n5671) );
  INVX1 U4074 ( .A(n17428), .Y(n5275) );
  NAND2X2 U4075 ( .A(n3472), .B(n3453), .Y(n13880) );
  NAND2X2 U4076 ( .A(n2871), .B(n2852), .Y(n17030) );
  NAND2X2 U4077 ( .A(n2629), .B(n2610), .Y(n18290) );
  NAND2X2 U4078 ( .A(n3231), .B(n3212), .Y(n15140) );
  NAND2X2 U4079 ( .A(n3170), .B(n3151), .Y(n15455) );
  NAND2X2 U4080 ( .A(n2568), .B(n2549), .Y(n18605) );
  NAND2X2 U4081 ( .A(n2932), .B(n2913), .Y(n16715) );
  NAND2X2 U4082 ( .A(n3292), .B(n3273), .Y(n14825) );
  NAND2X2 U4083 ( .A(n2993), .B(n2974), .Y(n16400) );
  NAND2X2 U4084 ( .A(n2690), .B(n2671), .Y(n17975) );
  NAND2X2 U4085 ( .A(n3353), .B(n3334), .Y(n14510) );
  NAND2X2 U4086 ( .A(n3051), .B(n3032), .Y(n16085) );
  NAND2X2 U4087 ( .A(n2750), .B(n2731), .Y(n17660) );
  NAND2X2 U4088 ( .A(n3411), .B(n3392), .Y(n14195) );
  NAND2X2 U4089 ( .A(n3112), .B(n3093), .Y(n15770) );
  NAND2X2 U4090 ( .A(n2811), .B(n2792), .Y(n17345) );
  NAND2X1 U4091 ( .A(n417), .B(n997), .Y(n17164) );
  NAND2X1 U4092 ( .A(n418), .B(n1136), .Y(n14014) );
  NAND2X1 U4093 ( .A(n420), .B(n1081), .Y(n15274) );
  NAND2X1 U4094 ( .A(n419), .B(n941), .Y(n18424) );
  NAND2X1 U4095 ( .A(n426), .B(n1067), .Y(n15589) );
  NAND2X1 U4096 ( .A(n430), .B(n1011), .Y(n16849) );
  NAND2X1 U4097 ( .A(n428), .B(n927), .Y(n18739) );
  NAND2X1 U4098 ( .A(n432), .B(n1095), .Y(n14959) );
  NAND2X1 U4099 ( .A(n425), .B(n1025), .Y(n16534) );
  NAND2X1 U4100 ( .A(n421), .B(n955), .Y(n18109) );
  NAND2X1 U4101 ( .A(n427), .B(n1109), .Y(n14644) );
  NAND2X1 U4102 ( .A(n422), .B(n1039), .Y(n16219) );
  NAND2X1 U4103 ( .A(n429), .B(n969), .Y(n17794) );
  NAND2X1 U4104 ( .A(n423), .B(n1123), .Y(n14329) );
  NAND2X1 U4105 ( .A(n431), .B(n1053), .Y(n15904) );
  NAND2X1 U4106 ( .A(n424), .B(n983), .Y(n17479) );
  NAND2X1 U4107 ( .A(n5378), .B(n1005), .Y(n17143) );
  NAND2X1 U4108 ( .A(n6149), .B(n1144), .Y(n13993) );
  NAND2X1 U4109 ( .A(n5850), .B(n1089), .Y(n15253) );
  NAND2X1 U4110 ( .A(n5024), .B(n949), .Y(n18403) );
  NAND2X1 U4111 ( .A(n5766), .B(n1075), .Y(n15568) );
  NAND2X1 U4112 ( .A(n5462), .B(n1019), .Y(n16828) );
  NAND2X1 U4113 ( .A(n4908), .B(n935), .Y(n18718) );
  NAND2X1 U4114 ( .A(n5926), .B(n1103), .Y(n14938) );
  NAND2X1 U4115 ( .A(n5538), .B(n1033), .Y(n16513) );
  NAND2X1 U4116 ( .A(n5108), .B(n963), .Y(n18088) );
  NAND2X1 U4117 ( .A(n6002), .B(n1117), .Y(n14623) );
  NAND2X1 U4118 ( .A(n5614), .B(n1047), .Y(n16198) );
  NAND2X1 U4119 ( .A(n5216), .B(n977), .Y(n17773) );
  NAND2X1 U4120 ( .A(n6078), .B(n1131), .Y(n14308) );
  NAND2X1 U4121 ( .A(n5690), .B(n1061), .Y(n15883) );
  NAND2X1 U4122 ( .A(n5294), .B(n991), .Y(n17458) );
  NAND2X1 U4123 ( .A(n993), .B(n9900), .Y(n10051) );
  NAND2X1 U4124 ( .A(n1135), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n237) );
  NAND2X1 U4125 ( .A(n937), .B(n11068), .Y(n11219) );
  NAND2X1 U4126 ( .A(n1077), .B(n8148), .Y(n8299) );
  NAND2X1 U4127 ( .A(n951), .B(n10776), .Y(n10927) );
  NAND2X1 U4128 ( .A(n1035), .B(n9024), .Y(n9175) );
  NAND2X1 U4129 ( .A(n1119), .B(n7272), .Y(n7423) );
  NAND2X1 U4130 ( .A(n979), .B(n10192), .Y(n10343) );
  NAND2X1 U4131 ( .A(n1021), .B(n9316), .Y(n9467) );
  NAND2X1 U4132 ( .A(n1063), .B(n8440), .Y(n8591) );
  NAND2X1 U4133 ( .A(n1105), .B(n7564), .Y(n7715) );
  NAND2X1 U4134 ( .A(n923), .B(n11360), .Y(n11511) );
  NAND2X1 U4135 ( .A(n965), .B(n10484), .Y(n10635) );
  NAND2X1 U4136 ( .A(n1007), .B(n9608), .Y(n9759) );
  NAND2X1 U4137 ( .A(n1049), .B(n8732), .Y(n8883) );
  NAND2X1 U4138 ( .A(n1091), .B(n7856), .Y(n8007) );
  NAND2X1 U4139 ( .A(n562), .B(n9970), .Y(n10013) );
  NAND2X1 U4140 ( .A(n561), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n199) );
  NAND2X1 U4141 ( .A(n563), .B(n11138), .Y(n11181) );
  NAND2X1 U4142 ( .A(n564), .B(n8218), .Y(n8261) );
  NAND2X1 U4143 ( .A(n565), .B(n10846), .Y(n10889) );
  NAND2X1 U4144 ( .A(n566), .B(n9094), .Y(n9137) );
  NAND2X1 U4145 ( .A(n567), .B(n7342), .Y(n7385) );
  NAND2X1 U4146 ( .A(n568), .B(n10262), .Y(n10305) );
  NAND2X1 U4147 ( .A(n569), .B(n9386), .Y(n9429) );
  NAND2X1 U4148 ( .A(n570), .B(n8510), .Y(n8553) );
  NAND2X1 U4149 ( .A(n571), .B(n7634), .Y(n7677) );
  NAND2X1 U4150 ( .A(n572), .B(n11430), .Y(n11473) );
  NAND2X1 U4151 ( .A(n573), .B(n10554), .Y(n10597) );
  NAND2X1 U4152 ( .A(n574), .B(n9678), .Y(n9721) );
  NAND2X1 U4153 ( .A(n575), .B(n8802), .Y(n8845) );
  NAND2X1 U4154 ( .A(n576), .B(n7926), .Y(n7969) );
  NAND2X1 U4155 ( .A(n513), .B(n993), .Y(n9949) );
  NAND2X1 U4156 ( .A(n514), .B(n1135), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n134) );
  NAND2X1 U4157 ( .A(n515), .B(n937), .Y(n11117) );
  NAND2X1 U4158 ( .A(n516), .B(n1077), .Y(n8197) );
  NAND2X1 U4159 ( .A(n522), .B(n951), .Y(n10825) );
  NAND2X1 U4160 ( .A(n524), .B(n1035), .Y(n9073) );
  NAND2X1 U4161 ( .A(n526), .B(n1119), .Y(n7321) );
  NAND2X1 U4162 ( .A(n528), .B(n979), .Y(n10241) );
  NAND2X1 U4163 ( .A(n521), .B(n1021), .Y(n9365) );
  NAND2X1 U4164 ( .A(n517), .B(n1063), .Y(n8489) );
  NAND2X1 U4165 ( .A(n523), .B(n1105), .Y(n7613) );
  NAND2X1 U4166 ( .A(n518), .B(n923), .Y(n11409) );
  NAND2X1 U4167 ( .A(n525), .B(n965), .Y(n10533) );
  NAND2X1 U4168 ( .A(n519), .B(n1007), .Y(n9657) );
  NAND2X1 U4169 ( .A(n527), .B(n1049), .Y(n8781) );
  NAND2X1 U4170 ( .A(n520), .B(n1091), .Y(n7905) );
  NAND2X1 U4171 ( .A(n1136), .B(n3482), .Y(n13876) );
  NAND2X1 U4172 ( .A(n997), .B(n2881), .Y(n17026) );
  NAND2X1 U4173 ( .A(n941), .B(n2639), .Y(n18286) );
  NAND2X1 U4174 ( .A(n1081), .B(n3241), .Y(n15136) );
  NAND2X1 U4175 ( .A(n1067), .B(n3180), .Y(n15451) );
  NAND2X1 U4176 ( .A(n927), .B(n2578), .Y(n18601) );
  NAND2X1 U4177 ( .A(n1011), .B(n2942), .Y(n16711) );
  NAND2X1 U4178 ( .A(n1095), .B(n3302), .Y(n14821) );
  NAND2X1 U4179 ( .A(n1025), .B(n3003), .Y(n16396) );
  NAND2X1 U4180 ( .A(n955), .B(n2700), .Y(n17971) );
  NAND2X1 U4181 ( .A(n1109), .B(n3363), .Y(n14506) );
  NAND2X1 U4182 ( .A(n1039), .B(n3061), .Y(n16081) );
  NAND2X1 U4183 ( .A(n969), .B(n2760), .Y(n17656) );
  NAND2X1 U4184 ( .A(n1123), .B(n3421), .Y(n14191) );
  NAND2X1 U4185 ( .A(n1053), .B(n3122), .Y(n15766) );
  NAND2X1 U4186 ( .A(n983), .B(n2821), .Y(n17341) );
  NAND2X1 U4187 ( .A(n5336), .B(n353), .Y(n9999) );
  NAND2X1 U4188 ( .A(n6132), .B(n354), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n185) );
  NAND2X1 U4189 ( .A(n4982), .B(n356), .Y(n11167) );
  NAND2X1 U4190 ( .A(n5808), .B(n355), .Y(n8247) );
  NAND2X1 U4191 ( .A(n5066), .B(n357), .Y(n10875) );
  NAND2X1 U4192 ( .A(n6036), .B(n358), .Y(n7371) );
  NAND2X1 U4193 ( .A(n5572), .B(n359), .Y(n9123) );
  NAND2X1 U4194 ( .A(n5252), .B(n360), .Y(n10291) );
  NAND2X1 U4195 ( .A(n5496), .B(n361), .Y(n9415) );
  NAND2X1 U4196 ( .A(n5724), .B(n362), .Y(n8539) );
  NAND2X1 U4197 ( .A(n5960), .B(n363), .Y(n7663) );
  NAND2X1 U4198 ( .A(n4866), .B(n364), .Y(n11459) );
  NAND2X1 U4199 ( .A(n5174), .B(n365), .Y(n10583) );
  NAND2X1 U4200 ( .A(n5420), .B(n366), .Y(n9707) );
  NAND2X1 U4201 ( .A(n5648), .B(n367), .Y(n8831) );
  NAND2X1 U4202 ( .A(n5884), .B(n368), .Y(n7955) );
  CLKINVX3 U4203 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n78), .Y(n6119) );
  CLKINVX3 U4204 ( .A(n9895), .Y(n5333) );
  CLKINVX3 U4205 ( .A(n11063), .Y(n4979) );
  CLKINVX3 U4206 ( .A(n8143), .Y(n5805) );
  CLKINVX3 U4207 ( .A(n10771), .Y(n5063) );
  CLKINVX3 U4208 ( .A(n7267), .Y(n6033) );
  CLKINVX3 U4209 ( .A(n9019), .Y(n5569) );
  CLKINVX3 U4210 ( .A(n10187), .Y(n5249) );
  CLKINVX3 U4211 ( .A(n9311), .Y(n5493) );
  CLKINVX3 U4212 ( .A(n8435), .Y(n5721) );
  CLKINVX3 U4213 ( .A(n7559), .Y(n5957) );
  CLKINVX3 U4214 ( .A(n11355), .Y(n4863) );
  CLKINVX3 U4215 ( .A(n10479), .Y(n5171) );
  CLKINVX3 U4216 ( .A(n9603), .Y(n5417) );
  CLKINVX3 U4217 ( .A(n8727), .Y(n5645) );
  CLKINVX3 U4218 ( .A(n7851), .Y(n5881) );
  CLKINVX3 U4219 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n101), .Y(n6166) );
  CLKINVX3 U4220 ( .A(n9917), .Y(n5376) );
  CLKINVX3 U4221 ( .A(n8165), .Y(n5848) );
  CLKINVX3 U4222 ( .A(n11085), .Y(n5022) );
  CLKINVX3 U4223 ( .A(n10793), .Y(n5106) );
  CLKINVX3 U4224 ( .A(n7289), .Y(n6076) );
  CLKINVX3 U4225 ( .A(n9041), .Y(n5612) );
  CLKINVX3 U4226 ( .A(n10209), .Y(n5292) );
  CLKINVX3 U4227 ( .A(n9333), .Y(n5536) );
  CLKINVX3 U4228 ( .A(n8457), .Y(n5764) );
  CLKINVX3 U4229 ( .A(n7581), .Y(n6000) );
  CLKINVX3 U4230 ( .A(n11377), .Y(n4906) );
  CLKINVX3 U4231 ( .A(n10501), .Y(n5214) );
  CLKINVX3 U4232 ( .A(n9625), .Y(n5460) );
  CLKINVX3 U4233 ( .A(n8749), .Y(n5688) );
  CLKINVX3 U4234 ( .A(n7873), .Y(n5924) );
  AOI21XL U4235 ( .A0(n9900), .A1(n546), .B0(n9986), .Y(n10062) );
  AOI21XL U4236 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .A1(n545), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n172), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n248) );
  AOI21XL U4237 ( .A0(n11068), .A1(n547), .B0(n11154), .Y(n11230) );
  AOI21XL U4238 ( .A0(n8148), .A1(n548), .B0(n8234), .Y(n8310) );
  AOI21XL U4239 ( .A0(n10776), .A1(n549), .B0(n10862), .Y(n10938) );
  AOI21XL U4240 ( .A0(n7272), .A1(n551), .B0(n7358), .Y(n7434) );
  AOI21XL U4241 ( .A0(n9024), .A1(n550), .B0(n9110), .Y(n9186) );
  AOI21XL U4242 ( .A0(n10192), .A1(n552), .B0(n10278), .Y(n10354) );
  AOI21XL U4243 ( .A0(n9316), .A1(n553), .B0(n9402), .Y(n9478) );
  AOI21XL U4244 ( .A0(n8440), .A1(n554), .B0(n8526), .Y(n8602) );
  AOI21XL U4245 ( .A0(n7564), .A1(n555), .B0(n7650), .Y(n7726) );
  AOI21XL U4246 ( .A0(n11360), .A1(n556), .B0(n11446), .Y(n11522) );
  AOI21XL U4247 ( .A0(n10484), .A1(n557), .B0(n10570), .Y(n10646) );
  AOI21XL U4248 ( .A0(n9608), .A1(n558), .B0(n9694), .Y(n9770) );
  AOI21XL U4249 ( .A0(n8732), .A1(n559), .B0(n8818), .Y(n8894) );
  AOI21XL U4250 ( .A0(n7856), .A1(n560), .B0(n7942), .Y(n8018) );
  NAND2X1 U4251 ( .A(n546), .B(n2893), .Y(n9957) );
  NAND2X1 U4252 ( .A(n545), .B(n3494), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n142) );
  NAND2X1 U4253 ( .A(n547), .B(n2650), .Y(n11125) );
  NAND2X1 U4254 ( .A(n548), .B(n3253), .Y(n8205) );
  NAND2X1 U4255 ( .A(n549), .B(n2711), .Y(n10833) );
  NAND2X1 U4256 ( .A(n550), .B(n3072), .Y(n9081) );
  NAND2X1 U4257 ( .A(n551), .B(n3433), .Y(n7329) );
  NAND2X1 U4258 ( .A(n552), .B(n2833), .Y(n10249) );
  NAND2X1 U4259 ( .A(n553), .B(n3015), .Y(n9373) );
  NAND2X1 U4260 ( .A(n554), .B(n3192), .Y(n8497) );
  NAND2X1 U4261 ( .A(n555), .B(n3375), .Y(n7621) );
  NAND2X1 U4262 ( .A(n556), .B(top_core_EC_ss_in[120]), .Y(n11417) );
  NAND2X1 U4263 ( .A(n557), .B(n2772), .Y(n10541) );
  NAND2X1 U4264 ( .A(n558), .B(n2954), .Y(n9665) );
  NAND2X1 U4265 ( .A(n559), .B(n3134), .Y(n8789) );
  NAND2X1 U4266 ( .A(n560), .B(n3314), .Y(n7913) );
  NAND2X1 U4267 ( .A(n5362), .B(n1309), .Y(n17113) );
  NAND2X1 U4268 ( .A(n6130), .B(n1279), .Y(n13963) );
  NAND2X1 U4269 ( .A(n5008), .B(n1321), .Y(n18373) );
  NAND2X1 U4270 ( .A(n5834), .B(n1291), .Y(n15223) );
  NAND2X1 U4271 ( .A(n5750), .B(n1294), .Y(n15538) );
  NAND2X1 U4272 ( .A(n4892), .B(n1324), .Y(n18688) );
  NAND2X1 U4273 ( .A(n5446), .B(n1306), .Y(n16798) );
  NAND2X1 U4274 ( .A(n5910), .B(n1288), .Y(n14908) );
  NAND2X1 U4275 ( .A(n5522), .B(n1303), .Y(n16483) );
  NAND2X1 U4276 ( .A(n5092), .B(n1318), .Y(n18058) );
  NAND2X1 U4277 ( .A(n5986), .B(n1285), .Y(n14593) );
  NAND2X1 U4278 ( .A(n5598), .B(n1300), .Y(n16168) );
  NAND2X1 U4279 ( .A(n5200), .B(n1315), .Y(n17743) );
  NAND2X1 U4280 ( .A(n6062), .B(n1282), .Y(n14278) );
  NAND2X1 U4281 ( .A(n5674), .B(n1297), .Y(n15853) );
  NAND2X1 U4282 ( .A(n5278), .B(n1312), .Y(n17428) );
  NAND2X1 U4283 ( .A(n481), .B(n546), .Y(n9947) );
  NAND2X1 U4284 ( .A(n482), .B(n545), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n132) );
  NAND2X1 U4285 ( .A(n483), .B(n547), .Y(n11115) );
  NAND2X1 U4286 ( .A(n484), .B(n548), .Y(n8195) );
  NAND2X1 U4287 ( .A(n485), .B(n549), .Y(n10823) );
  NAND2X1 U4288 ( .A(n487), .B(n551), .Y(n7319) );
  NAND2X1 U4289 ( .A(n486), .B(n550), .Y(n9071) );
  NAND2X1 U4290 ( .A(n488), .B(n552), .Y(n10239) );
  NAND2X1 U4291 ( .A(n489), .B(n553), .Y(n9363) );
  NAND2X1 U4292 ( .A(n490), .B(n554), .Y(n8487) );
  NAND2X1 U4293 ( .A(n491), .B(n555), .Y(n7611) );
  NAND2X1 U4294 ( .A(n492), .B(n556), .Y(n11407) );
  NAND2X1 U4295 ( .A(n493), .B(n557), .Y(n10531) );
  NAND2X1 U4296 ( .A(n494), .B(n558), .Y(n9655) );
  NAND2X1 U4297 ( .A(n495), .B(n559), .Y(n8779) );
  NAND2X1 U4298 ( .A(n496), .B(n560), .Y(n7903) );
  NAND2X1 U4299 ( .A(n562), .B(n353), .Y(n9930) );
  NAND2X1 U4300 ( .A(n561), .B(n354), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n115) );
  NAND2X1 U4301 ( .A(n563), .B(n356), .Y(n11098) );
  NAND2X1 U4302 ( .A(n564), .B(n355), .Y(n8178) );
  NAND2X1 U4303 ( .A(n565), .B(n357), .Y(n10806) );
  NAND2X1 U4304 ( .A(n566), .B(n359), .Y(n9054) );
  NAND2X1 U4305 ( .A(n567), .B(n358), .Y(n7302) );
  NAND2X1 U4306 ( .A(n568), .B(n360), .Y(n10222) );
  NAND2X1 U4307 ( .A(n569), .B(n361), .Y(n9346) );
  NAND2X1 U4308 ( .A(n570), .B(n362), .Y(n8470) );
  NAND2X1 U4309 ( .A(n571), .B(n363), .Y(n7594) );
  NAND2X1 U4310 ( .A(n572), .B(n364), .Y(n11390) );
  NAND2X1 U4311 ( .A(n573), .B(n365), .Y(n10514) );
  NAND2X1 U4312 ( .A(n574), .B(n366), .Y(n9638) );
  NAND2X1 U4313 ( .A(n575), .B(n367), .Y(n8762) );
  NAND2X1 U4314 ( .A(n576), .B(n368), .Y(n7886) );
  NAND2X1 U4315 ( .A(n514), .B(n6130), .Y(n13979) );
  NAND2X1 U4316 ( .A(n513), .B(n5362), .Y(n17129) );
  NAND2X1 U4317 ( .A(n515), .B(n5008), .Y(n18389) );
  NAND2X1 U4318 ( .A(n516), .B(n5834), .Y(n15239) );
  NAND2X1 U4319 ( .A(n517), .B(n5750), .Y(n15554) );
  NAND2X1 U4320 ( .A(n518), .B(n4892), .Y(n18704) );
  NAND2X1 U4321 ( .A(n519), .B(n5446), .Y(n16814) );
  NAND2X1 U4322 ( .A(n520), .B(n5910), .Y(n14924) );
  NAND2X1 U4323 ( .A(n521), .B(n5522), .Y(n16499) );
  NAND2X1 U4324 ( .A(n522), .B(n5092), .Y(n18074) );
  NAND2X1 U4325 ( .A(n523), .B(n5986), .Y(n14609) );
  NAND2X1 U4326 ( .A(n524), .B(n5598), .Y(n16184) );
  NAND2X1 U4327 ( .A(n525), .B(n5200), .Y(n17759) );
  NAND2X1 U4328 ( .A(n526), .B(n6062), .Y(n14294) );
  NAND2X1 U4329 ( .A(n527), .B(n5674), .Y(n15869) );
  NAND2X1 U4330 ( .A(n528), .B(n5278), .Y(n17444) );
  AOI21XL U4331 ( .A0(n2871), .A1(n9891), .B0(n417), .Y(n9945) );
  AOI21XL U4332 ( .A0(n3472), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), 
        .B0(n418), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n130) );
  AOI21XL U4333 ( .A0(n2629), .A1(n11059), .B0(n419), .Y(n11113) );
  AOI21XL U4334 ( .A0(n3231), .A1(n8139), .B0(n420), .Y(n8193) );
  AOI21XL U4335 ( .A0(n2690), .A1(n10767), .B0(n421), .Y(n10821) );
  AOI21XL U4336 ( .A0(n3051), .A1(n9015), .B0(n422), .Y(n9069) );
  AOI21XL U4337 ( .A0(n3411), .A1(n7263), .B0(n423), .Y(n7317) );
  AOI21XL U4338 ( .A0(n2811), .A1(n10183), .B0(n424), .Y(n10237) );
  AOI21XL U4339 ( .A0(n2993), .A1(n9307), .B0(n425), .Y(n9361) );
  AOI21XL U4340 ( .A0(n3170), .A1(n8431), .B0(n426), .Y(n8485) );
  AOI21XL U4341 ( .A0(n3353), .A1(n7555), .B0(n427), .Y(n7609) );
  AOI21XL U4342 ( .A0(n2568), .A1(n11351), .B0(n428), .Y(n11405) );
  AOI21XL U4343 ( .A0(n2750), .A1(n10475), .B0(n429), .Y(n10529) );
  AOI21XL U4344 ( .A0(n2932), .A1(n9599), .B0(n430), .Y(n9653) );
  AOI21XL U4345 ( .A0(n3112), .A1(n8723), .B0(n431), .Y(n8777) );
  AOI21XL U4346 ( .A0(n3292), .A1(n7847), .B0(n432), .Y(n7901) );
  NAND2X1 U4347 ( .A(n1141), .B(n6130), .Y(n13877) );
  NAND2X1 U4348 ( .A(n1002), .B(n5362), .Y(n17027) );
  NAND2X1 U4349 ( .A(n946), .B(n5008), .Y(n18287) );
  NAND2X1 U4350 ( .A(n1086), .B(n5834), .Y(n15137) );
  NAND2X1 U4351 ( .A(n1072), .B(n5750), .Y(n15452) );
  NAND2X1 U4352 ( .A(n932), .B(n4892), .Y(n18602) );
  NAND2X1 U4353 ( .A(n1016), .B(n5446), .Y(n16712) );
  NAND2X1 U4354 ( .A(n1100), .B(n5910), .Y(n14822) );
  NAND2X1 U4355 ( .A(n1030), .B(n5522), .Y(n16397) );
  NAND2X1 U4356 ( .A(n960), .B(n5092), .Y(n17972) );
  NAND2X1 U4357 ( .A(n1114), .B(n5986), .Y(n14507) );
  NAND2X1 U4358 ( .A(n1044), .B(n5598), .Y(n16082) );
  NAND2X1 U4359 ( .A(n974), .B(n5200), .Y(n17657) );
  NAND2X1 U4360 ( .A(n1128), .B(n6062), .Y(n14192) );
  NAND2X1 U4361 ( .A(n1058), .B(n5674), .Y(n15767) );
  NAND2X1 U4362 ( .A(n988), .B(n5278), .Y(n17342) );
  NOR2X1 U4363 ( .A(n17065), .B(n401), .Y(n17092) );
  NOR2X1 U4364 ( .A(n13915), .B(n402), .Y(n13942) );
  NOR2X1 U4365 ( .A(n18325), .B(n403), .Y(n18352) );
  NOR2X1 U4366 ( .A(n15175), .B(n404), .Y(n15202) );
  NOR2X1 U4367 ( .A(n15490), .B(n410), .Y(n15517) );
  NOR2X1 U4368 ( .A(n18640), .B(n412), .Y(n18667) );
  NOR2X1 U4369 ( .A(n16750), .B(n414), .Y(n16777) );
  NOR2X1 U4370 ( .A(n14860), .B(n416), .Y(n14887) );
  NOR2X1 U4371 ( .A(n16435), .B(n409), .Y(n16462) );
  NOR2X1 U4372 ( .A(n18010), .B(n405), .Y(n18037) );
  NOR2X1 U4373 ( .A(n14545), .B(n411), .Y(n14572) );
  NOR2X1 U4374 ( .A(n16120), .B(n406), .Y(n16147) );
  NOR2X1 U4375 ( .A(n17695), .B(n413), .Y(n17722) );
  NOR2X1 U4376 ( .A(n14230), .B(n407), .Y(n14257) );
  NOR2X1 U4377 ( .A(n15805), .B(n415), .Y(n15832) );
  NOR2X1 U4378 ( .A(n17380), .B(n408), .Y(n17407) );
  AOI31X1 U4379 ( .A0(n13964), .A1(n14014), .A2(n13877), .B0(n3454), .Y(n14102) );
  AOI31X1 U4380 ( .A0(n17114), .A1(n17164), .A2(n17027), .B0(n2853), .Y(n17252) );
  AOI31X1 U4381 ( .A0(n18374), .A1(n18424), .A2(n18287), .B0(n2611), .Y(n18512) );
  AOI31X1 U4382 ( .A0(n15224), .A1(n15274), .A2(n15137), .B0(n3213), .Y(n15362) );
  AOI31X1 U4383 ( .A0(n15539), .A1(n15589), .A2(n15452), .B0(n3152), .Y(n15677) );
  AOI31X1 U4384 ( .A0(n18689), .A1(n18739), .A2(n18602), .B0(n2550), .Y(n18827) );
  AOI31X1 U4385 ( .A0(n16799), .A1(n16849), .A2(n16712), .B0(n2914), .Y(n16937) );
  AOI31X1 U4386 ( .A0(n14909), .A1(n14959), .A2(n14822), .B0(n3274), .Y(n15047) );
  AOI31X1 U4387 ( .A0(n16484), .A1(n16534), .A2(n16397), .B0(n2975), .Y(n16622) );
  AOI31X1 U4388 ( .A0(n18059), .A1(n18109), .A2(n17972), .B0(n2672), .Y(n18197) );
  AOI31X1 U4389 ( .A0(n14594), .A1(n14644), .A2(n14507), .B0(n3335), .Y(n14732) );
  AOI31X1 U4390 ( .A0(n16169), .A1(n16219), .A2(n16082), .B0(n3033), .Y(n16307) );
  AOI31X1 U4391 ( .A0(n17744), .A1(n17794), .A2(n17657), .B0(n2732), .Y(n17882) );
  AOI31X1 U4392 ( .A0(n14279), .A1(n14329), .A2(n14192), .B0(n3393), .Y(n14417) );
  AOI31X1 U4393 ( .A0(n15854), .A1(n15904), .A2(n15767), .B0(n3094), .Y(n15992) );
  AOI31X1 U4394 ( .A0(n17429), .A1(n17479), .A2(n17342), .B0(n2793), .Y(n17567) );
  INVX1 U4395 ( .A(n17035), .Y(n5335) );
  INVX1 U4396 ( .A(n13885), .Y(n6118) );
  INVX1 U4397 ( .A(n18295), .Y(n4981) );
  INVX1 U4398 ( .A(n15145), .Y(n5807) );
  INVX1 U4399 ( .A(n15460), .Y(n5723) );
  INVX1 U4400 ( .A(n18610), .Y(n4865) );
  INVX1 U4401 ( .A(n16720), .Y(n5419) );
  INVX1 U4402 ( .A(n14830), .Y(n5883) );
  INVX1 U4403 ( .A(n16405), .Y(n5495) );
  INVX1 U4404 ( .A(n17980), .Y(n5065) );
  INVX1 U4405 ( .A(n14515), .Y(n5959) );
  INVX1 U4406 ( .A(n16090), .Y(n5571) );
  INVX1 U4407 ( .A(n17665), .Y(n5173) );
  INVX1 U4408 ( .A(n14200), .Y(n6035) );
  INVX1 U4409 ( .A(n15775), .Y(n5647) );
  INVX1 U4410 ( .A(n17350), .Y(n5251) );
  NOR2X1 U4411 ( .A(n305), .B(n433), .Y(n17285) );
  XNOR2X1 U4412 ( .A(n2871), .B(n2892), .Y(n305) );
  NOR2X1 U4413 ( .A(n306), .B(n434), .Y(n14135) );
  XNOR2X1 U4414 ( .A(n3472), .B(n3493), .Y(n306) );
  NOR2X1 U4415 ( .A(n307), .B(n436), .Y(n15395) );
  XNOR2X1 U4416 ( .A(n3231), .B(n3252), .Y(n307) );
  NOR2X1 U4417 ( .A(n308), .B(n435), .Y(n18545) );
  XNOR2X1 U4418 ( .A(n2629), .B(n2661), .Y(n308) );
  NOR2X1 U4419 ( .A(n309), .B(n437), .Y(n15710) );
  XNOR2X1 U4420 ( .A(n3170), .B(n3191), .Y(n309) );
  NOR2X1 U4421 ( .A(n310), .B(n438), .Y(n16970) );
  XNOR2X1 U4422 ( .A(n2932), .B(n2953), .Y(n310) );
  NOR2X1 U4423 ( .A(n311), .B(n439), .Y(n18860) );
  XNOR2X1 U4424 ( .A(n2568), .B(n2589), .Y(n311) );
  NOR2X1 U4425 ( .A(n312), .B(n440), .Y(n15080) );
  XNOR2X1 U4426 ( .A(n3292), .B(n3313), .Y(n312) );
  NOR2X1 U4427 ( .A(n313), .B(n441), .Y(n16655) );
  XNOR2X1 U4428 ( .A(n2993), .B(n3014), .Y(n313) );
  NOR2X1 U4429 ( .A(n314), .B(n442), .Y(n18230) );
  XNOR2X1 U4430 ( .A(n2690), .B(n2710), .Y(n314) );
  NOR2X1 U4431 ( .A(n315), .B(n443), .Y(n14765) );
  XNOR2X1 U4432 ( .A(n3353), .B(n3374), .Y(n315) );
  NOR2X1 U4433 ( .A(n316), .B(n444), .Y(n16340) );
  XNOR2X1 U4434 ( .A(n3051), .B(n3083), .Y(n316) );
  NOR2X1 U4435 ( .A(n317), .B(n445), .Y(n17915) );
  XNOR2X1 U4436 ( .A(n2750), .B(n2771), .Y(n317) );
  NOR2X1 U4437 ( .A(n318), .B(n446), .Y(n14450) );
  XNOR2X1 U4438 ( .A(n3411), .B(n3432), .Y(n318) );
  NOR2X1 U4439 ( .A(n319), .B(n447), .Y(n16025) );
  XNOR2X1 U4440 ( .A(n3112), .B(n3133), .Y(n319) );
  NOR2X1 U4441 ( .A(n320), .B(n448), .Y(n17600) );
  XNOR2X1 U4442 ( .A(n2811), .B(n2832), .Y(n320) );
  NAND2X1 U4443 ( .A(n5362), .B(n1003), .Y(n17082) );
  NAND2X1 U4444 ( .A(n6130), .B(n1142), .Y(n13932) );
  NAND2X1 U4445 ( .A(n5008), .B(n947), .Y(n18342) );
  NAND2X1 U4446 ( .A(n5834), .B(n1087), .Y(n15192) );
  NAND2X1 U4447 ( .A(n5750), .B(n1073), .Y(n15507) );
  NAND2X1 U4448 ( .A(n5446), .B(n1017), .Y(n16767) );
  NAND2X1 U4449 ( .A(n4892), .B(n933), .Y(n18657) );
  NAND2X1 U4450 ( .A(n5910), .B(n1101), .Y(n14877) );
  NAND2X1 U4451 ( .A(n5522), .B(n1031), .Y(n16452) );
  NAND2X1 U4452 ( .A(n5092), .B(n961), .Y(n18027) );
  NAND2X1 U4453 ( .A(n5986), .B(n1115), .Y(n14562) );
  NAND2X1 U4454 ( .A(n5598), .B(n1045), .Y(n16137) );
  NAND2X1 U4455 ( .A(n5200), .B(n975), .Y(n17712) );
  NAND2X1 U4456 ( .A(n6062), .B(n1129), .Y(n14247) );
  NAND2X1 U4457 ( .A(n5674), .B(n1059), .Y(n15822) );
  NAND2X1 U4458 ( .A(n5278), .B(n989), .Y(n17397) );
  NAND2X1 U4459 ( .A(n5376), .B(n2893), .Y(n17081) );
  NAND2X1 U4460 ( .A(n6166), .B(n3494), .Y(n13931) );
  NAND2X1 U4461 ( .A(n5022), .B(n2650), .Y(n18341) );
  NAND2X1 U4462 ( .A(n5848), .B(n3253), .Y(n15191) );
  NAND2X1 U4463 ( .A(n5764), .B(n3192), .Y(n15506) );
  NAND2X1 U4464 ( .A(n5460), .B(n2954), .Y(n16766) );
  NAND2X1 U4465 ( .A(n4906), .B(n2599), .Y(n18656) );
  NAND2X1 U4466 ( .A(n5924), .B(n3314), .Y(n14876) );
  NAND2X1 U4467 ( .A(n5536), .B(n3015), .Y(n16451) );
  NAND2X1 U4468 ( .A(n5106), .B(n2711), .Y(n18026) );
  NAND2X1 U4469 ( .A(n6000), .B(n3375), .Y(n14561) );
  NAND2X1 U4470 ( .A(n5612), .B(n3072), .Y(n16136) );
  NAND2X1 U4471 ( .A(n5214), .B(n2772), .Y(n17711) );
  NAND2X1 U4472 ( .A(n6076), .B(n3433), .Y(n14246) );
  NAND2X1 U4473 ( .A(n5688), .B(n3134), .Y(n15821) );
  NAND2X1 U4474 ( .A(n5292), .B(n2833), .Y(n17396) );
  INVX1 U4475 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n108), .Y(n6155) );
  INVX1 U4476 ( .A(n9923), .Y(n5365) );
  INVX1 U4477 ( .A(n11091), .Y(n5011) );
  INVX1 U4478 ( .A(n8171), .Y(n5837) );
  INVX1 U4479 ( .A(n10799), .Y(n5095) );
  INVX1 U4480 ( .A(n9047), .Y(n5601) );
  INVX1 U4481 ( .A(n7295), .Y(n6065) );
  INVX1 U4482 ( .A(n10215), .Y(n5281) );
  INVX1 U4483 ( .A(n9339), .Y(n5525) );
  INVX1 U4484 ( .A(n8463), .Y(n5753) );
  INVX1 U4485 ( .A(n7587), .Y(n5989) );
  INVX1 U4486 ( .A(n11383), .Y(n4895) );
  INVX1 U4487 ( .A(n10507), .Y(n5203) );
  INVX1 U4488 ( .A(n9631), .Y(n5449) );
  INVX1 U4489 ( .A(n8755), .Y(n5677) );
  INVX1 U4490 ( .A(n7879), .Y(n5913) );
  OAI21XL U4491 ( .A0(n5376), .A1(n546), .B0(n9913), .Y(n10152) );
  OAI21XL U4492 ( .A0(n6166), .A1(n545), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n338) );
  OAI21XL U4493 ( .A0(n5848), .A1(n548), .B0(n8161), .Y(n8400) );
  OAI21XL U4494 ( .A0(n5022), .A1(n547), .B0(n11081), .Y(n11320) );
  OAI21XL U4495 ( .A0(n5106), .A1(n549), .B0(n10789), .Y(n11028) );
  OAI21XL U4496 ( .A0(n6076), .A1(n551), .B0(n7285), .Y(n7524) );
  OAI21XL U4497 ( .A0(n5612), .A1(n550), .B0(n9037), .Y(n9276) );
  OAI21XL U4498 ( .A0(n5292), .A1(n552), .B0(n10205), .Y(n10444) );
  OAI21XL U4499 ( .A0(n5536), .A1(n553), .B0(n9329), .Y(n9568) );
  OAI21XL U4500 ( .A0(n5764), .A1(n554), .B0(n8453), .Y(n8692) );
  OAI21XL U4501 ( .A0(n6000), .A1(n555), .B0(n7577), .Y(n7816) );
  OAI21XL U4502 ( .A0(n4906), .A1(n556), .B0(n11373), .Y(n11612) );
  OAI21XL U4503 ( .A0(n5214), .A1(n557), .B0(n10497), .Y(n10736) );
  OAI21XL U4504 ( .A0(n5460), .A1(n558), .B0(n9621), .Y(n9860) );
  OAI21XL U4505 ( .A0(n5688), .A1(n559), .B0(n8745), .Y(n8984) );
  OAI21XL U4506 ( .A0(n5924), .A1(n560), .B0(n7869), .Y(n8108) );
  INVX1 U4507 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n197), .Y(n6135) );
  INVX1 U4508 ( .A(n10011), .Y(n5339) );
  INVX1 U4509 ( .A(n11179), .Y(n4985) );
  INVX1 U4510 ( .A(n8259), .Y(n5811) );
  INVX1 U4511 ( .A(n10887), .Y(n5069) );
  INVX1 U4512 ( .A(n9135), .Y(n5575) );
  INVX1 U4513 ( .A(n7383), .Y(n6039) );
  INVX1 U4514 ( .A(n10303), .Y(n5255) );
  INVX1 U4515 ( .A(n9427), .Y(n5499) );
  INVX1 U4516 ( .A(n8551), .Y(n5727) );
  INVX1 U4517 ( .A(n7675), .Y(n5963) );
  INVX1 U4518 ( .A(n11471), .Y(n4869) );
  INVX1 U4519 ( .A(n10595), .Y(n5177) );
  INVX1 U4520 ( .A(n9719), .Y(n5423) );
  INVX1 U4521 ( .A(n8843), .Y(n5651) );
  INVX1 U4522 ( .A(n7967), .Y(n5887) );
  NOR2XL U4523 ( .A(n10035), .B(n5365), .Y(n10053) );
  NOR2XL U4524 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n221), .B(n6155), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n239) );
  NOR2XL U4525 ( .A(n11203), .B(n5011), .Y(n11221) );
  NOR2XL U4526 ( .A(n8283), .B(n5837), .Y(n8301) );
  NOR2XL U4527 ( .A(n10911), .B(n5095), .Y(n10929) );
  NOR2XL U4528 ( .A(n9159), .B(n5601), .Y(n9177) );
  NOR2XL U4529 ( .A(n7407), .B(n6065), .Y(n7425) );
  NOR2XL U4530 ( .A(n10327), .B(n5281), .Y(n10345) );
  NOR2XL U4531 ( .A(n9451), .B(n5525), .Y(n9469) );
  NOR2XL U4532 ( .A(n8575), .B(n5753), .Y(n8593) );
  NOR2XL U4533 ( .A(n7699), .B(n5989), .Y(n7717) );
  NOR2XL U4534 ( .A(n11495), .B(n4895), .Y(n11513) );
  NOR2XL U4535 ( .A(n10619), .B(n5203), .Y(n10637) );
  NOR2XL U4536 ( .A(n9743), .B(n5449), .Y(n9761) );
  NOR2XL U4537 ( .A(n8867), .B(n5677), .Y(n8885) );
  NOR2XL U4538 ( .A(n7991), .B(n5913), .Y(n8009) );
  INVX1 U4539 ( .A(n9912), .Y(n5371) );
  INVX1 U4540 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n96), .Y(n6161) );
  INVX1 U4541 ( .A(n8160), .Y(n5843) );
  INVX1 U4542 ( .A(n11080), .Y(n5017) );
  INVX1 U4543 ( .A(n10788), .Y(n5101) );
  INVX1 U4544 ( .A(n7284), .Y(n6071) );
  INVX1 U4545 ( .A(n9036), .Y(n5607) );
  INVX1 U4546 ( .A(n10204), .Y(n5287) );
  INVX1 U4547 ( .A(n9328), .Y(n5531) );
  INVX1 U4548 ( .A(n8452), .Y(n5759) );
  INVX1 U4549 ( .A(n7576), .Y(n5995) );
  INVX1 U4550 ( .A(n11372), .Y(n4901) );
  INVX1 U4551 ( .A(n10496), .Y(n5209) );
  INVX1 U4552 ( .A(n9620), .Y(n5455) );
  INVX1 U4553 ( .A(n8744), .Y(n5683) );
  INVX1 U4554 ( .A(n7868), .Y(n5919) );
  AND2X2 U4555 ( .A(n2880), .B(n2893), .Y(n353) );
  AND2X2 U4556 ( .A(n3481), .B(n3494), .Y(n354) );
  AND2X2 U4557 ( .A(n3240), .B(n3253), .Y(n355) );
  AND2X2 U4558 ( .A(n2638), .B(n2650), .Y(n356) );
  AND2X2 U4559 ( .A(n2699), .B(n2711), .Y(n357) );
  AND2X2 U4560 ( .A(n3420), .B(n3433), .Y(n358) );
  AND2X2 U4561 ( .A(n3060), .B(n3072), .Y(n359) );
  AND2X2 U4562 ( .A(n2820), .B(n2833), .Y(n360) );
  AND2X2 U4563 ( .A(n3002), .B(n3015), .Y(n361) );
  AND2X2 U4564 ( .A(n3179), .B(n3192), .Y(n362) );
  AND2X2 U4565 ( .A(n3362), .B(n3375), .Y(n363) );
  AND2X2 U4566 ( .A(n2577), .B(n2590), .Y(n364) );
  AND2X2 U4567 ( .A(n2759), .B(n2772), .Y(n365) );
  AND2X2 U4568 ( .A(n2941), .B(n2954), .Y(n366) );
  AND2X2 U4569 ( .A(n3121), .B(n3134), .Y(n367) );
  AND2X2 U4570 ( .A(n3301), .B(n3314), .Y(n368) );
  OAI21XL U4571 ( .A0(n338), .A1(n14073), .B0(n14108), .Y(n14107) );
  OAI21XL U4572 ( .A0(n6149), .A1(n6130), .B0(n3494), .Y(n14108) );
  OAI21XL U4573 ( .A0(n337), .A1(n17223), .B0(n17258), .Y(n17257) );
  OAI21XL U4574 ( .A0(n5378), .A1(n5362), .B0(n2893), .Y(n17258) );
  OAI21XL U4575 ( .A0(n339), .A1(n18483), .B0(n18518), .Y(n18517) );
  OAI21XL U4576 ( .A0(n5024), .A1(n5008), .B0(n2650), .Y(n18518) );
  OAI21XL U4577 ( .A0(n340), .A1(n15333), .B0(n15368), .Y(n15367) );
  OAI21XL U4578 ( .A0(n5850), .A1(n5834), .B0(n3253), .Y(n15368) );
  OAI21XL U4579 ( .A0(n341), .A1(n15648), .B0(n15683), .Y(n15682) );
  OAI21XL U4580 ( .A0(n5766), .A1(n5750), .B0(n3192), .Y(n15683) );
  OAI21XL U4581 ( .A0(n343), .A1(n18798), .B0(n18833), .Y(n18832) );
  OAI21XL U4582 ( .A0(n4908), .A1(n4892), .B0(n2590), .Y(n18833) );
  OAI21XL U4583 ( .A0(n342), .A1(n16908), .B0(n16943), .Y(n16942) );
  OAI21XL U4584 ( .A0(n5462), .A1(n5446), .B0(n2954), .Y(n16943) );
  OAI21XL U4585 ( .A0(n344), .A1(n15018), .B0(n15053), .Y(n15052) );
  OAI21XL U4586 ( .A0(n5926), .A1(n5910), .B0(n3314), .Y(n15053) );
  OAI21XL U4587 ( .A0(n345), .A1(n16593), .B0(n16628), .Y(n16627) );
  OAI21XL U4588 ( .A0(n5538), .A1(n5522), .B0(n3015), .Y(n16628) );
  OAI21XL U4589 ( .A0(n346), .A1(n18168), .B0(n18203), .Y(n18202) );
  OAI21XL U4590 ( .A0(n5108), .A1(n5092), .B0(n2711), .Y(n18203) );
  OAI21XL U4591 ( .A0(n347), .A1(n14703), .B0(n14738), .Y(n14737) );
  OAI21XL U4592 ( .A0(n6002), .A1(n5986), .B0(n3375), .Y(n14738) );
  OAI21XL U4593 ( .A0(n348), .A1(n16278), .B0(n16313), .Y(n16312) );
  OAI21XL U4594 ( .A0(n5614), .A1(n5598), .B0(n3072), .Y(n16313) );
  OAI21XL U4595 ( .A0(n349), .A1(n17853), .B0(n17888), .Y(n17887) );
  OAI21XL U4596 ( .A0(n5216), .A1(n5200), .B0(n2772), .Y(n17888) );
  OAI21XL U4597 ( .A0(n350), .A1(n14388), .B0(n14423), .Y(n14422) );
  OAI21XL U4598 ( .A0(n6078), .A1(n6062), .B0(n3433), .Y(n14423) );
  OAI21XL U4599 ( .A0(n351), .A1(n15963), .B0(n15998), .Y(n15997) );
  OAI21XL U4600 ( .A0(n5690), .A1(n5674), .B0(n3134), .Y(n15998) );
  OAI21XL U4601 ( .A0(n352), .A1(n17538), .B0(n17573), .Y(n17572) );
  OAI21XL U4602 ( .A0(n5294), .A1(n5278), .B0(n2833), .Y(n17573) );
  CLKINVX3 U4603 ( .A(n2346), .Y(n2340) );
  CLKINVX3 U4604 ( .A(n2346), .Y(n2343) );
  CLKINVX3 U4605 ( .A(n2345), .Y(n2342) );
  CLKINVX3 U4606 ( .A(n2345), .Y(n2341) );
  INVX1 U4607 ( .A(n9950), .Y(n5369) );
  INVX1 U4608 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n135), .Y(n6159) );
  INVX1 U4609 ( .A(n11118), .Y(n5015) );
  INVX1 U4610 ( .A(n8198), .Y(n5841) );
  INVX1 U4611 ( .A(n10826), .Y(n5099) );
  INVX1 U4612 ( .A(n7322), .Y(n6069) );
  INVX1 U4613 ( .A(n9074), .Y(n5605) );
  INVX1 U4614 ( .A(n10242), .Y(n5285) );
  INVX1 U4615 ( .A(n9366), .Y(n5529) );
  INVX1 U4616 ( .A(n8490), .Y(n5757) );
  INVX1 U4617 ( .A(n7614), .Y(n5993) );
  INVX1 U4618 ( .A(n11410), .Y(n4899) );
  INVX1 U4619 ( .A(n10534), .Y(n5207) );
  INVX1 U4620 ( .A(n9658), .Y(n5453) );
  INVX1 U4621 ( .A(n8782), .Y(n5681) );
  INVX1 U4622 ( .A(n7906), .Y(n5917) );
  CLKINVX3 U4623 ( .A(n238), .Y(n3629) );
  CLKINVX3 U4624 ( .A(n238), .Y(n3630) );
  CLKINVX3 U4625 ( .A(n238), .Y(n3631) );
  CLKINVX3 U4626 ( .A(n238), .Y(n3632) );
  CLKINVX3 U4627 ( .A(n238), .Y(n3633) );
  CLKINVX3 U4628 ( .A(n238), .Y(n3634) );
  CLKINVX3 U4629 ( .A(n238), .Y(n3635) );
  CLKINVX3 U4630 ( .A(n617), .Y(n3637) );
  CLKINVX3 U4631 ( .A(n617), .Y(n3638) );
  CLKINVX3 U4632 ( .A(n617), .Y(n3639) );
  CLKINVX3 U4633 ( .A(n617), .Y(n3640) );
  CLKINVX3 U4634 ( .A(n617), .Y(n3641) );
  CLKINVX3 U4635 ( .A(n617), .Y(n3642) );
  CLKINVX3 U4636 ( .A(n617), .Y(n3643) );
  CLKINVX3 U4637 ( .A(n2346), .Y(n2339) );
  CLKINVX3 U4638 ( .A(n2346), .Y(n2338) );
  CLKINVX3 U4639 ( .A(n2346), .Y(n2337) );
  INVX1 U4640 ( .A(n10065), .Y(n5340) );
  INVX1 U4641 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n251), .Y(n6136) );
  INVX1 U4642 ( .A(n8313), .Y(n5812) );
  INVX1 U4643 ( .A(n11233), .Y(n4986) );
  INVX1 U4644 ( .A(n10941), .Y(n5070) );
  INVX1 U4645 ( .A(n7437), .Y(n6040) );
  INVX1 U4646 ( .A(n9189), .Y(n5576) );
  INVX1 U4647 ( .A(n10357), .Y(n5256) );
  INVX1 U4648 ( .A(n9481), .Y(n5500) );
  INVX1 U4649 ( .A(n8605), .Y(n5728) );
  INVX1 U4650 ( .A(n7729), .Y(n5964) );
  INVX1 U4651 ( .A(n11525), .Y(n4870) );
  INVX1 U4652 ( .A(n10649), .Y(n5178) );
  INVX1 U4653 ( .A(n9773), .Y(n5424) );
  INVX1 U4654 ( .A(n8897), .Y(n5652) );
  INVX1 U4655 ( .A(n8021), .Y(n5888) );
  INVX1 U4656 ( .A(n13302), .Y(n6548) );
  INVX1 U4657 ( .A(n12672), .Y(n6843) );
  INVX1 U4658 ( .A(n12987), .Y(n6889) );
  CLKINVX3 U4659 ( .A(n3608), .Y(n3587) );
  INVX1 U4660 ( .A(n9955), .Y(n5364) );
  INVX1 U4661 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n140), .Y(n6154) );
  INVX1 U4662 ( .A(n11123), .Y(n5010) );
  INVX1 U4663 ( .A(n8203), .Y(n5836) );
  INVX1 U4664 ( .A(n10831), .Y(n5094) );
  INVX1 U4665 ( .A(n9079), .Y(n5600) );
  INVX1 U4666 ( .A(n7327), .Y(n6064) );
  INVX1 U4667 ( .A(n10247), .Y(n5280) );
  INVX1 U4668 ( .A(n9371), .Y(n5524) );
  INVX1 U4669 ( .A(n8495), .Y(n5752) );
  INVX1 U4670 ( .A(n7619), .Y(n5988) );
  INVX1 U4671 ( .A(n11415), .Y(n4894) );
  INVX1 U4672 ( .A(n10539), .Y(n5202) );
  INVX1 U4673 ( .A(n9663), .Y(n5448) );
  INVX1 U4674 ( .A(n8787), .Y(n5676) );
  INVX1 U4675 ( .A(n7911), .Y(n5912) );
  AND2X2 U4676 ( .A(n3493), .B(n3482), .Y(n369) );
  AND2X2 U4677 ( .A(n2892), .B(n2881), .Y(n370) );
  AND2X2 U4678 ( .A(n2651), .B(n2639), .Y(n371) );
  AND2X2 U4679 ( .A(n3252), .B(n3241), .Y(n372) );
  AND2X2 U4680 ( .A(n3191), .B(n3180), .Y(n373) );
  AND2X2 U4681 ( .A(n2589), .B(n2578), .Y(n374) );
  AND2X2 U4682 ( .A(n2953), .B(n2942), .Y(n375) );
  AND2X2 U4683 ( .A(n3313), .B(n3302), .Y(n376) );
  AND2X2 U4684 ( .A(n3014), .B(n3003), .Y(n377) );
  AND2X2 U4685 ( .A(n2710), .B(n2700), .Y(n378) );
  AND2X2 U4686 ( .A(n3374), .B(n3363), .Y(n379) );
  AND2X2 U4687 ( .A(n3073), .B(n3061), .Y(n380) );
  AND2X2 U4688 ( .A(n2771), .B(n2760), .Y(n381) );
  AND2X2 U4689 ( .A(n3432), .B(n3421), .Y(n382) );
  AND2X2 U4690 ( .A(n3133), .B(n3122), .Y(n383) );
  AND2X2 U4691 ( .A(n2832), .B(n2821), .Y(n384) );
  AND2X2 U4692 ( .A(n3493), .B(n3482), .Y(n385) );
  AND2X2 U4693 ( .A(n2892), .B(n2881), .Y(n386) );
  AND2X2 U4694 ( .A(n2651), .B(n2639), .Y(n387) );
  AND2X2 U4695 ( .A(n3252), .B(n3241), .Y(n388) );
  AND2X2 U4696 ( .A(n3191), .B(n3180), .Y(n389) );
  AND2X2 U4697 ( .A(n2589), .B(n2578), .Y(n390) );
  AND2X2 U4698 ( .A(n2953), .B(n2942), .Y(n391) );
  AND2X2 U4699 ( .A(n3313), .B(n3302), .Y(n392) );
  AND2X2 U4700 ( .A(n3014), .B(n3003), .Y(n393) );
  AND2X2 U4701 ( .A(n2710), .B(n2700), .Y(n394) );
  AND2X2 U4702 ( .A(n3374), .B(n3363), .Y(n395) );
  AND2X2 U4703 ( .A(n3073), .B(n3061), .Y(n396) );
  AND2X2 U4704 ( .A(n2771), .B(n2760), .Y(n397) );
  AND2X2 U4705 ( .A(n3432), .B(n3421), .Y(n398) );
  AND2X2 U4706 ( .A(n3133), .B(n3122), .Y(n399) );
  AND2X2 U4707 ( .A(n2832), .B(n2821), .Y(n400) );
  INVX1 U4708 ( .A(n17155), .Y(n5360) );
  INVX1 U4709 ( .A(n14005), .Y(n6128) );
  INVX1 U4710 ( .A(n18415), .Y(n5006) );
  INVX1 U4711 ( .A(n15265), .Y(n5832) );
  INVX1 U4712 ( .A(n15580), .Y(n5748) );
  INVX1 U4713 ( .A(n18730), .Y(n4890) );
  INVX1 U4714 ( .A(n16840), .Y(n5444) );
  INVX1 U4715 ( .A(n14950), .Y(n5908) );
  INVX1 U4716 ( .A(n16525), .Y(n5520) );
  INVX1 U4717 ( .A(n18100), .Y(n5090) );
  INVX1 U4718 ( .A(n14635), .Y(n5984) );
  INVX1 U4719 ( .A(n16210), .Y(n5596) );
  INVX1 U4720 ( .A(n17785), .Y(n5198) );
  INVX1 U4721 ( .A(n14320), .Y(n6060) );
  INVX1 U4722 ( .A(n15895), .Y(n5672) );
  INVX1 U4723 ( .A(n17470), .Y(n5276) );
  INVX1 U4724 ( .A(n10021), .Y(n5349) );
  INVX1 U4725 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n207), .Y(n6145) );
  INVX1 U4726 ( .A(n11189), .Y(n4995) );
  INVX1 U4727 ( .A(n8269), .Y(n5821) );
  INVX1 U4728 ( .A(n10897), .Y(n5079) );
  INVX1 U4729 ( .A(n9145), .Y(n5585) );
  INVX1 U4730 ( .A(n7393), .Y(n6049) );
  INVX1 U4731 ( .A(n10313), .Y(n5265) );
  INVX1 U4732 ( .A(n9437), .Y(n5509) );
  INVX1 U4733 ( .A(n8561), .Y(n5737) );
  INVX1 U4734 ( .A(n7685), .Y(n5973) );
  INVX1 U4735 ( .A(n11481), .Y(n4879) );
  INVX1 U4736 ( .A(n10605), .Y(n5187) );
  INVX1 U4737 ( .A(n9729), .Y(n5433) );
  INVX1 U4738 ( .A(n8853), .Y(n5661) );
  INVX1 U4739 ( .A(n7977), .Y(n5897) );
  INVX1 U4740 ( .A(n9904), .Y(n5343) );
  INVX1 U4741 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n87), .Y(n6139) );
  INVX1 U4742 ( .A(n8152), .Y(n5815) );
  INVX1 U4743 ( .A(n11072), .Y(n4989) );
  INVX1 U4744 ( .A(n10780), .Y(n5073) );
  INVX1 U4745 ( .A(n7276), .Y(n6043) );
  INVX1 U4746 ( .A(n9028), .Y(n5579) );
  INVX1 U4747 ( .A(n10196), .Y(n5259) );
  INVX1 U4748 ( .A(n9320), .Y(n5503) );
  INVX1 U4749 ( .A(n8444), .Y(n5731) );
  INVX1 U4750 ( .A(n7568), .Y(n5967) );
  INVX1 U4751 ( .A(n11364), .Y(n4873) );
  INVX1 U4752 ( .A(n10488), .Y(n5181) );
  INVX1 U4753 ( .A(n9612), .Y(n5427) );
  INVX1 U4754 ( .A(n8736), .Y(n5655) );
  INVX1 U4755 ( .A(n7860), .Y(n5891) );
  INVX1 U4756 ( .A(n2345), .Y(n2344) );
  INVX1 U4757 ( .A(n3615), .Y(n3606) );
  INVX1 U4758 ( .A(n3622), .Y(n3607) );
  INVX1 U4759 ( .A(n3620), .Y(n3596) );
  INVX1 U4760 ( .A(n3623), .Y(n3589) );
  INVX1 U4761 ( .A(n3618), .Y(n3602) );
  INVX1 U4762 ( .A(n3619), .Y(n3597) );
  INVX1 U4763 ( .A(n3620), .Y(n3595) );
  INVX1 U4764 ( .A(n3614), .Y(n3611) );
  INVX1 U4765 ( .A(n3621), .Y(n3591) );
  INVX1 U4766 ( .A(n3617), .Y(n3605) );
  INVX1 U4767 ( .A(n3620), .Y(n3594) );
  INVX1 U4768 ( .A(n3621), .Y(n3593) );
  INVX1 U4769 ( .A(n3618), .Y(n3601) );
  INVX1 U4770 ( .A(n3618), .Y(n3600) );
  INVX1 U4771 ( .A(n3619), .Y(n3598) );
  INVX1 U4772 ( .A(n3617), .Y(n3603) );
  INVX1 U4773 ( .A(n3617), .Y(n3604) );
  INVX1 U4774 ( .A(n3619), .Y(n3599) );
  INVX1 U4775 ( .A(n3621), .Y(n3592) );
  INVX1 U4776 ( .A(n3623), .Y(n3590) );
  INVX1 U4777 ( .A(n3623), .Y(n3588) );
  INVX1 U4778 ( .A(n3614), .Y(n3613) );
  INVX1 U4779 ( .A(n3614), .Y(n3612) );
  INVX1 U4780 ( .A(n3616), .Y(n3610) );
  INVX1 U4781 ( .A(n3616), .Y(n3609) );
  INVX1 U4782 ( .A(n3616), .Y(n3608) );
  NOR2X2 U4783 ( .A(n3472), .B(n3457), .Y(n13858) );
  NOR2X2 U4784 ( .A(n2871), .B(n2862), .Y(n17008) );
  NOR2X2 U4785 ( .A(n2629), .B(n2614), .Y(n18268) );
  NOR2X2 U4786 ( .A(n3231), .B(n3222), .Y(n15118) );
  NOR2X2 U4787 ( .A(n3170), .B(n3155), .Y(n15433) );
  NOR2X2 U4788 ( .A(n2932), .B(n2917), .Y(n16693) );
  NOR2X2 U4789 ( .A(n2568), .B(n2553), .Y(n18583) );
  NOR2X2 U4790 ( .A(n3292), .B(n3277), .Y(n14803) );
  NOR2X2 U4791 ( .A(n2993), .B(n2978), .Y(n16378) );
  NOR2X2 U4792 ( .A(n2690), .B(n2681), .Y(n17953) );
  NOR2X2 U4793 ( .A(n3353), .B(n3338), .Y(n14488) );
  NOR2X2 U4794 ( .A(n3051), .B(n3036), .Y(n16063) );
  NOR2X2 U4795 ( .A(n2750), .B(n2741), .Y(n17638) );
  NOR2X2 U4796 ( .A(n3411), .B(n3396), .Y(n14173) );
  NOR2X2 U4797 ( .A(n3112), .B(n3103), .Y(n15748) );
  NOR2X2 U4798 ( .A(n2811), .B(n2796), .Y(n17323) );
  NAND2X2 U4799 ( .A(n586), .B(n9913), .Y(n9958) );
  NAND2X2 U4800 ( .A(n585), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n143) );
  NAND2X2 U4801 ( .A(n587), .B(n11081), .Y(n11126) );
  NAND2X2 U4802 ( .A(n588), .B(n8161), .Y(n8206) );
  NAND2X2 U4803 ( .A(n589), .B(n10789), .Y(n10834) );
  NAND2X2 U4804 ( .A(n590), .B(n9037), .Y(n9082) );
  NAND2X2 U4805 ( .A(n591), .B(n7285), .Y(n7330) );
  NAND2X2 U4806 ( .A(n592), .B(n10205), .Y(n10250) );
  NAND2X2 U4807 ( .A(n593), .B(n9329), .Y(n9374) );
  NAND2X2 U4808 ( .A(n594), .B(n8453), .Y(n8498) );
  NAND2X2 U4809 ( .A(n595), .B(n7577), .Y(n7622) );
  NAND2X2 U4810 ( .A(n596), .B(n11373), .Y(n11418) );
  NAND2X2 U4811 ( .A(n597), .B(n10497), .Y(n10542) );
  NAND2X2 U4812 ( .A(n598), .B(n9621), .Y(n9666) );
  NAND2X2 U4813 ( .A(n599), .B(n8745), .Y(n8790) );
  NAND2X2 U4814 ( .A(n600), .B(n7869), .Y(n7914) );
  NAND2X2 U4815 ( .A(n2875), .B(n2867), .Y(n9917) );
  NAND2X2 U4816 ( .A(n3478), .B(n3467), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n101) );
  NAND2X2 U4817 ( .A(n2633), .B(n2625), .Y(n11085) );
  NAND2X2 U4818 ( .A(n3234), .B(n3227), .Y(n8165) );
  NAND2X2 U4819 ( .A(n2694), .B(n2686), .Y(n10793) );
  NAND2X2 U4820 ( .A(n3055), .B(n3047), .Y(n9041) );
  NAND2X2 U4821 ( .A(n3415), .B(n3407), .Y(n7289) );
  NAND2X2 U4822 ( .A(n2817), .B(n2807), .Y(n10209) );
  NAND2X2 U4823 ( .A(n2997), .B(n2989), .Y(n9333) );
  NAND2X2 U4824 ( .A(n3173), .B(n3166), .Y(n8457) );
  NAND2X2 U4825 ( .A(n3356), .B(n3349), .Y(n7581) );
  NAND2X2 U4826 ( .A(n2572), .B(n2564), .Y(n11377) );
  NAND2X2 U4827 ( .A(n2753), .B(n2746), .Y(n10501) );
  NAND2X2 U4828 ( .A(n2936), .B(n2928), .Y(n9625) );
  NAND2X2 U4829 ( .A(n3116), .B(n3108), .Y(n8749) );
  NAND2X2 U4830 ( .A(n3298), .B(n3288), .Y(n7873) );
  NAND2X2 U4831 ( .A(n2856), .B(n2872), .Y(n17035) );
  NAND2X2 U4832 ( .A(n3456), .B(n3473), .Y(n13885) );
  NAND2X2 U4833 ( .A(n2619), .B(n2630), .Y(n18295) );
  NAND2X2 U4834 ( .A(n3216), .B(n3232), .Y(n15145) );
  NAND2X2 U4835 ( .A(n3160), .B(n3171), .Y(n15460) );
  NAND2X2 U4836 ( .A(n2560), .B(n2569), .Y(n18610) );
  NAND2X2 U4837 ( .A(n2922), .B(n2933), .Y(n16720) );
  NAND2X2 U4838 ( .A(n3282), .B(n3293), .Y(n14830) );
  NAND2X2 U4839 ( .A(n2983), .B(n2994), .Y(n16405) );
  NAND2X2 U4840 ( .A(n2675), .B(n2691), .Y(n17980) );
  NAND2X2 U4841 ( .A(n3343), .B(n3354), .Y(n14515) );
  NAND2X2 U4842 ( .A(n3041), .B(n3052), .Y(n16090) );
  NAND2X2 U4843 ( .A(n2735), .B(n2751), .Y(n17665) );
  NAND2X2 U4844 ( .A(n3401), .B(n3412), .Y(n14200) );
  NAND2X2 U4845 ( .A(n3097), .B(n3113), .Y(n15775) );
  NAND2X2 U4846 ( .A(n2801), .B(n2812), .Y(n17350) );
  NAND2X2 U4847 ( .A(n3464), .B(n3492), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n78) );
  NAND2X2 U4848 ( .A(n2856), .B(n2891), .Y(n9895) );
  NAND2X2 U4849 ( .A(n2614), .B(n2641), .Y(n11063) );
  NAND2X2 U4850 ( .A(n3216), .B(n3248), .Y(n8143) );
  NAND2X2 U4851 ( .A(n2675), .B(n2703), .Y(n10771) );
  NAND2X2 U4852 ( .A(n3036), .B(n3063), .Y(n9019) );
  NAND2X2 U4853 ( .A(n3396), .B(n3423), .Y(n7267) );
  NAND2X2 U4854 ( .A(n2796), .B(n2823), .Y(n10187) );
  NAND2X2 U4855 ( .A(n2978), .B(n3010), .Y(n9311) );
  NAND2X2 U4856 ( .A(n3155), .B(n3183), .Y(n8435) );
  NAND2X2 U4857 ( .A(n3338), .B(n3366), .Y(n7559) );
  NAND2X2 U4858 ( .A(n2551), .B(n2581), .Y(n11355) );
  NAND2X2 U4859 ( .A(n2735), .B(n2763), .Y(n10479) );
  NAND2X2 U4860 ( .A(n2917), .B(n2944), .Y(n9603) );
  NAND2X2 U4861 ( .A(n3097), .B(n3125), .Y(n8727) );
  NAND2X2 U4862 ( .A(n3277), .B(n3309), .Y(n7851) );
  NAND2X1 U4863 ( .A(n586), .B(n9900), .Y(n9950) );
  NAND2X1 U4864 ( .A(n585), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n135) );
  NAND2X1 U4865 ( .A(n587), .B(n11068), .Y(n11118) );
  NAND2X1 U4866 ( .A(n588), .B(n8148), .Y(n8198) );
  NAND2X1 U4867 ( .A(n589), .B(n10776), .Y(n10826) );
  NAND2X1 U4868 ( .A(n590), .B(n9024), .Y(n9074) );
  NAND2X1 U4869 ( .A(n591), .B(n7272), .Y(n7322) );
  NAND2X1 U4870 ( .A(n592), .B(n10192), .Y(n10242) );
  NAND2X1 U4871 ( .A(n593), .B(n9316), .Y(n9366) );
  NAND2X1 U4872 ( .A(n594), .B(n8440), .Y(n8490) );
  NAND2X1 U4873 ( .A(n595), .B(n7564), .Y(n7614) );
  NAND2X1 U4874 ( .A(n596), .B(n11360), .Y(n11410) );
  NAND2X1 U4875 ( .A(n597), .B(n10484), .Y(n10534) );
  NAND2X1 U4876 ( .A(n598), .B(n9608), .Y(n9658) );
  NAND2X1 U4877 ( .A(n599), .B(n8732), .Y(n8782) );
  NAND2X1 U4878 ( .A(n600), .B(n7856), .Y(n7906) );
  NOR2X1 U4879 ( .A(n57), .B(n513), .Y(n17020) );
  NOR2X1 U4880 ( .A(n58), .B(n514), .Y(n13870) );
  NOR2X1 U4881 ( .A(n59), .B(n515), .Y(n18280) );
  NOR2X1 U4882 ( .A(n60), .B(n516), .Y(n15130) );
  NOR2X1 U4883 ( .A(n61), .B(n517), .Y(n15445) );
  NOR2X1 U4884 ( .A(n63), .B(n518), .Y(n18595) );
  NOR2X1 U4885 ( .A(n62), .B(n519), .Y(n16705) );
  NOR2X1 U4886 ( .A(n64), .B(n520), .Y(n14815) );
  NOR2X1 U4887 ( .A(n65), .B(n521), .Y(n16390) );
  NOR2X1 U4888 ( .A(n66), .B(n522), .Y(n17965) );
  NOR2X1 U4889 ( .A(n67), .B(n523), .Y(n14500) );
  NOR2X1 U4890 ( .A(n68), .B(n524), .Y(n16075) );
  NOR2X1 U4891 ( .A(n69), .B(n525), .Y(n17650) );
  NOR2X1 U4892 ( .A(n70), .B(n526), .Y(n14185) );
  NOR2X1 U4893 ( .A(n71), .B(n527), .Y(n15760) );
  NOR2X1 U4894 ( .A(n72), .B(n528), .Y(n17335) );
  NOR2X1 U4895 ( .A(n2871), .B(n2866), .Y(n17175) );
  NOR2X1 U4896 ( .A(n3472), .B(n3467), .Y(n14025) );
  NOR2X1 U4897 ( .A(n2629), .B(n2624), .Y(n18435) );
  NOR2X1 U4898 ( .A(n3231), .B(n3226), .Y(n15285) );
  NOR2X1 U4899 ( .A(n3170), .B(n3165), .Y(n15600) );
  NOR2X1 U4900 ( .A(n2932), .B(n2927), .Y(n16860) );
  NOR2X1 U4901 ( .A(n2568), .B(n2563), .Y(n18750) );
  NOR2X1 U4902 ( .A(n3292), .B(n3287), .Y(n14970) );
  NOR2X1 U4903 ( .A(n2993), .B(n2988), .Y(n16545) );
  NOR2X1 U4904 ( .A(n2690), .B(n2685), .Y(n18120) );
  NOR2X1 U4905 ( .A(n3353), .B(n3348), .Y(n14655) );
  NOR2X1 U4906 ( .A(n3051), .B(n3046), .Y(n16230) );
  NOR2X1 U4907 ( .A(n2750), .B(n2745), .Y(n17805) );
  NOR2X1 U4908 ( .A(n3411), .B(n3406), .Y(n14340) );
  NOR2X1 U4909 ( .A(n3112), .B(n3107), .Y(n15915) );
  NOR2X1 U4910 ( .A(n2811), .B(n2806), .Y(n17490) );
  NOR2X1 U4911 ( .A(n450), .B(n2874), .Y(n17065) );
  NOR2X1 U4912 ( .A(n449), .B(n3474), .Y(n13915) );
  NOR2X1 U4913 ( .A(n452), .B(n3233), .Y(n15175) );
  NOR2X1 U4914 ( .A(n451), .B(n2632), .Y(n18325) );
  NOR2X1 U4915 ( .A(n453), .B(n3172), .Y(n15490) );
  NOR2X1 U4916 ( .A(n454), .B(n2571), .Y(n18640) );
  NOR2X1 U4917 ( .A(n455), .B(n2939), .Y(n16750) );
  NOR2X1 U4918 ( .A(n456), .B(n3298), .Y(n14860) );
  NOR2X1 U4919 ( .A(n457), .B(n3000), .Y(n16435) );
  NOR2X1 U4920 ( .A(n458), .B(n2697), .Y(n18010) );
  NOR2X1 U4921 ( .A(n459), .B(n3355), .Y(n14545) );
  NOR2X1 U4922 ( .A(n460), .B(n3054), .Y(n16120) );
  NOR2X1 U4923 ( .A(n461), .B(n2752), .Y(n17695) );
  NOR2X1 U4924 ( .A(n462), .B(n3418), .Y(n14230) );
  NOR2X1 U4925 ( .A(n463), .B(n3115), .Y(n15805) );
  NOR2X1 U4926 ( .A(n464), .B(n2817), .Y(n17380) );
  NOR2X1 U4927 ( .A(n1137), .B(n6125), .Y(n14073) );
  NOR2X1 U4928 ( .A(n998), .B(n5357), .Y(n17223) );
  NOR2X1 U4929 ( .A(n942), .B(n5003), .Y(n18483) );
  NOR2X1 U4930 ( .A(n1082), .B(n5829), .Y(n15333) );
  NOR2X1 U4931 ( .A(n1068), .B(n5745), .Y(n15648) );
  NOR2X1 U4932 ( .A(n928), .B(n4887), .Y(n18798) );
  NOR2X1 U4933 ( .A(n1012), .B(n5441), .Y(n16908) );
  NOR2X1 U4934 ( .A(n1096), .B(n5905), .Y(n15018) );
  NOR2X1 U4935 ( .A(n1026), .B(n5517), .Y(n16593) );
  NOR2X1 U4936 ( .A(n956), .B(n5087), .Y(n18168) );
  NOR2X1 U4937 ( .A(n1110), .B(n5981), .Y(n14703) );
  NOR2X1 U4938 ( .A(n1040), .B(n5593), .Y(n16278) );
  NOR2X1 U4939 ( .A(n970), .B(n5195), .Y(n17853) );
  NOR2X1 U4940 ( .A(n1124), .B(n6057), .Y(n14388) );
  NOR2X1 U4941 ( .A(n1054), .B(n5669), .Y(n15963) );
  NOR2X1 U4942 ( .A(n984), .B(n5273), .Y(n17538) );
  NOR2X1 U4943 ( .A(n17014), .B(n1003), .Y(n17058) );
  NOR2X1 U4944 ( .A(n13864), .B(n1142), .Y(n13908) );
  NOR2X1 U4945 ( .A(n18274), .B(n947), .Y(n18318) );
  NOR2X1 U4946 ( .A(n15124), .B(n1087), .Y(n15168) );
  NOR2X1 U4947 ( .A(n15439), .B(n1073), .Y(n15483) );
  NOR2X1 U4948 ( .A(n18589), .B(n933), .Y(n18633) );
  NOR2X1 U4949 ( .A(n16699), .B(n1017), .Y(n16743) );
  NOR2X1 U4950 ( .A(n14809), .B(n1101), .Y(n14853) );
  NOR2X1 U4951 ( .A(n16384), .B(n1031), .Y(n16428) );
  NOR2X1 U4952 ( .A(n17959), .B(n961), .Y(n18003) );
  NOR2X1 U4953 ( .A(n14494), .B(n1115), .Y(n14538) );
  NOR2X1 U4954 ( .A(n16069), .B(n1045), .Y(n16113) );
  NOR2X1 U4955 ( .A(n17644), .B(n975), .Y(n17688) );
  NOR2X1 U4956 ( .A(n14179), .B(n1129), .Y(n14223) );
  NOR2X1 U4957 ( .A(n15754), .B(n1059), .Y(n15798) );
  NOR2X1 U4958 ( .A(n17329), .B(n989), .Y(n17373) );
  NAND2X1 U4959 ( .A(n529), .B(n5341), .Y(n9885) );
  NAND2X1 U4960 ( .A(n530), .B(n6137), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n67) );
  NAND2X1 U4961 ( .A(n531), .B(n4987), .Y(n11053) );
  NAND2X1 U4962 ( .A(n532), .B(n5813), .Y(n8133) );
  NAND2X1 U4963 ( .A(n533), .B(n5071), .Y(n10761) );
  NAND2X1 U4964 ( .A(n534), .B(n5577), .Y(n9009) );
  NAND2X1 U4965 ( .A(n535), .B(n6041), .Y(n7257) );
  NAND2X1 U4966 ( .A(n536), .B(n5257), .Y(n10177) );
  NAND2X1 U4967 ( .A(n537), .B(n5501), .Y(n9301) );
  NAND2X1 U4968 ( .A(n538), .B(n5729), .Y(n8425) );
  NAND2X1 U4969 ( .A(n539), .B(n5965), .Y(n7549) );
  NAND2X1 U4970 ( .A(n540), .B(n4871), .Y(n11345) );
  NAND2X1 U4971 ( .A(n541), .B(n5179), .Y(n10469) );
  NAND2X1 U4972 ( .A(n542), .B(n5425), .Y(n9593) );
  NAND2X1 U4973 ( .A(n543), .B(n5653), .Y(n8717) );
  NAND2X1 U4974 ( .A(n544), .B(n5889), .Y(n7841) );
  NOR2X1 U4975 ( .A(n450), .B(n2854), .Y(n17010) );
  NOR2X1 U4976 ( .A(n449), .B(n3457), .Y(n13860) );
  NOR2X1 U4977 ( .A(n451), .B(n2614), .Y(n18270) );
  NOR2X1 U4978 ( .A(n452), .B(n3214), .Y(n15120) );
  NOR2X1 U4979 ( .A(n453), .B(n3155), .Y(n15435) );
  NOR2X1 U4980 ( .A(n455), .B(n2917), .Y(n16695) );
  NOR2X1 U4981 ( .A(n454), .B(n2553), .Y(n18585) );
  NOR2X1 U4982 ( .A(n456), .B(n3277), .Y(n14805) );
  NOR2X1 U4983 ( .A(n457), .B(n2978), .Y(n16380) );
  NOR2X1 U4984 ( .A(n458), .B(n2673), .Y(n17955) );
  NOR2X1 U4985 ( .A(n459), .B(n3338), .Y(n14490) );
  NOR2X1 U4986 ( .A(n460), .B(n3036), .Y(n16065) );
  NOR2X1 U4987 ( .A(n461), .B(n2733), .Y(n17640) );
  NOR2X1 U4988 ( .A(n462), .B(n3396), .Y(n14175) );
  NOR2X1 U4989 ( .A(n463), .B(n3095), .Y(n15750) );
  NOR2X1 U4990 ( .A(n464), .B(n2796), .Y(n17325) );
  NAND2X1 U4991 ( .A(n5341), .B(n2904), .Y(n10011) );
  NAND2X1 U4992 ( .A(n6137), .B(n3506), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n197) );
  NAND2X1 U4993 ( .A(n4987), .B(n2662), .Y(n11179) );
  NAND2X1 U4994 ( .A(n5813), .B(n3264), .Y(n8259) );
  NAND2X1 U4995 ( .A(n5071), .B(n2722), .Y(n10887) );
  NAND2X1 U4996 ( .A(n5577), .B(n3084), .Y(n9135) );
  NAND2X1 U4997 ( .A(n6041), .B(n3444), .Y(n7383) );
  NAND2X1 U4998 ( .A(n5257), .B(n2845), .Y(n10303) );
  NAND2X1 U4999 ( .A(n5501), .B(n3024), .Y(n9427) );
  NAND2X1 U5000 ( .A(n5729), .B(n3203), .Y(n8551) );
  NAND2X1 U5001 ( .A(n5965), .B(n3384), .Y(n7675) );
  NAND2X1 U5002 ( .A(n4871), .B(n2601), .Y(n11471) );
  NAND2X1 U5003 ( .A(n5179), .B(n2777), .Y(n10595) );
  NAND2X1 U5004 ( .A(n5425), .B(n2965), .Y(n9719) );
  NAND2X1 U5005 ( .A(n5653), .B(n3143), .Y(n8843) );
  NAND2X1 U5006 ( .A(n5889), .B(n3315), .Y(n7967) );
  NAND2X1 U5007 ( .A(n998), .B(n1003), .Y(n17114) );
  NAND2X1 U5008 ( .A(n1137), .B(n1142), .Y(n13964) );
  NAND2X1 U5009 ( .A(n942), .B(n947), .Y(n18374) );
  NAND2X1 U5010 ( .A(n1082), .B(n1087), .Y(n15224) );
  NAND2X1 U5011 ( .A(n1068), .B(n1073), .Y(n15539) );
  NAND2X1 U5012 ( .A(n928), .B(n933), .Y(n18689) );
  NAND2X1 U5013 ( .A(n1012), .B(n1017), .Y(n16799) );
  NAND2X1 U5014 ( .A(n1096), .B(n1101), .Y(n14909) );
  NAND2X1 U5015 ( .A(n1026), .B(n1031), .Y(n16484) );
  NAND2X1 U5016 ( .A(n956), .B(n961), .Y(n18059) );
  NAND2X1 U5017 ( .A(n1110), .B(n1115), .Y(n14594) );
  NAND2X1 U5018 ( .A(n1040), .B(n1045), .Y(n16169) );
  NAND2X1 U5019 ( .A(n970), .B(n975), .Y(n17744) );
  NAND2X1 U5020 ( .A(n1124), .B(n1129), .Y(n14279) );
  NAND2X1 U5021 ( .A(n1054), .B(n1059), .Y(n15854) );
  NAND2X1 U5022 ( .A(n984), .B(n989), .Y(n17429) );
  NAND2X1 U5023 ( .A(n1137), .B(n3493), .Y(n13941) );
  NAND2X1 U5024 ( .A(n998), .B(n2893), .Y(n17091) );
  NAND2X1 U5025 ( .A(n942), .B(n2650), .Y(n18351) );
  NAND2X1 U5026 ( .A(n1082), .B(n3253), .Y(n15201) );
  NAND2X1 U5027 ( .A(n1068), .B(n3192), .Y(n15516) );
  NAND2X1 U5028 ( .A(n1012), .B(n2954), .Y(n16776) );
  NAND2X1 U5029 ( .A(n928), .B(n2598), .Y(n18666) );
  NAND2X1 U5030 ( .A(n1096), .B(n3314), .Y(n14886) );
  NAND2X1 U5031 ( .A(n1026), .B(n3015), .Y(n16461) );
  NAND2X1 U5032 ( .A(n956), .B(n2711), .Y(n18036) );
  NAND2X1 U5033 ( .A(n1110), .B(n3375), .Y(n14571) );
  NAND2X1 U5034 ( .A(n1040), .B(n3072), .Y(n16146) );
  NAND2X1 U5035 ( .A(n970), .B(n2772), .Y(n17721) );
  NAND2X1 U5036 ( .A(n1124), .B(n3433), .Y(n14256) );
  NAND2X1 U5037 ( .A(n1054), .B(n3134), .Y(n15831) );
  NAND2X1 U5038 ( .A(n984), .B(n2833), .Y(n17406) );
  NOR2XL U5039 ( .A(n57), .B(n337), .Y(n17121) );
  NOR2XL U5040 ( .A(n58), .B(n338), .Y(n13971) );
  NOR2XL U5041 ( .A(n59), .B(n339), .Y(n18381) );
  NOR2XL U5042 ( .A(n60), .B(n340), .Y(n15231) );
  NOR2XL U5043 ( .A(n61), .B(n341), .Y(n15546) );
  NOR2XL U5044 ( .A(n62), .B(n342), .Y(n16806) );
  NOR2XL U5045 ( .A(n63), .B(n343), .Y(n18696) );
  NOR2XL U5046 ( .A(n64), .B(n344), .Y(n14916) );
  NOR2XL U5047 ( .A(n65), .B(n345), .Y(n16491) );
  NOR2XL U5048 ( .A(n66), .B(n346), .Y(n18066) );
  NOR2XL U5049 ( .A(n67), .B(n347), .Y(n14601) );
  NOR2XL U5050 ( .A(n68), .B(n348), .Y(n16176) );
  NOR2XL U5051 ( .A(n69), .B(n349), .Y(n17751) );
  NOR2XL U5052 ( .A(n70), .B(n350), .Y(n14286) );
  NOR2XL U5053 ( .A(n71), .B(n351), .Y(n15861) );
  NOR2XL U5054 ( .A(n72), .B(n352), .Y(n17436) );
  AOI31X1 U5055 ( .A0(n3495), .A1(n3453), .A2(n1136), .B0(n13862), .Y(n14119)
         );
  AOI31X1 U5056 ( .A0(n2895), .A1(n2852), .A2(n997), .B0(n17012), .Y(n17269)
         );
  AOI31X1 U5057 ( .A0(n2652), .A1(n2610), .A2(n941), .B0(n18272), .Y(n18529)
         );
  AOI31X1 U5058 ( .A0(n3255), .A1(n3212), .A2(n1081), .B0(n15122), .Y(n15379)
         );
  AOI31X1 U5059 ( .A0(n3194), .A1(n3151), .A2(n1067), .B0(n15437), .Y(n15694)
         );
  AOI31X1 U5060 ( .A0(n2591), .A1(n2549), .A2(n927), .B0(n18587), .Y(n18844)
         );
  AOI31X1 U5061 ( .A0(n2956), .A1(n2913), .A2(n1011), .B0(n16697), .Y(n16954)
         );
  AOI31X1 U5062 ( .A0(n3317), .A1(n3273), .A2(n1095), .B0(n14807), .Y(n15064)
         );
  AOI31X1 U5063 ( .A0(n3019), .A1(n2974), .A2(n1025), .B0(n16382), .Y(n16639)
         );
  AOI31X1 U5064 ( .A0(n2712), .A1(n2671), .A2(n955), .B0(n17957), .Y(n18214)
         );
  AOI31X1 U5065 ( .A0(n3379), .A1(n3334), .A2(n1109), .B0(n14492), .Y(n14749)
         );
  AOI31X1 U5066 ( .A0(n3074), .A1(n3032), .A2(n1039), .B0(n16067), .Y(n16324)
         );
  AOI31X1 U5067 ( .A0(n2778), .A1(n2731), .A2(n969), .B0(n17642), .Y(n17899)
         );
  AOI31X1 U5068 ( .A0(n3434), .A1(n3392), .A2(n1123), .B0(n14177), .Y(n14434)
         );
  AOI31X1 U5069 ( .A0(n3138), .A1(n3093), .A2(n1053), .B0(n15752), .Y(n16009)
         );
  AOI31X1 U5070 ( .A0(n2838), .A1(n2792), .A2(n983), .B0(n17327), .Y(n17584)
         );
  NAND2X1 U5071 ( .A(n5341), .B(n2881), .Y(n10065) );
  NAND2X1 U5072 ( .A(n6137), .B(n3482), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n251) );
  NAND2X1 U5073 ( .A(n4987), .B(n2639), .Y(n11233) );
  NAND2X1 U5074 ( .A(n5813), .B(n3241), .Y(n8313) );
  NAND2X1 U5075 ( .A(n5071), .B(n2700), .Y(n10941) );
  NAND2X1 U5076 ( .A(n6041), .B(n3421), .Y(n7437) );
  NAND2X1 U5077 ( .A(n5577), .B(n3061), .Y(n9189) );
  NAND2X1 U5078 ( .A(n5257), .B(n2821), .Y(n10357) );
  NAND2X1 U5079 ( .A(n5501), .B(n3003), .Y(n9481) );
  NAND2X1 U5080 ( .A(n5729), .B(n3180), .Y(n8605) );
  NAND2X1 U5081 ( .A(n5965), .B(n3363), .Y(n7729) );
  NAND2X1 U5082 ( .A(n4871), .B(n2578), .Y(n11525) );
  NAND2X1 U5083 ( .A(n5179), .B(n2760), .Y(n10649) );
  NAND2X1 U5084 ( .A(n5425), .B(n2942), .Y(n9773) );
  NAND2X1 U5085 ( .A(n5653), .B(n3122), .Y(n8897) );
  NAND2X1 U5086 ( .A(n5889), .B(n3302), .Y(n8021) );
  NAND2X1 U5087 ( .A(n5362), .B(n2904), .Y(n17155) );
  NAND2X1 U5088 ( .A(n6130), .B(n3496), .Y(n14005) );
  NAND2X1 U5089 ( .A(n5008), .B(n2662), .Y(n18415) );
  NAND2X1 U5090 ( .A(n5834), .B(n3264), .Y(n15265) );
  NAND2X1 U5091 ( .A(n5750), .B(n3203), .Y(n15580) );
  NAND2X1 U5092 ( .A(n4892), .B(n2601), .Y(n18730) );
  NAND2X1 U5093 ( .A(n5446), .B(n2965), .Y(n16840) );
  NAND2X1 U5094 ( .A(n5910), .B(n3319), .Y(n14950) );
  NAND2X1 U5095 ( .A(n5522), .B(n3024), .Y(n16525) );
  NAND2X1 U5096 ( .A(n5092), .B(n2722), .Y(n18100) );
  NAND2X1 U5097 ( .A(n5986), .B(n3384), .Y(n14635) );
  NAND2X1 U5098 ( .A(n5598), .B(n3084), .Y(n16210) );
  NAND2X1 U5099 ( .A(n5200), .B(n2781), .Y(n17785) );
  NAND2X1 U5100 ( .A(n6062), .B(n3444), .Y(n14320) );
  NAND2X1 U5101 ( .A(n5674), .B(n3143), .Y(n15895) );
  NAND2X1 U5102 ( .A(n5278), .B(n2845), .Y(n17470) );
  AOI22X1 U5103 ( .A0(n450), .A1(n996), .B0(n353), .B1(n5350), .Y(n10099) );
  AOI22X1 U5104 ( .A0(n449), .A1(n1139), .B0(n354), .B1(n6146), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n285) );
  AOI22X1 U5105 ( .A0(n452), .A1(n1080), .B0(n355), .B1(n5822), .Y(n8347) );
  AOI22X1 U5106 ( .A0(n451), .A1(n940), .B0(n356), .B1(n4996), .Y(n11267) );
  AOI22X1 U5107 ( .A0(n458), .A1(n954), .B0(n357), .B1(n5080), .Y(n10975) );
  AOI22X1 U5108 ( .A0(n462), .A1(n1122), .B0(n358), .B1(n6050), .Y(n7471) );
  AOI22X1 U5109 ( .A0(n460), .A1(n1038), .B0(n359), .B1(n5586), .Y(n9223) );
  AOI22X1 U5110 ( .A0(n464), .A1(n982), .B0(n360), .B1(n5266), .Y(n10391) );
  AOI22X1 U5111 ( .A0(n457), .A1(n1024), .B0(n361), .B1(n5510), .Y(n9515) );
  AOI22X1 U5112 ( .A0(n453), .A1(n1066), .B0(n362), .B1(n5738), .Y(n8639) );
  AOI22X1 U5113 ( .A0(n459), .A1(n1108), .B0(n363), .B1(n5974), .Y(n7763) );
  AOI22X1 U5114 ( .A0(n454), .A1(n926), .B0(n364), .B1(n4880), .Y(n11559) );
  AOI22X1 U5115 ( .A0(n461), .A1(n968), .B0(n365), .B1(n5188), .Y(n10683) );
  AOI22X1 U5116 ( .A0(n455), .A1(n1010), .B0(n366), .B1(n5434), .Y(n9807) );
  AOI22X1 U5117 ( .A0(n463), .A1(n1052), .B0(n367), .B1(n5662), .Y(n8931) );
  AOI22X1 U5118 ( .A0(n456), .A1(n1094), .B0(n368), .B1(n5898), .Y(n8055) );
  AOI31X1 U5119 ( .A0(n386), .A1(n2867), .A2(n17008), .B0(n5331), .Y(n17281)
         );
  INVX1 U5120 ( .A(n17085), .Y(n5331) );
  AOI31X1 U5121 ( .A0(n385), .A1(n3468), .A2(n13858), .B0(n6115), .Y(n14131)
         );
  INVX1 U5122 ( .A(n13935), .Y(n6115) );
  AOI31X1 U5123 ( .A0(n388), .A1(n3227), .A2(n15118), .B0(n5803), .Y(n15391)
         );
  INVX1 U5124 ( .A(n15195), .Y(n5803) );
  AOI31X1 U5125 ( .A0(n387), .A1(n2625), .A2(n18268), .B0(n4977), .Y(n18541)
         );
  INVX1 U5126 ( .A(n18345), .Y(n4977) );
  AOI31X1 U5127 ( .A0(n389), .A1(n3166), .A2(n15433), .B0(n5719), .Y(n15706)
         );
  INVX1 U5128 ( .A(n15510), .Y(n5719) );
  AOI31X1 U5129 ( .A0(n391), .A1(n2928), .A2(n16693), .B0(n5415), .Y(n16966)
         );
  INVX1 U5130 ( .A(n16770), .Y(n5415) );
  AOI31X1 U5131 ( .A0(n390), .A1(n2564), .A2(n18583), .B0(n4861), .Y(n18856)
         );
  INVX1 U5132 ( .A(n18660), .Y(n4861) );
  AOI31X1 U5133 ( .A0(n392), .A1(n3288), .A2(n14803), .B0(n5879), .Y(n15076)
         );
  INVX1 U5134 ( .A(n14880), .Y(n5879) );
  AOI31X1 U5135 ( .A0(n393), .A1(n2989), .A2(n16378), .B0(n5491), .Y(n16651)
         );
  INVX1 U5136 ( .A(n16455), .Y(n5491) );
  AOI31X1 U5137 ( .A0(n394), .A1(n2686), .A2(n17953), .B0(n5061), .Y(n18226)
         );
  INVX1 U5138 ( .A(n18030), .Y(n5061) );
  AOI31X1 U5139 ( .A0(n395), .A1(n3349), .A2(n14488), .B0(n5955), .Y(n14761)
         );
  INVX1 U5140 ( .A(n14565), .Y(n5955) );
  AOI31X1 U5141 ( .A0(n396), .A1(n3047), .A2(n16063), .B0(n5567), .Y(n16336)
         );
  INVX1 U5142 ( .A(n16140), .Y(n5567) );
  AOI31X1 U5143 ( .A0(n397), .A1(n2746), .A2(n17638), .B0(n5169), .Y(n17911)
         );
  INVX1 U5144 ( .A(n17715), .Y(n5169) );
  AOI31X1 U5145 ( .A0(n398), .A1(n3407), .A2(n14173), .B0(n6031), .Y(n14446)
         );
  INVX1 U5146 ( .A(n14250), .Y(n6031) );
  AOI31X1 U5147 ( .A0(n399), .A1(n3108), .A2(n15748), .B0(n5643), .Y(n16021)
         );
  INVX1 U5148 ( .A(n15825), .Y(n5643) );
  AOI31X1 U5149 ( .A0(n400), .A1(n2807), .A2(n17323), .B0(n5247), .Y(n17596)
         );
  INVX1 U5150 ( .A(n17400), .Y(n5247) );
  NAND2X1 U5151 ( .A(n1133), .B(n3482), .Y(n13863) );
  NAND2X1 U5152 ( .A(n994), .B(n2881), .Y(n17013) );
  NAND2X1 U5153 ( .A(n938), .B(n2639), .Y(n18273) );
  NAND2X1 U5154 ( .A(n1078), .B(n3241), .Y(n15123) );
  NAND2X1 U5155 ( .A(n1064), .B(n3180), .Y(n15438) );
  NAND2X1 U5156 ( .A(n1008), .B(n2942), .Y(n16698) );
  NAND2X1 U5157 ( .A(n924), .B(n2578), .Y(n18588) );
  NAND2X1 U5158 ( .A(n1092), .B(n3302), .Y(n14808) );
  NAND2X1 U5159 ( .A(n1022), .B(n3003), .Y(n16383) );
  NAND2X1 U5160 ( .A(n952), .B(n2700), .Y(n17958) );
  NAND2X1 U5161 ( .A(n1106), .B(n3363), .Y(n14493) );
  NAND2X1 U5162 ( .A(n1036), .B(n3061), .Y(n16068) );
  NAND2X1 U5163 ( .A(n966), .B(n2760), .Y(n17643) );
  NAND2X1 U5164 ( .A(n1120), .B(n3421), .Y(n14178) );
  NAND2X1 U5165 ( .A(n1050), .B(n3122), .Y(n15753) );
  NAND2X1 U5166 ( .A(n980), .B(n2821), .Y(n17328) );
  NAND2X1 U5167 ( .A(n2875), .B(n2866), .Y(n17090) );
  NAND2X1 U5168 ( .A(n2633), .B(n2624), .Y(n18350) );
  NAND2X1 U5169 ( .A(n3235), .B(n3226), .Y(n15200) );
  NAND2X1 U5170 ( .A(n3174), .B(n3165), .Y(n15515) );
  NAND2X1 U5171 ( .A(n2936), .B(n2927), .Y(n16775) );
  NAND2X1 U5172 ( .A(n2572), .B(n2563), .Y(n18665) );
  NAND2X1 U5173 ( .A(n3295), .B(n3287), .Y(n14885) );
  NAND2X1 U5174 ( .A(n2997), .B(n2988), .Y(n16460) );
  NAND2X1 U5175 ( .A(n2694), .B(n2685), .Y(n18035) );
  NAND2X1 U5176 ( .A(n3357), .B(n3348), .Y(n14570) );
  NAND2X1 U5177 ( .A(n3055), .B(n3046), .Y(n16145) );
  NAND2X1 U5178 ( .A(n2754), .B(n2745), .Y(n17720) );
  NAND2X1 U5179 ( .A(n3415), .B(n3406), .Y(n14255) );
  NAND2X1 U5180 ( .A(n3116), .B(n3107), .Y(n15830) );
  NAND2X1 U5181 ( .A(n2814), .B(n2806), .Y(n17405) );
  NAND2X1 U5182 ( .A(n3477), .B(n3468), .Y(n13940) );
  NAND2X1 U5183 ( .A(n1135), .B(n3497), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n87) );
  NAND2X1 U5184 ( .A(n993), .B(n2899), .Y(n9904) );
  NAND2X1 U5185 ( .A(n1077), .B(n3259), .Y(n8152) );
  NAND2X1 U5186 ( .A(n937), .B(n2658), .Y(n11072) );
  NAND2X1 U5187 ( .A(n951), .B(n2713), .Y(n10780) );
  NAND2X1 U5188 ( .A(n1119), .B(n3435), .Y(n7276) );
  NAND2X1 U5189 ( .A(n1035), .B(n3080), .Y(n9028) );
  NAND2X1 U5190 ( .A(n979), .B(n2837), .Y(n10196) );
  NAND2X1 U5191 ( .A(n1021), .B(n3018), .Y(n9320) );
  NAND2X1 U5192 ( .A(n1063), .B(n3198), .Y(n8444) );
  NAND2X1 U5193 ( .A(n1105), .B(n3378), .Y(n7568) );
  NAND2X1 U5194 ( .A(n923), .B(n2597), .Y(n11364) );
  NAND2X1 U5195 ( .A(n965), .B(n2776), .Y(n10488) );
  NAND2X1 U5196 ( .A(n1007), .B(n2960), .Y(n9612) );
  NAND2X1 U5197 ( .A(n1049), .B(n3137), .Y(n8736) );
  NAND2X1 U5198 ( .A(n1091), .B(n3317), .Y(n7860) );
  NAND2X1 U5199 ( .A(n6146), .B(n3482), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n133) );
  NAND2X1 U5200 ( .A(n5350), .B(n2881), .Y(n9948) );
  NAND2X1 U5201 ( .A(n4996), .B(n2639), .Y(n11116) );
  NAND2X1 U5202 ( .A(n5822), .B(n3241), .Y(n8196) );
  NAND2X1 U5203 ( .A(n5080), .B(n2700), .Y(n10824) );
  NAND2X1 U5204 ( .A(n5586), .B(n3061), .Y(n9072) );
  NAND2X1 U5205 ( .A(n6050), .B(n3421), .Y(n7320) );
  NAND2X1 U5206 ( .A(n5266), .B(n2821), .Y(n10240) );
  NAND2X1 U5207 ( .A(n5510), .B(n3003), .Y(n9364) );
  NAND2X1 U5208 ( .A(n5738), .B(n3180), .Y(n8488) );
  NAND2X1 U5209 ( .A(n5974), .B(n3363), .Y(n7612) );
  NAND2X1 U5210 ( .A(n4880), .B(n2578), .Y(n11408) );
  NAND2X1 U5211 ( .A(n5188), .B(n2760), .Y(n10532) );
  NAND2X1 U5212 ( .A(n5434), .B(n2942), .Y(n9656) );
  NAND2X1 U5213 ( .A(n5662), .B(n3122), .Y(n8780) );
  NAND2X1 U5214 ( .A(n5898), .B(n3302), .Y(n7904) );
  AOI22XL U5215 ( .A0(n2880), .A1(n5362), .B0(n1311), .B1(n994), .Y(n17220) );
  AOI22XL U5216 ( .A0(n3481), .A1(n6130), .B0(n1281), .B1(n1133), .Y(n14070)
         );
  AOI22XL U5217 ( .A0(n3240), .A1(n5834), .B0(n1293), .B1(n1078), .Y(n15330)
         );
  AOI22XL U5218 ( .A0(n2638), .A1(n5008), .B0(n1323), .B1(n938), .Y(n18480) );
  AOI22XL U5219 ( .A0(n3179), .A1(n5750), .B0(n1296), .B1(n1064), .Y(n15645)
         );
  AOI22XL U5220 ( .A0(n2941), .A1(n5446), .B0(n1308), .B1(n1008), .Y(n16905)
         );
  AOI22XL U5221 ( .A0(n2577), .A1(n4892), .B0(n1326), .B1(n924), .Y(n18795) );
  AOI22XL U5222 ( .A0(n3301), .A1(n5910), .B0(n1290), .B1(n1092), .Y(n15015)
         );
  AOI22XL U5223 ( .A0(n3002), .A1(n5522), .B0(n1305), .B1(n1022), .Y(n16590)
         );
  AOI22XL U5224 ( .A0(n2699), .A1(n5092), .B0(n1320), .B1(n952), .Y(n18165) );
  AOI22XL U5225 ( .A0(n3362), .A1(n5986), .B0(n1287), .B1(n1106), .Y(n14700)
         );
  AOI22XL U5226 ( .A0(n3060), .A1(n5598), .B0(n1302), .B1(n1036), .Y(n16275)
         );
  AOI22XL U5227 ( .A0(n2759), .A1(n5200), .B0(n1317), .B1(n966), .Y(n17850) );
  AOI22XL U5228 ( .A0(n3420), .A1(n6062), .B0(n1284), .B1(n1120), .Y(n14385)
         );
  AOI22XL U5229 ( .A0(n3121), .A1(n5674), .B0(n1299), .B1(n1050), .Y(n15960)
         );
  AOI22XL U5230 ( .A0(n2820), .A1(n5278), .B0(n1314), .B1(n980), .Y(n17535) );
  NAND2X1 U5231 ( .A(n6156), .B(n402), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n140) );
  NAND2X1 U5232 ( .A(n5366), .B(n401), .Y(n9955) );
  NAND2X1 U5233 ( .A(n5012), .B(n403), .Y(n11123) );
  NAND2X1 U5234 ( .A(n5838), .B(n404), .Y(n8203) );
  NAND2X1 U5235 ( .A(n5096), .B(n405), .Y(n10831) );
  NAND2X1 U5236 ( .A(n5602), .B(n406), .Y(n9079) );
  NAND2X1 U5237 ( .A(n6066), .B(n407), .Y(n7327) );
  NAND2X1 U5238 ( .A(n5282), .B(n408), .Y(n10247) );
  NAND2X1 U5239 ( .A(n5526), .B(n409), .Y(n9371) );
  NAND2X1 U5240 ( .A(n5754), .B(n410), .Y(n8495) );
  NAND2X1 U5241 ( .A(n5990), .B(n411), .Y(n7619) );
  NAND2X1 U5242 ( .A(n4896), .B(n412), .Y(n11415) );
  NAND2X1 U5243 ( .A(n5204), .B(n413), .Y(n10539) );
  NAND2X1 U5244 ( .A(n5450), .B(n414), .Y(n9663) );
  NAND2X1 U5245 ( .A(n5678), .B(n415), .Y(n8787) );
  NAND2X1 U5246 ( .A(n5914), .B(n416), .Y(n7911) );
  AOI22XL U5247 ( .A0(n17061), .A1(n994), .B0(n529), .B1(n5376), .Y(n17077) );
  AOI22XL U5248 ( .A0(n13911), .A1(n1133), .B0(n530), .B1(n6166), .Y(n13927)
         );
  AOI22XL U5249 ( .A0(n18321), .A1(n938), .B0(n531), .B1(n5022), .Y(n18337) );
  AOI22XL U5250 ( .A0(n15171), .A1(n1078), .B0(n532), .B1(n5848), .Y(n15187)
         );
  AOI22XL U5251 ( .A0(n15486), .A1(n1064), .B0(n538), .B1(n5764), .Y(n15502)
         );
  AOI22XL U5252 ( .A0(n18636), .A1(n924), .B0(n540), .B1(n4906), .Y(n18652) );
  AOI22XL U5253 ( .A0(n16746), .A1(n1008), .B0(n542), .B1(n5460), .Y(n16762)
         );
  AOI22XL U5254 ( .A0(n14856), .A1(n1092), .B0(n544), .B1(n5924), .Y(n14872)
         );
  AOI22XL U5255 ( .A0(n16431), .A1(n1022), .B0(n537), .B1(n5536), .Y(n16447)
         );
  AOI22XL U5256 ( .A0(n18006), .A1(n952), .B0(n533), .B1(n5106), .Y(n18022) );
  AOI22XL U5257 ( .A0(n14541), .A1(n1106), .B0(n539), .B1(n6000), .Y(n14557)
         );
  AOI22XL U5258 ( .A0(n16116), .A1(n1036), .B0(n534), .B1(n5612), .Y(n16132)
         );
  AOI22XL U5259 ( .A0(n17691), .A1(n966), .B0(n541), .B1(n5214), .Y(n17707) );
  AOI22XL U5260 ( .A0(n14226), .A1(n1120), .B0(n535), .B1(n6076), .Y(n14242)
         );
  AOI22XL U5261 ( .A0(n15801), .A1(n1050), .B0(n543), .B1(n5688), .Y(n15817)
         );
  AOI22XL U5262 ( .A0(n17376), .A1(n980), .B0(n536), .B1(n5292), .Y(n17392) );
  NAND2X1 U5263 ( .A(n417), .B(n5366), .Y(n9923) );
  NAND2X1 U5264 ( .A(n418), .B(n6156), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n108) );
  NAND2X1 U5265 ( .A(n419), .B(n5012), .Y(n11091) );
  NAND2X1 U5266 ( .A(n420), .B(n5838), .Y(n8171) );
  NAND2X1 U5267 ( .A(n421), .B(n5096), .Y(n10799) );
  NAND2X1 U5268 ( .A(n422), .B(n5602), .Y(n9047) );
  NAND2X1 U5269 ( .A(n423), .B(n6066), .Y(n7295) );
  NAND2X1 U5270 ( .A(n424), .B(n5282), .Y(n10215) );
  NAND2X1 U5271 ( .A(n425), .B(n5526), .Y(n9339) );
  NAND2X1 U5272 ( .A(n426), .B(n5754), .Y(n8463) );
  NAND2X1 U5273 ( .A(n427), .B(n5990), .Y(n7587) );
  NAND2X1 U5274 ( .A(n428), .B(n4896), .Y(n11383) );
  NAND2X1 U5275 ( .A(n429), .B(n5204), .Y(n10507) );
  NAND2X1 U5276 ( .A(n430), .B(n5450), .Y(n9631) );
  NAND2X1 U5277 ( .A(n431), .B(n5678), .Y(n8755) );
  NAND2X1 U5278 ( .A(n432), .B(n5914), .Y(n7879) );
  OAI21XL U5279 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n71), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n143), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n75) );
  OAI21XL U5280 ( .A0(n9970), .A1(n9889), .B0(n9958), .Y(n9892) );
  OAI21XL U5281 ( .A0(n11138), .A1(n11057), .B0(n11126), .Y(n11060) );
  OAI21XL U5282 ( .A0(n8218), .A1(n8137), .B0(n8206), .Y(n8140) );
  OAI21XL U5283 ( .A0(n10846), .A1(n10765), .B0(n10834), .Y(n10768) );
  OAI21XL U5284 ( .A0(n7342), .A1(n7261), .B0(n7330), .Y(n7264) );
  OAI21XL U5285 ( .A0(n9094), .A1(n9013), .B0(n9082), .Y(n9016) );
  OAI21XL U5286 ( .A0(n10262), .A1(n10181), .B0(n10250), .Y(n10184) );
  OAI21XL U5287 ( .A0(n9386), .A1(n9305), .B0(n9374), .Y(n9308) );
  OAI21XL U5288 ( .A0(n8510), .A1(n8429), .B0(n8498), .Y(n8432) );
  OAI21XL U5289 ( .A0(n7634), .A1(n7553), .B0(n7622), .Y(n7556) );
  OAI21XL U5290 ( .A0(n11430), .A1(n11349), .B0(n11418), .Y(n11352) );
  OAI21XL U5291 ( .A0(n10554), .A1(n10473), .B0(n10542), .Y(n10476) );
  OAI21XL U5292 ( .A0(n9678), .A1(n9597), .B0(n9666), .Y(n9600) );
  OAI21XL U5293 ( .A0(n8802), .A1(n8721), .B0(n8790), .Y(n8724) );
  OAI21XL U5294 ( .A0(n7926), .A1(n7845), .B0(n7914), .Y(n7848) );
  NAND2X1 U5295 ( .A(n2866), .B(n2872), .Y(n9912) );
  NAND2X1 U5296 ( .A(n3467), .B(n3473), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n96) );
  NAND2X1 U5297 ( .A(n3226), .B(n3232), .Y(n8160) );
  NAND2X1 U5298 ( .A(n2624), .B(n2630), .Y(n11080) );
  NAND2X1 U5299 ( .A(n2685), .B(n2691), .Y(n10788) );
  NAND2X1 U5300 ( .A(n3406), .B(n3412), .Y(n7284) );
  NAND2X1 U5301 ( .A(n3046), .B(n3052), .Y(n9036) );
  NAND2X1 U5302 ( .A(n2806), .B(n2812), .Y(n10204) );
  NAND2X1 U5303 ( .A(n2988), .B(n2994), .Y(n9328) );
  NAND2X1 U5304 ( .A(n3165), .B(n3171), .Y(n8452) );
  NAND2X1 U5305 ( .A(n3348), .B(n3354), .Y(n7576) );
  NAND2X1 U5306 ( .A(n2563), .B(n2569), .Y(n11372) );
  NAND2X1 U5307 ( .A(n2745), .B(n2751), .Y(n10496) );
  NAND2X1 U5308 ( .A(n2927), .B(n2933), .Y(n9620) );
  NAND2X1 U5309 ( .A(n3107), .B(n3113), .Y(n8744) );
  NAND2X1 U5310 ( .A(n3287), .B(n3293), .Y(n7868) );
  NAND2X1 U5311 ( .A(n1001), .B(n5341), .Y(n10045) );
  NAND2X1 U5312 ( .A(n1143), .B(n6137), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n231) );
  NAND2X1 U5313 ( .A(n945), .B(n4987), .Y(n11213) );
  NAND2X1 U5314 ( .A(n1085), .B(n5813), .Y(n8293) );
  NAND2X1 U5315 ( .A(n959), .B(n5071), .Y(n10921) );
  NAND2X1 U5316 ( .A(n1043), .B(n5577), .Y(n9169) );
  NAND2X1 U5317 ( .A(n1127), .B(n6041), .Y(n7417) );
  NAND2X1 U5318 ( .A(n987), .B(n5257), .Y(n10337) );
  NAND2X1 U5319 ( .A(n1029), .B(n5501), .Y(n9461) );
  NAND2X1 U5320 ( .A(n1071), .B(n5729), .Y(n8585) );
  NAND2X1 U5321 ( .A(n1113), .B(n5965), .Y(n7709) );
  NAND2X1 U5322 ( .A(n931), .B(n4871), .Y(n11505) );
  NAND2X1 U5323 ( .A(n973), .B(n5179), .Y(n10629) );
  NAND2X1 U5324 ( .A(n1015), .B(n5425), .Y(n9753) );
  NAND2X1 U5325 ( .A(n1057), .B(n5653), .Y(n8877) );
  NAND2X1 U5326 ( .A(n1099), .B(n5889), .Y(n8001) );
  AOI21X1 U5327 ( .A0(n466), .A1(n1139), .B0(n6137), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n274) );
  AOI21X1 U5328 ( .A0(n465), .A1(n996), .B0(n5341), .Y(n10088) );
  AOI21X1 U5329 ( .A0(n467), .A1(n940), .B0(n4987), .Y(n11256) );
  AOI21X1 U5330 ( .A0(n468), .A1(n1080), .B0(n5813), .Y(n8336) );
  AOI21X1 U5331 ( .A0(n474), .A1(n954), .B0(n5071), .Y(n10964) );
  AOI21X1 U5332 ( .A0(n476), .A1(n1038), .B0(n5577), .Y(n9212) );
  AOI21X1 U5333 ( .A0(n478), .A1(n1122), .B0(n6041), .Y(n7460) );
  AOI21X1 U5334 ( .A0(n480), .A1(n982), .B0(n5257), .Y(n10380) );
  AOI21X1 U5335 ( .A0(n473), .A1(n1024), .B0(n5501), .Y(n9504) );
  AOI21X1 U5336 ( .A0(n469), .A1(n1066), .B0(n5729), .Y(n8628) );
  AOI21X1 U5337 ( .A0(n475), .A1(n1108), .B0(n5965), .Y(n7752) );
  AOI21X1 U5338 ( .A0(n471), .A1(n926), .B0(n4871), .Y(n11548) );
  AOI21X1 U5339 ( .A0(n477), .A1(n968), .B0(n5179), .Y(n10672) );
  AOI21X1 U5340 ( .A0(n470), .A1(n1010), .B0(n5425), .Y(n9796) );
  AOI21X1 U5341 ( .A0(n479), .A1(n1052), .B0(n5653), .Y(n8920) );
  AOI21X1 U5342 ( .A0(n472), .A1(n1094), .B0(n5889), .Y(n8044) );
  NAND2X1 U5343 ( .A(n686), .B(n6549), .Y(n13349) );
  NAND2X1 U5344 ( .A(n688), .B(n6844), .Y(n12719) );
  NAND2X1 U5345 ( .A(n687), .B(n6890), .Y(n13034) );
  NAND2X1 U5346 ( .A(n1137), .B(n13857), .Y(n13875) );
  NAND2X1 U5347 ( .A(n998), .B(n17007), .Y(n17025) );
  NAND2X1 U5348 ( .A(n942), .B(n18267), .Y(n18285) );
  NAND2X1 U5349 ( .A(n1082), .B(n15117), .Y(n15135) );
  NAND2X1 U5350 ( .A(n1068), .B(n15432), .Y(n15450) );
  NAND2X1 U5351 ( .A(n928), .B(n18582), .Y(n18600) );
  NAND2X1 U5352 ( .A(n1012), .B(n16692), .Y(n16710) );
  NAND2X1 U5353 ( .A(n1096), .B(n14802), .Y(n14820) );
  NAND2X1 U5354 ( .A(n1026), .B(n16377), .Y(n16395) );
  NAND2X1 U5355 ( .A(n956), .B(n17952), .Y(n17970) );
  NAND2X1 U5356 ( .A(n1110), .B(n14487), .Y(n14505) );
  NAND2X1 U5357 ( .A(n1040), .B(n16062), .Y(n16080) );
  NAND2X1 U5358 ( .A(n970), .B(n17637), .Y(n17655) );
  NAND2X1 U5359 ( .A(n1124), .B(n14172), .Y(n14190) );
  NAND2X1 U5360 ( .A(n1054), .B(n15747), .Y(n15765) );
  NAND2X1 U5361 ( .A(n984), .B(n17322), .Y(n17340) );
  NAND2X1 U5362 ( .A(n586), .B(n2892), .Y(n10074) );
  NAND2X1 U5363 ( .A(n587), .B(n2661), .Y(n11242) );
  NAND2X1 U5364 ( .A(n588), .B(n3252), .Y(n8322) );
  NAND2X1 U5365 ( .A(n589), .B(n2710), .Y(n10950) );
  NAND2X1 U5366 ( .A(n591), .B(n3432), .Y(n7446) );
  NAND2X1 U5367 ( .A(n590), .B(n3083), .Y(n9198) );
  NAND2X1 U5368 ( .A(n592), .B(n2832), .Y(n10366) );
  NAND2X1 U5369 ( .A(n593), .B(n3014), .Y(n9490) );
  NAND2X1 U5370 ( .A(n594), .B(n3191), .Y(n8614) );
  NAND2X1 U5371 ( .A(n595), .B(n3374), .Y(n7738) );
  NAND2X1 U5372 ( .A(n596), .B(n2589), .Y(n11534) );
  NAND2X1 U5373 ( .A(n597), .B(n2771), .Y(n10658) );
  NAND2X1 U5374 ( .A(n598), .B(n2953), .Y(n9782) );
  NAND2X1 U5375 ( .A(n599), .B(n3133), .Y(n8906) );
  NAND2X1 U5376 ( .A(n600), .B(n3313), .Y(n8030) );
  NAND2X1 U5377 ( .A(n585), .B(n3494), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n260) );
  CLKINVX3 U5378 ( .A(n9914), .Y(n5336) );
  CLKINVX3 U5379 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n98), .Y(n6132) );
  CLKINVX3 U5380 ( .A(n8162), .Y(n5808) );
  CLKINVX3 U5381 ( .A(n11082), .Y(n4982) );
  CLKINVX3 U5382 ( .A(n10790), .Y(n5066) );
  CLKINVX3 U5383 ( .A(n7286), .Y(n6036) );
  CLKINVX3 U5384 ( .A(n9038), .Y(n5572) );
  CLKINVX3 U5385 ( .A(n10206), .Y(n5252) );
  CLKINVX3 U5386 ( .A(n9330), .Y(n5496) );
  CLKINVX3 U5387 ( .A(n8454), .Y(n5724) );
  CLKINVX3 U5388 ( .A(n7578), .Y(n5960) );
  CLKINVX3 U5389 ( .A(n11374), .Y(n4866) );
  CLKINVX3 U5390 ( .A(n10498), .Y(n5174) );
  CLKINVX3 U5391 ( .A(n9622), .Y(n5420) );
  CLKINVX3 U5392 ( .A(n8746), .Y(n5648) );
  CLKINVX3 U5393 ( .A(n7870), .Y(n5884) );
  NAND2X1 U5394 ( .A(n1133), .B(n1141), .Y(n13854) );
  NAND2X1 U5395 ( .A(n994), .B(n1002), .Y(n17004) );
  NAND2X1 U5396 ( .A(n938), .B(n946), .Y(n18264) );
  NAND2X1 U5397 ( .A(n1078), .B(n1086), .Y(n15114) );
  NAND2X1 U5398 ( .A(n1064), .B(n1072), .Y(n15429) );
  NAND2X1 U5399 ( .A(n924), .B(n932), .Y(n18579) );
  NAND2X1 U5400 ( .A(n1008), .B(n1016), .Y(n16689) );
  NAND2X1 U5401 ( .A(n1092), .B(n1100), .Y(n14799) );
  NAND2X1 U5402 ( .A(n1022), .B(n1030), .Y(n16374) );
  NAND2X1 U5403 ( .A(n952), .B(n960), .Y(n17949) );
  NAND2X1 U5404 ( .A(n1106), .B(n1114), .Y(n14484) );
  NAND2X1 U5405 ( .A(n1036), .B(n1044), .Y(n16059) );
  NAND2X1 U5406 ( .A(n966), .B(n974), .Y(n17634) );
  NAND2X1 U5407 ( .A(n1120), .B(n1128), .Y(n14169) );
  NAND2X1 U5408 ( .A(n1050), .B(n1058), .Y(n15744) );
  NAND2X1 U5409 ( .A(n980), .B(n988), .Y(n17319) );
  NAND2X1 U5410 ( .A(n1172), .B(n6549), .Y(n13248) );
  NAND2X1 U5411 ( .A(n1212), .B(n6844), .Y(n12618) );
  NAND2X1 U5412 ( .A(n1218), .B(n6890), .Y(n12933) );
  AOI21XL U5413 ( .A0(n9970), .A1(n5362), .B0(n17235), .Y(n17045) );
  AOI21XL U5414 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .A1(n6130), 
        .B0(n14085), .Y(n13895) );
  AOI21XL U5415 ( .A0(n8218), .A1(n5834), .B0(n15345), .Y(n15155) );
  AOI21XL U5416 ( .A0(n11138), .A1(n5008), .B0(n18495), .Y(n18305) );
  AOI21XL U5417 ( .A0(n11430), .A1(n4892), .B0(n18810), .Y(n18620) );
  AOI21XL U5418 ( .A0(n8510), .A1(n5750), .B0(n15660), .Y(n15470) );
  AOI21XL U5419 ( .A0(n9678), .A1(n5446), .B0(n16920), .Y(n16730) );
  AOI21XL U5420 ( .A0(n7926), .A1(n5910), .B0(n15030), .Y(n14840) );
  AOI21XL U5421 ( .A0(n9386), .A1(n5522), .B0(n16605), .Y(n16415) );
  AOI21XL U5422 ( .A0(n10846), .A1(n5092), .B0(n18180), .Y(n17990) );
  AOI21XL U5423 ( .A0(n7634), .A1(n5986), .B0(n14715), .Y(n14525) );
  AOI21XL U5424 ( .A0(n9094), .A1(n5598), .B0(n16290), .Y(n16100) );
  AOI21XL U5425 ( .A0(n10554), .A1(n5200), .B0(n17865), .Y(n17675) );
  AOI21XL U5426 ( .A0(n7342), .A1(n6062), .B0(n14400), .Y(n14210) );
  AOI21XL U5427 ( .A0(n8802), .A1(n5674), .B0(n15975), .Y(n15785) );
  AOI21XL U5428 ( .A0(n10262), .A1(n5278), .B0(n17550), .Y(n17360) );
  NAND3X1 U5429 ( .A(n2867), .B(n2872), .C(n370), .Y(n17163) );
  NAND3X1 U5430 ( .A(n3468), .B(n3473), .C(n369), .Y(n14013) );
  NAND3X1 U5431 ( .A(n2625), .B(n2630), .C(n371), .Y(n18423) );
  NAND3X1 U5432 ( .A(n3227), .B(n3232), .C(n372), .Y(n15273) );
  NAND3X1 U5433 ( .A(n3166), .B(n3171), .C(n373), .Y(n15588) );
  NAND3X1 U5434 ( .A(n2928), .B(n2933), .C(n375), .Y(n16848) );
  NAND3X1 U5435 ( .A(n2564), .B(n2569), .C(n374), .Y(n18738) );
  NAND3X1 U5436 ( .A(n3288), .B(n3293), .C(n376), .Y(n14958) );
  NAND3X1 U5437 ( .A(n2989), .B(n2994), .C(n377), .Y(n16533) );
  NAND3X1 U5438 ( .A(n2686), .B(n2691), .C(n378), .Y(n18108) );
  NAND3X1 U5439 ( .A(n3349), .B(n3354), .C(n379), .Y(n14643) );
  NAND3X1 U5440 ( .A(n3047), .B(n3052), .C(n380), .Y(n16218) );
  NAND3X1 U5441 ( .A(n2746), .B(n2751), .C(n381), .Y(n17793) );
  NAND3X1 U5442 ( .A(n3407), .B(n3412), .C(n382), .Y(n14328) );
  NAND3X1 U5443 ( .A(n3108), .B(n3113), .C(n383), .Y(n15903) );
  NAND3X1 U5444 ( .A(n2807), .B(n2812), .C(n384), .Y(n17478) );
  CLKINVX3 U5445 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n171), .Y(n6105) );
  CLKINVX3 U5446 ( .A(n9985), .Y(n5321) );
  CLKINVX3 U5447 ( .A(n11153), .Y(n4967) );
  CLKINVX3 U5448 ( .A(n8233), .Y(n5793) );
  CLKINVX3 U5449 ( .A(n10861), .Y(n5051) );
  CLKINVX3 U5450 ( .A(n9109), .Y(n5557) );
  CLKINVX3 U5451 ( .A(n7357), .Y(n6021) );
  CLKINVX3 U5452 ( .A(n10277), .Y(n5237) );
  CLKINVX3 U5453 ( .A(n9401), .Y(n5481) );
  CLKINVX3 U5454 ( .A(n8525), .Y(n5709) );
  CLKINVX3 U5455 ( .A(n7649), .Y(n5945) );
  CLKINVX3 U5456 ( .A(n11445), .Y(n4851) );
  CLKINVX3 U5457 ( .A(n10569), .Y(n5159) );
  CLKINVX3 U5458 ( .A(n9693), .Y(n5405) );
  CLKINVX3 U5459 ( .A(n8817), .Y(n5633) );
  CLKINVX3 U5460 ( .A(n7941), .Y(n5869) );
  NOR2X1 U5461 ( .A(n562), .B(n5350), .Y(n10003) );
  NOR2X1 U5462 ( .A(n561), .B(n6146), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n189) );
  NOR2X1 U5463 ( .A(n563), .B(n4996), .Y(n11171) );
  NOR2X1 U5464 ( .A(n564), .B(n5822), .Y(n8251) );
  NOR2X1 U5465 ( .A(n565), .B(n5080), .Y(n10879) );
  NOR2X1 U5466 ( .A(n567), .B(n6050), .Y(n7375) );
  NOR2X1 U5467 ( .A(n566), .B(n5586), .Y(n9127) );
  NOR2X1 U5468 ( .A(n568), .B(n5266), .Y(n10295) );
  NOR2X1 U5469 ( .A(n569), .B(n5510), .Y(n9419) );
  NOR2X1 U5470 ( .A(n570), .B(n5738), .Y(n8543) );
  NOR2X1 U5471 ( .A(n571), .B(n5974), .Y(n7667) );
  NOR2X1 U5472 ( .A(n572), .B(n4880), .Y(n11463) );
  NOR2X1 U5473 ( .A(n573), .B(n5188), .Y(n10587) );
  NOR2X1 U5474 ( .A(n574), .B(n5434), .Y(n9711) );
  NOR2X1 U5475 ( .A(n575), .B(n5662), .Y(n8835) );
  NOR2X1 U5476 ( .A(n576), .B(n5898), .Y(n7959) );
  NAND3X1 U5477 ( .A(n1004), .B(n2857), .C(n5366), .Y(n9974) );
  NAND3X1 U5478 ( .A(n1145), .B(n3458), .C(n6156), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n160) );
  NAND3X1 U5479 ( .A(n948), .B(n2615), .C(n5012), .Y(n11142) );
  NAND3X1 U5480 ( .A(n1088), .B(n3217), .C(n5838), .Y(n8222) );
  NAND3X1 U5481 ( .A(n962), .B(n2676), .C(n5096), .Y(n10850) );
  NAND3X1 U5482 ( .A(n1046), .B(n3037), .C(n5602), .Y(n9098) );
  NAND3X1 U5483 ( .A(n1130), .B(n3397), .C(n6066), .Y(n7346) );
  NAND3X1 U5484 ( .A(n990), .B(n2797), .C(n5282), .Y(n10266) );
  NAND3X1 U5485 ( .A(n1032), .B(n2979), .C(n5526), .Y(n9390) );
  NAND3X1 U5486 ( .A(n1074), .B(n3156), .C(n5754), .Y(n8514) );
  NAND3X1 U5487 ( .A(n1116), .B(n3339), .C(n5990), .Y(n7638) );
  NAND3X1 U5488 ( .A(n934), .B(n2554), .C(n4896), .Y(n11434) );
  NAND3X1 U5489 ( .A(n976), .B(n2736), .C(n5204), .Y(n10558) );
  NAND3X1 U5490 ( .A(n1018), .B(n2918), .C(n5450), .Y(n9682) );
  NAND3X1 U5491 ( .A(n1060), .B(n3098), .C(n5678), .Y(n8806) );
  NAND3X1 U5492 ( .A(n1102), .B(n3278), .C(n5914), .Y(n7930) );
  NOR2XL U5493 ( .A(n1310), .B(n2876), .Y(n17059) );
  NOR2XL U5494 ( .A(n1280), .B(n3474), .Y(n13909) );
  NOR2XL U5495 ( .A(n1292), .B(n3237), .Y(n15169) );
  NOR2XL U5496 ( .A(n1322), .B(n2634), .Y(n18319) );
  NOR2XL U5497 ( .A(n1295), .B(n3176), .Y(n15484) );
  NOR2XL U5498 ( .A(n1307), .B(n2937), .Y(n16744) );
  NOR2XL U5499 ( .A(n1325), .B(n2573), .Y(n18634) );
  NOR2XL U5500 ( .A(n1289), .B(n3296), .Y(n14854) );
  NOR2XL U5501 ( .A(n1304), .B(n2998), .Y(n16429) );
  NOR2XL U5502 ( .A(n1319), .B(n2695), .Y(n18004) );
  NOR2XL U5503 ( .A(n1286), .B(n3359), .Y(n14539) );
  NOR2XL U5504 ( .A(n1301), .B(n3056), .Y(n16114) );
  NOR2XL U5505 ( .A(n1316), .B(n2756), .Y(n17689) );
  NOR2XL U5506 ( .A(n1283), .B(n3416), .Y(n14224) );
  NOR2XL U5507 ( .A(n1298), .B(n3117), .Y(n15799) );
  NOR2XL U5508 ( .A(n1313), .B(n2815), .Y(n17374) );
  CLKINVX3 U5509 ( .A(n17073), .Y(n5362) );
  CLKINVX3 U5510 ( .A(n13923), .Y(n6130) );
  CLKINVX3 U5511 ( .A(n18333), .Y(n5008) );
  CLKINVX3 U5512 ( .A(n15183), .Y(n5834) );
  CLKINVX3 U5513 ( .A(n15498), .Y(n5750) );
  CLKINVX3 U5514 ( .A(n16758), .Y(n5446) );
  CLKINVX3 U5515 ( .A(n14868), .Y(n5910) );
  CLKINVX3 U5516 ( .A(n18648), .Y(n4892) );
  CLKINVX3 U5517 ( .A(n16443), .Y(n5522) );
  CLKINVX3 U5518 ( .A(n18018), .Y(n5092) );
  CLKINVX3 U5519 ( .A(n14553), .Y(n5986) );
  CLKINVX3 U5520 ( .A(n16128), .Y(n5598) );
  CLKINVX3 U5521 ( .A(n17703), .Y(n5200) );
  CLKINVX3 U5522 ( .A(n14238), .Y(n6062) );
  CLKINVX3 U5523 ( .A(n15813), .Y(n5674) );
  CLKINVX3 U5524 ( .A(n17388), .Y(n5278) );
  INVX1 U5525 ( .A(n14085), .Y(n6153) );
  INVX1 U5526 ( .A(n17235), .Y(n5382) );
  INVX1 U5527 ( .A(n18495), .Y(n5028) );
  INVX1 U5528 ( .A(n15345), .Y(n5854) );
  INVX1 U5529 ( .A(n15660), .Y(n5770) );
  INVX1 U5530 ( .A(n16920), .Y(n5466) );
  INVX1 U5531 ( .A(n18810), .Y(n4912) );
  INVX1 U5532 ( .A(n15030), .Y(n5930) );
  INVX1 U5533 ( .A(n16605), .Y(n5542) );
  INVX1 U5534 ( .A(n18180), .Y(n5112) );
  INVX1 U5535 ( .A(n14715), .Y(n6006) );
  INVX1 U5536 ( .A(n16290), .Y(n5618) );
  INVX1 U5537 ( .A(n17865), .Y(n5220) );
  INVX1 U5538 ( .A(n14400), .Y(n6082) );
  INVX1 U5539 ( .A(n15975), .Y(n5694) );
  INVX1 U5540 ( .A(n17550), .Y(n5298) );
  AOI22XL U5541 ( .A0(n9996), .A1(n1246), .B0(n546), .B1(n401), .Y(n10078) );
  AOI22XL U5542 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n182), .A1(n1328), 
        .B0(n545), .B1(n402), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n264) );
  AOI22XL U5543 ( .A0(n11164), .A1(n1254), .B0(n547), .B1(n403), .Y(n11246) );
  AOI22XL U5544 ( .A0(n8244), .A1(n1234), .B0(n548), .B1(n404), .Y(n8326) );
  AOI22XL U5545 ( .A0(n10872), .A1(n1252), .B0(n549), .B1(n405), .Y(n10954) );
  AOI22XL U5546 ( .A0(n7368), .A1(n1228), .B0(n551), .B1(n407), .Y(n7450) );
  AOI22XL U5547 ( .A0(n9120), .A1(n1240), .B0(n550), .B1(n406), .Y(n9202) );
  AOI22XL U5548 ( .A0(n10288), .A1(n1248), .B0(n552), .B1(n408), .Y(n10370) );
  AOI22XL U5549 ( .A0(n9412), .A1(n1242), .B0(n553), .B1(n409), .Y(n9494) );
  AOI22XL U5550 ( .A0(n8536), .A1(n1236), .B0(n554), .B1(n410), .Y(n8618) );
  AOI22XL U5551 ( .A0(n7660), .A1(n1230), .B0(n555), .B1(n411), .Y(n7742) );
  AOI22XL U5552 ( .A0(n11456), .A1(n1256), .B0(n556), .B1(n412), .Y(n11538) );
  AOI22XL U5553 ( .A0(n10580), .A1(n1250), .B0(n557), .B1(n413), .Y(n10662) );
  AOI22XL U5554 ( .A0(n9704), .A1(n1244), .B0(n558), .B1(n414), .Y(n9786) );
  AOI22XL U5555 ( .A0(n8828), .A1(n1238), .B0(n559), .B1(n415), .Y(n8910) );
  AOI22XL U5556 ( .A0(n7952), .A1(n1232), .B0(n560), .B1(n416), .Y(n8034) );
  NAND2X1 U5557 ( .A(n5329), .B(n1005), .Y(n17041) );
  NAND2X1 U5558 ( .A(n6113), .B(n1144), .Y(n13891) );
  NAND2X1 U5559 ( .A(n4975), .B(n949), .Y(n18301) );
  NAND2X1 U5560 ( .A(n5801), .B(n1089), .Y(n15151) );
  NAND2X1 U5561 ( .A(n5717), .B(n1075), .Y(n15466) );
  NAND2X1 U5562 ( .A(n5413), .B(n1019), .Y(n16726) );
  NAND2X1 U5563 ( .A(n4859), .B(n935), .Y(n18616) );
  NAND2X1 U5564 ( .A(n5877), .B(n1103), .Y(n14836) );
  NAND2X1 U5565 ( .A(n5489), .B(n1033), .Y(n16411) );
  NAND2X1 U5566 ( .A(n5059), .B(n963), .Y(n17986) );
  NAND2X1 U5567 ( .A(n5953), .B(n1117), .Y(n14521) );
  NAND2X1 U5568 ( .A(n5565), .B(n1047), .Y(n16096) );
  NAND2X1 U5569 ( .A(n5167), .B(n977), .Y(n17671) );
  NAND2X1 U5570 ( .A(n6029), .B(n1131), .Y(n14206) );
  NAND2X1 U5571 ( .A(n5641), .B(n1061), .Y(n15781) );
  NAND2X1 U5572 ( .A(n5245), .B(n991), .Y(n17356) );
  NAND2X1 U5573 ( .A(n6549), .B(n1173), .Y(n13302) );
  NAND2X1 U5574 ( .A(n6844), .B(n1213), .Y(n12672) );
  NAND2X1 U5575 ( .A(n6890), .B(n1219), .Y(n12987) );
  AOI22X1 U5576 ( .A0(n513), .A1(n5350), .B0(n5366), .B1(n2883), .Y(n10097) );
  AOI22X1 U5577 ( .A0(n514), .A1(n6146), .B0(n6156), .B1(n3484), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n283) );
  AOI22X1 U5578 ( .A0(n516), .A1(n5822), .B0(n5838), .B1(n3247), .Y(n8345) );
  AOI22X1 U5579 ( .A0(n515), .A1(n4996), .B0(n5012), .B1(n2641), .Y(n11265) );
  AOI22X1 U5580 ( .A0(n522), .A1(n5080), .B0(n5096), .B1(n2708), .Y(n10973) );
  AOI22X1 U5581 ( .A0(n526), .A1(n6050), .B0(n6066), .B1(n3423), .Y(n7469) );
  AOI22X1 U5582 ( .A0(n524), .A1(n5586), .B0(n5602), .B1(n3063), .Y(n9221) );
  AOI22X1 U5583 ( .A0(n528), .A1(n5266), .B0(n5282), .B1(n2823), .Y(n10389) );
  AOI22X1 U5584 ( .A0(n521), .A1(n5510), .B0(n5526), .B1(n3009), .Y(n9513) );
  AOI22X1 U5585 ( .A0(n517), .A1(n5738), .B0(n5754), .B1(n3188), .Y(n8637) );
  AOI22X1 U5586 ( .A0(n523), .A1(n5974), .B0(n5990), .B1(n3371), .Y(n7761) );
  AOI22X1 U5587 ( .A0(n518), .A1(n4880), .B0(n4896), .B1(n2586), .Y(n11557) );
  AOI22X1 U5588 ( .A0(n525), .A1(n5188), .B0(n5204), .B1(n2768), .Y(n10681) );
  AOI22X1 U5589 ( .A0(n519), .A1(n5434), .B0(n5450), .B1(n2944), .Y(n9805) );
  AOI22X1 U5590 ( .A0(n527), .A1(n5662), .B0(n5678), .B1(n3130), .Y(n8929) );
  AOI22X1 U5591 ( .A0(n520), .A1(n5898), .B0(n5914), .B1(n3308), .Y(n8053) );
  CLKINVX3 U5592 ( .A(n17014), .Y(n5357) );
  CLKINVX3 U5593 ( .A(n13864), .Y(n6125) );
  CLKINVX3 U5594 ( .A(n18274), .Y(n5003) );
  CLKINVX3 U5595 ( .A(n15124), .Y(n5829) );
  CLKINVX3 U5596 ( .A(n15439), .Y(n5745) );
  CLKINVX3 U5597 ( .A(n18589), .Y(n4887) );
  CLKINVX3 U5598 ( .A(n16699), .Y(n5441) );
  CLKINVX3 U5599 ( .A(n14809), .Y(n5905) );
  CLKINVX3 U5600 ( .A(n16384), .Y(n5517) );
  CLKINVX3 U5601 ( .A(n17959), .Y(n5087) );
  CLKINVX3 U5602 ( .A(n14494), .Y(n5981) );
  CLKINVX3 U5603 ( .A(n16069), .Y(n5593) );
  CLKINVX3 U5604 ( .A(n17644), .Y(n5195) );
  CLKINVX3 U5605 ( .A(n14179), .Y(n6057) );
  CLKINVX3 U5606 ( .A(n15754), .Y(n5669) );
  CLKINVX3 U5607 ( .A(n17329), .Y(n5273) );
  AND2X2 U5608 ( .A(n2885), .B(n2894), .Y(n401) );
  AND2X2 U5609 ( .A(n3486), .B(n3499), .Y(n402) );
  AND2X2 U5610 ( .A(n2649), .B(n2664), .Y(n403) );
  AND2X2 U5611 ( .A(n3246), .B(n3254), .Y(n404) );
  AND2X2 U5612 ( .A(n2708), .B(n2723), .Y(n405) );
  AND2X2 U5613 ( .A(n3071), .B(n3086), .Y(n406) );
  AND2X2 U5614 ( .A(n3431), .B(n3445), .Y(n407) );
  AND2X2 U5615 ( .A(n2831), .B(n2835), .Y(n408) );
  AND2X2 U5616 ( .A(n3008), .B(n3025), .Y(n409) );
  AND2X2 U5617 ( .A(n3188), .B(n3193), .Y(n410) );
  AND2X2 U5618 ( .A(n3371), .B(n3385), .Y(n411) );
  AND2X2 U5619 ( .A(n2586), .B(n2603), .Y(n412) );
  AND2X2 U5620 ( .A(n2768), .B(n2785), .Y(n413) );
  AND2X2 U5621 ( .A(n2952), .B(n2955), .Y(n414) );
  AND2X2 U5622 ( .A(n3130), .B(n3144), .Y(n415) );
  AND2X2 U5623 ( .A(n3307), .B(n3327), .Y(n416) );
  INVX1 U5624 ( .A(n16997), .Y(n5326) );
  INVX1 U5625 ( .A(n18257), .Y(n4972) );
  INVX1 U5626 ( .A(n15107), .Y(n5798) );
  INVX1 U5627 ( .A(n13847), .Y(n6108) );
  INVX1 U5628 ( .A(n15422), .Y(n5714) );
  INVX1 U5629 ( .A(n18572), .Y(n4856) );
  INVX1 U5630 ( .A(n16682), .Y(n5410) );
  INVX1 U5631 ( .A(n14792), .Y(n5874) );
  INVX1 U5632 ( .A(n16367), .Y(n5486) );
  INVX1 U5633 ( .A(n17942), .Y(n5056) );
  INVX1 U5634 ( .A(n14477), .Y(n5950) );
  INVX1 U5635 ( .A(n16052), .Y(n5562) );
  INVX1 U5636 ( .A(n17627), .Y(n5164) );
  INVX1 U5637 ( .A(n14162), .Y(n6026) );
  INVX1 U5638 ( .A(n15737), .Y(n5638) );
  INVX1 U5639 ( .A(n17312), .Y(n5242) );
  AOI22X1 U5640 ( .A0(n5350), .A1(n401), .B0(n450), .B1(n5341), .Y(n10061) );
  AOI22X1 U5641 ( .A0(n6146), .A1(n402), .B0(n449), .B1(n6137), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n247) );
  AOI22X1 U5642 ( .A0(n4996), .A1(n403), .B0(n451), .B1(n4987), .Y(n11229) );
  AOI22X1 U5643 ( .A0(n5822), .A1(n404), .B0(n452), .B1(n5813), .Y(n8309) );
  AOI22X1 U5644 ( .A0(n5080), .A1(n405), .B0(n458), .B1(n5071), .Y(n10937) );
  AOI22X1 U5645 ( .A0(n6050), .A1(n407), .B0(n462), .B1(n6041), .Y(n7433) );
  AOI22X1 U5646 ( .A0(n5586), .A1(n406), .B0(n460), .B1(n5577), .Y(n9185) );
  AOI22X1 U5647 ( .A0(n5266), .A1(n408), .B0(n464), .B1(n5257), .Y(n10353) );
  AOI22X1 U5648 ( .A0(n5510), .A1(n409), .B0(n457), .B1(n5501), .Y(n9477) );
  AOI22X1 U5649 ( .A0(n5738), .A1(n410), .B0(n453), .B1(n5729), .Y(n8601) );
  AOI22X1 U5650 ( .A0(n5974), .A1(n411), .B0(n459), .B1(n5965), .Y(n7725) );
  AOI22X1 U5651 ( .A0(n4880), .A1(n412), .B0(n454), .B1(n4871), .Y(n11521) );
  AOI22X1 U5652 ( .A0(n5188), .A1(n413), .B0(n461), .B1(n5179), .Y(n10645) );
  AOI22X1 U5653 ( .A0(n5434), .A1(n414), .B0(n455), .B1(n5425), .Y(n9769) );
  AOI22X1 U5654 ( .A0(n5662), .A1(n415), .B0(n463), .B1(n5653), .Y(n8893) );
  AOI22X1 U5655 ( .A0(n5898), .A1(n416), .B0(n456), .B1(n5889), .Y(n8017) );
  INVX1 U5656 ( .A(n13937), .Y(n6107) );
  INVX1 U5657 ( .A(n17087), .Y(n5325) );
  INVX1 U5658 ( .A(n18347), .Y(n4971) );
  INVX1 U5659 ( .A(n15197), .Y(n5797) );
  INVX1 U5660 ( .A(n15512), .Y(n5713) );
  INVX1 U5661 ( .A(n18662), .Y(n4855) );
  INVX1 U5662 ( .A(n16772), .Y(n5409) );
  INVX1 U5663 ( .A(n14882), .Y(n5873) );
  INVX1 U5664 ( .A(n16457), .Y(n5485) );
  INVX1 U5665 ( .A(n18032), .Y(n5055) );
  INVX1 U5666 ( .A(n14567), .Y(n5949) );
  INVX1 U5667 ( .A(n16142), .Y(n5561) );
  INVX1 U5668 ( .A(n17717), .Y(n5163) );
  INVX1 U5669 ( .A(n14252), .Y(n6025) );
  INVX1 U5670 ( .A(n15827), .Y(n5637) );
  INVX1 U5671 ( .A(n17402), .Y(n5241) );
  AOI22X1 U5672 ( .A0(n3493), .A1(n13848), .B0(n6125), .B1(n434), .Y(n13846)
         );
  AOI22X1 U5673 ( .A0(n2892), .A1(n16998), .B0(n5357), .B1(n433), .Y(n16996)
         );
  AOI22X1 U5674 ( .A0(n2659), .A1(n18258), .B0(n5003), .B1(n435), .Y(n18256)
         );
  AOI22X1 U5675 ( .A0(n3252), .A1(n15108), .B0(n5829), .B1(n436), .Y(n15106)
         );
  AOI22X1 U5676 ( .A0(n3191), .A1(n15423), .B0(n5745), .B1(n437), .Y(n15421)
         );
  AOI22X1 U5677 ( .A0(n2589), .A1(n18573), .B0(n4887), .B1(n439), .Y(n18571)
         );
  AOI22X1 U5678 ( .A0(n2953), .A1(n16683), .B0(n5441), .B1(n438), .Y(n16681)
         );
  AOI22X1 U5679 ( .A0(n3313), .A1(n14793), .B0(n5905), .B1(n440), .Y(n14791)
         );
  AOI22X1 U5680 ( .A0(n3014), .A1(n16368), .B0(n5517), .B1(n441), .Y(n16366)
         );
  AOI22X1 U5681 ( .A0(n2710), .A1(n17943), .B0(n5087), .B1(n442), .Y(n17941)
         );
  AOI22X1 U5682 ( .A0(n3374), .A1(n14478), .B0(n5981), .B1(n443), .Y(n14476)
         );
  AOI22X1 U5683 ( .A0(n3081), .A1(n16053), .B0(n5593), .B1(n444), .Y(n16051)
         );
  AOI22X1 U5684 ( .A0(n2771), .A1(n17628), .B0(n5195), .B1(n445), .Y(n17626)
         );
  AOI22X1 U5685 ( .A0(n3432), .A1(n14163), .B0(n6057), .B1(n446), .Y(n14161)
         );
  AOI22X1 U5686 ( .A0(n3133), .A1(n15738), .B0(n5669), .B1(n447), .Y(n15736)
         );
  AOI22X1 U5687 ( .A0(n2832), .A1(n17313), .B0(n5273), .B1(n448), .Y(n17311)
         );
  CLKINVX3 U5688 ( .A(n3491), .Y(n3481) );
  CLKINVX3 U5689 ( .A(n2890), .Y(n2880) );
  CLKINVX3 U5690 ( .A(n2645), .Y(n2638) );
  CLKINVX3 U5691 ( .A(n3244), .Y(n3240) );
  CLKINVX3 U5692 ( .A(n3183), .Y(n3179) );
  CLKINVX3 U5693 ( .A(n2581), .Y(n2577) );
  CLKINVX3 U5694 ( .A(n2948), .Y(n2941) );
  CLKINVX3 U5695 ( .A(n3305), .Y(n3301) );
  CLKINVX3 U5696 ( .A(n3006), .Y(n3002) );
  CLKINVX3 U5697 ( .A(n2703), .Y(n2699) );
  CLKINVX3 U5698 ( .A(n3366), .Y(n3362) );
  CLKINVX3 U5699 ( .A(n3067), .Y(n3060) );
  CLKINVX3 U5700 ( .A(n2763), .Y(n2759) );
  CLKINVX3 U5701 ( .A(n3427), .Y(n3420) );
  CLKINVX3 U5702 ( .A(n3125), .Y(n3121) );
  CLKINVX3 U5703 ( .A(n2827), .Y(n2820) );
  AND2X2 U5704 ( .A(n2880), .B(n2894), .Y(n417) );
  AND2X2 U5705 ( .A(n3481), .B(n3507), .Y(n418) );
  AND2X2 U5706 ( .A(n2638), .B(n2656), .Y(n419) );
  AND2X2 U5707 ( .A(n3240), .B(n3254), .Y(n420) );
  AND2X2 U5708 ( .A(n2699), .B(n2717), .Y(n421) );
  AND2X2 U5709 ( .A(n3060), .B(n3078), .Y(n422) );
  AND2X2 U5710 ( .A(n3420), .B(n3439), .Y(n423) );
  AND2X2 U5711 ( .A(n2820), .B(n2840), .Y(n424) );
  AND2X2 U5712 ( .A(n3002), .B(n3025), .Y(n425) );
  AND2X2 U5713 ( .A(n3179), .B(n3193), .Y(n426) );
  AND2X2 U5714 ( .A(n3362), .B(n3385), .Y(n427) );
  AND2X2 U5715 ( .A(n2577), .B(n2595), .Y(n428) );
  AND2X2 U5716 ( .A(n2759), .B(n2777), .Y(n429) );
  AND2X2 U5717 ( .A(n2941), .B(n2955), .Y(n430) );
  AND2X2 U5718 ( .A(n3121), .B(n3144), .Y(n431) );
  AND2X2 U5719 ( .A(n3301), .B(n3318), .Y(n432) );
  NOR2X1 U5720 ( .A(n5346), .B(n9903), .Y(n10014) );
  NOR2X1 U5721 ( .A(n6142), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n86), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n200) );
  NOR2X1 U5722 ( .A(n4992), .B(n11071), .Y(n11182) );
  NOR2X1 U5723 ( .A(n5818), .B(n8151), .Y(n8262) );
  NOR2X1 U5724 ( .A(n5076), .B(n10779), .Y(n10890) );
  NOR2X1 U5725 ( .A(n5582), .B(n9027), .Y(n9138) );
  NOR2X1 U5726 ( .A(n6046), .B(n7275), .Y(n7386) );
  NOR2X1 U5727 ( .A(n5262), .B(n10195), .Y(n10306) );
  NOR2X1 U5728 ( .A(n5506), .B(n9319), .Y(n9430) );
  NOR2X1 U5729 ( .A(n5734), .B(n8443), .Y(n8554) );
  NOR2X1 U5730 ( .A(n5970), .B(n7567), .Y(n7678) );
  NOR2X1 U5731 ( .A(n4876), .B(n11363), .Y(n11474) );
  NOR2X1 U5732 ( .A(n5184), .B(n10487), .Y(n10598) );
  NOR2X1 U5733 ( .A(n5430), .B(n9611), .Y(n9722) );
  NOR2X1 U5734 ( .A(n5658), .B(n8735), .Y(n8846) );
  NOR2X1 U5735 ( .A(n5894), .B(n7859), .Y(n7970) );
  NOR2XL U5736 ( .A(n10000), .B(n9926), .Y(n10109) );
  NOR2XL U5737 ( .A(n265), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n111), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n295) );
  NOR2XL U5738 ( .A(n264), .B(n8174), .Y(n8357) );
  NOR2XL U5739 ( .A(n11168), .B(n11094), .Y(n11277) );
  NOR2XL U5740 ( .A(n10876), .B(n10802), .Y(n10985) );
  NOR2XL U5741 ( .A(n7372), .B(n7298), .Y(n7481) );
  NOR2XL U5742 ( .A(n9124), .B(n9050), .Y(n9233) );
  NOR2XL U5743 ( .A(n10292), .B(n10218), .Y(n10401) );
  NOR2XL U5744 ( .A(n9416), .B(n9342), .Y(n9525) );
  NOR2XL U5745 ( .A(n8540), .B(n8466), .Y(n8649) );
  NOR2XL U5746 ( .A(n7664), .B(n7590), .Y(n7773) );
  NOR2XL U5747 ( .A(n11460), .B(n11386), .Y(n11569) );
  NOR2XL U5748 ( .A(n10584), .B(n10510), .Y(n10693) );
  NOR2XL U5749 ( .A(n9708), .B(n9634), .Y(n9817) );
  NOR2XL U5750 ( .A(n8832), .B(n8758), .Y(n8941) );
  NOR2XL U5751 ( .A(n7956), .B(n7882), .Y(n8065) );
  INVX1 U5752 ( .A(n17033), .Y(n5328) );
  INVX1 U5753 ( .A(n13883), .Y(n6112) );
  INVX1 U5754 ( .A(n18293), .Y(n4974) );
  INVX1 U5755 ( .A(n15143), .Y(n5800) );
  INVX1 U5756 ( .A(n15458), .Y(n5716) );
  INVX1 U5757 ( .A(n18608), .Y(n4858) );
  INVX1 U5758 ( .A(n16718), .Y(n5412) );
  INVX1 U5759 ( .A(n14828), .Y(n5876) );
  INVX1 U5760 ( .A(n16403), .Y(n5488) );
  INVX1 U5761 ( .A(n17978), .Y(n5058) );
  INVX1 U5762 ( .A(n14513), .Y(n5952) );
  INVX1 U5763 ( .A(n16088), .Y(n5564) );
  INVX1 U5764 ( .A(n17663), .Y(n5166) );
  INVX1 U5765 ( .A(n14198), .Y(n6028) );
  INVX1 U5766 ( .A(n15773), .Y(n5640) );
  INVX1 U5767 ( .A(n17348), .Y(n5244) );
  AOI2BB1X1 U5768 ( .A0N(n10003), .A1N(n2903), .B0(n10004), .Y(n10001) );
  AOI2BB1X1 U5769 ( .A0N(top_core_EC_ss_gen_tbox_0__sboxs_r_n189), .A1N(n3503), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n190), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n187) );
  AOI2BB1X1 U5770 ( .A0N(n11171), .A1N(n2651), .B0(n11172), .Y(n11169) );
  AOI2BB1X1 U5771 ( .A0N(n8251), .A1N(n3263), .B0(n8252), .Y(n8249) );
  AOI2BB1X1 U5772 ( .A0N(n10879), .A1N(n2711), .B0(n10880), .Y(n10877) );
  AOI2BB1X1 U5773 ( .A0N(n9127), .A1N(n3073), .B0(n9128), .Y(n9125) );
  AOI2BB1X1 U5774 ( .A0N(n7375), .A1N(n3433), .B0(n7376), .Y(n7373) );
  AOI2BB1X1 U5775 ( .A0N(n10295), .A1N(n2834), .B0(n10296), .Y(n10293) );
  AOI2BB1X1 U5776 ( .A0N(n9419), .A1N(n3016), .B0(n9420), .Y(n9417) );
  AOI2BB1X1 U5777 ( .A0N(n8543), .A1N(n3202), .B0(n8544), .Y(n8541) );
  AOI2BB1X1 U5778 ( .A0N(n7667), .A1N(n3376), .B0(n7668), .Y(n7665) );
  AOI2BB1X1 U5779 ( .A0N(n11463), .A1N(n2590), .B0(n11464), .Y(n11461) );
  AOI2BB1X1 U5780 ( .A0N(n10587), .A1N(n2773), .B0(n10588), .Y(n10585) );
  AOI2BB1X1 U5781 ( .A0N(n9711), .A1N(n2964), .B0(n9712), .Y(n9709) );
  AOI2BB1X1 U5782 ( .A0N(n8835), .A1N(n3135), .B0(n8836), .Y(n8833) );
  AOI2BB1X1 U5783 ( .A0N(n7959), .A1N(n3325), .B0(n7960), .Y(n7957) );
  CLKINVX3 U5784 ( .A(n2486), .Y(n2373) );
  CLKINVX3 U5785 ( .A(n2487), .Y(n2374) );
  CLKINVX3 U5786 ( .A(n2485), .Y(n2368) );
  CLKINVX3 U5787 ( .A(n2485), .Y(n2369) );
  CLKINVX3 U5788 ( .A(n2486), .Y(n2372) );
  CLKINVX3 U5789 ( .A(n2485), .Y(n2370) );
  CLKINVX3 U5790 ( .A(n2486), .Y(n2371) );
  CLKINVX3 U5791 ( .A(n2488), .Y(n2378) );
  CLKINVX3 U5792 ( .A(n2489), .Y(n2381) );
  CLKINVX3 U5793 ( .A(n2489), .Y(n2382) );
  CLKINVX3 U5794 ( .A(n2490), .Y(n2383) );
  CLKINVX3 U5795 ( .A(n2489), .Y(n2380) );
  CLKINVX3 U5796 ( .A(n2488), .Y(n2379) );
  CLKINVX3 U5797 ( .A(n2487), .Y(n2375) );
  CLKINVX3 U5798 ( .A(n2487), .Y(n2376) );
  CLKINVX3 U5799 ( .A(n2488), .Y(n2377) );
  CLKINVX3 U5800 ( .A(n2490), .Y(n2384) );
  CLKINVX3 U5801 ( .A(n2491), .Y(n2386) );
  CLKINVX3 U5802 ( .A(n2492), .Y(n2391) );
  CLKINVX3 U5803 ( .A(n2493), .Y(n2392) );
  CLKINVX3 U5804 ( .A(n2491), .Y(n2388) );
  CLKINVX3 U5805 ( .A(n2491), .Y(n2387) );
  CLKINVX3 U5806 ( .A(n2492), .Y(n2389) );
  CLKINVX3 U5807 ( .A(n2490), .Y(n2385) );
  CLKINVX3 U5808 ( .A(n2492), .Y(n2390) );
  CLKINVX3 U5809 ( .A(n2493), .Y(n2393) );
  CLKINVX3 U5810 ( .A(n2493), .Y(n2394) );
  NAND2XL U5811 ( .A(n9896), .B(n15), .Y(n10081) );
  NAND2XL U5812 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .B(n14), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n267) );
  NAND2XL U5813 ( .A(n8144), .B(n17), .Y(n8329) );
  NAND2XL U5814 ( .A(n11064), .B(n16), .Y(n11249) );
  NAND2XL U5815 ( .A(n10772), .B(n18), .Y(n10957) );
  NAND2XL U5816 ( .A(n7268), .B(n20), .Y(n7453) );
  NAND2XL U5817 ( .A(n9020), .B(n19), .Y(n9205) );
  NAND2XL U5818 ( .A(n10188), .B(n21), .Y(n10373) );
  NAND2XL U5819 ( .A(n9312), .B(n22), .Y(n9497) );
  NAND2XL U5820 ( .A(n8436), .B(n23), .Y(n8621) );
  NAND2XL U5821 ( .A(n7560), .B(n24), .Y(n7745) );
  NAND2XL U5822 ( .A(n11356), .B(n25), .Y(n11541) );
  NAND2XL U5823 ( .A(n10480), .B(n26), .Y(n10665) );
  NAND2XL U5824 ( .A(n9604), .B(n27), .Y(n9789) );
  NAND2XL U5825 ( .A(n8728), .B(n28), .Y(n8913) );
  NAND2XL U5826 ( .A(n7852), .B(n29), .Y(n8037) );
  CLKINVX3 U5827 ( .A(n2896), .Y(n2893) );
  CLKINVX3 U5828 ( .A(n3499), .Y(n3494) );
  CLKINVX3 U5829 ( .A(n2653), .Y(n2650) );
  CLKINVX3 U5830 ( .A(n3256), .Y(n3253) );
  CLKINVX3 U5831 ( .A(n3195), .Y(n3192) );
  CLKINVX3 U5832 ( .A(n2957), .Y(n2954) );
  CLKINVX3 U5833 ( .A(n3020), .Y(n3015) );
  CLKINVX3 U5834 ( .A(n2714), .Y(n2711) );
  CLKINVX3 U5835 ( .A(n3380), .Y(n3375) );
  CLKINVX3 U5836 ( .A(n3075), .Y(n3072) );
  CLKINVX3 U5837 ( .A(n2779), .Y(n2772) );
  CLKINVX3 U5838 ( .A(n3436), .Y(n3433) );
  CLKINVX3 U5839 ( .A(n3139), .Y(n3134) );
  CLKINVX3 U5840 ( .A(n2839), .Y(n2833) );
  CLKINVX3 U5841 ( .A(n3319), .Y(n3314) );
  AOI21XL U5842 ( .A0(n135), .A1(n513), .B0(n10012), .Y(n10008) );
  AOI21XL U5843 ( .A0(n136), .A1(n514), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n198), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n194) );
  AOI21XL U5844 ( .A0(n137), .A1(n515), .B0(n11180), .Y(n11176) );
  AOI21XL U5845 ( .A0(n138), .A1(n516), .B0(n8260), .Y(n8256) );
  AOI21XL U5846 ( .A0(n139), .A1(n522), .B0(n10888), .Y(n10884) );
  AOI21XL U5847 ( .A0(n140), .A1(n524), .B0(n9136), .Y(n9132) );
  AOI21XL U5848 ( .A0(n141), .A1(n526), .B0(n7384), .Y(n7380) );
  AOI21XL U5849 ( .A0(n142), .A1(n528), .B0(n10304), .Y(n10300) );
  AOI21XL U5850 ( .A0(n143), .A1(n521), .B0(n9428), .Y(n9424) );
  AOI21XL U5851 ( .A0(n144), .A1(n517), .B0(n8552), .Y(n8548) );
  AOI21XL U5852 ( .A0(n145), .A1(n523), .B0(n7676), .Y(n7672) );
  AOI21XL U5853 ( .A0(n146), .A1(n518), .B0(n11472), .Y(n11468) );
  AOI21XL U5854 ( .A0(n147), .A1(n525), .B0(n10596), .Y(n10592) );
  AOI21XL U5855 ( .A0(n148), .A1(n519), .B0(n9720), .Y(n9716) );
  AOI21XL U5856 ( .A0(n149), .A1(n527), .B0(n8844), .Y(n8840) );
  AOI21XL U5857 ( .A0(n150), .A1(n520), .B0(n7968), .Y(n7964) );
  INVX1 U5858 ( .A(n10041), .Y(n5392) );
  INVX1 U5859 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n227), .Y(n6176) );
  INVX1 U5860 ( .A(n11209), .Y(n5038) );
  INVX1 U5861 ( .A(n8289), .Y(n5864) );
  INVX1 U5862 ( .A(n10917), .Y(n5122) );
  INVX1 U5863 ( .A(n9165), .Y(n5628) );
  INVX1 U5864 ( .A(n7413), .Y(n6092) );
  INVX1 U5865 ( .A(n10333), .Y(n5308) );
  INVX1 U5866 ( .A(n9457), .Y(n5552) );
  INVX1 U5867 ( .A(n8581), .Y(n5780) );
  INVX1 U5868 ( .A(n7705), .Y(n6016) );
  INVX1 U5869 ( .A(n11501), .Y(n4922) );
  INVX1 U5870 ( .A(n10625), .Y(n5230) );
  INVX1 U5871 ( .A(n9749), .Y(n5476) );
  INVX1 U5872 ( .A(n8873), .Y(n5704) );
  INVX1 U5873 ( .A(n7997), .Y(n5940) );
  AOI21X1 U5874 ( .A0(n10113), .A1(n2851), .B0(n10114), .Y(n10089) );
  AOI21X1 U5875 ( .A0(n10115), .A1(n10116), .B0(n2852), .Y(n10114) );
  NAND4X1 U5876 ( .A(n10051), .B(n9958), .C(n10117), .D(n10118), .Y(n10113) );
  AOI21X1 U5877 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n299), .A1(n3452), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n300), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n275) );
  AOI21X1 U5878 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n301), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n302), .B0(n3453), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n300) );
  NAND4X1 U5879 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n237), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n143), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n303), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n304), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n299) );
  AOI21X1 U5880 ( .A0(n8361), .A1(n3211), .B0(n8362), .Y(n8337) );
  AOI21X1 U5881 ( .A0(n8363), .A1(n8364), .B0(n3212), .Y(n8362) );
  NAND4X1 U5882 ( .A(n8299), .B(n8206), .C(n8365), .D(n8366), .Y(n8361) );
  AOI21X1 U5883 ( .A0(n11281), .A1(n2609), .B0(n11282), .Y(n11257) );
  AOI21X1 U5884 ( .A0(n11283), .A1(n11284), .B0(n2610), .Y(n11282) );
  NAND4X1 U5885 ( .A(n11219), .B(n11126), .C(n11285), .D(n11286), .Y(n11281)
         );
  AOI21X1 U5886 ( .A0(n10989), .A1(n2670), .B0(n10990), .Y(n10965) );
  AOI21X1 U5887 ( .A0(n10991), .A1(n10992), .B0(n2671), .Y(n10990) );
  NAND4X1 U5888 ( .A(n10927), .B(n10834), .C(n10993), .D(n10994), .Y(n10989)
         );
  AOI21X1 U5889 ( .A0(n7485), .A1(n3391), .B0(n7486), .Y(n7461) );
  AOI21X1 U5890 ( .A0(n7487), .A1(n7488), .B0(n3392), .Y(n7486) );
  NAND4X1 U5891 ( .A(n7423), .B(n7330), .C(n7489), .D(n7490), .Y(n7485) );
  AOI21X1 U5892 ( .A0(n9237), .A1(n3031), .B0(n9238), .Y(n9213) );
  AOI21X1 U5893 ( .A0(n9239), .A1(n9240), .B0(n3032), .Y(n9238) );
  NAND4X1 U5894 ( .A(n9175), .B(n9082), .C(n9241), .D(n9242), .Y(n9237) );
  AOI21X1 U5895 ( .A0(n10405), .A1(n2791), .B0(n10406), .Y(n10381) );
  AOI21X1 U5896 ( .A0(n10407), .A1(n10408), .B0(n2792), .Y(n10406) );
  NAND4X1 U5897 ( .A(n10343), .B(n10250), .C(n10409), .D(n10410), .Y(n10405)
         );
  AOI21X1 U5898 ( .A0(n9529), .A1(n2973), .B0(n9530), .Y(n9505) );
  AOI21X1 U5899 ( .A0(n9531), .A1(n9532), .B0(n2974), .Y(n9530) );
  NAND4X1 U5900 ( .A(n9467), .B(n9374), .C(n9533), .D(n9534), .Y(n9529) );
  AOI21X1 U5901 ( .A0(n8653), .A1(n3150), .B0(n8654), .Y(n8629) );
  AOI21X1 U5902 ( .A0(n8655), .A1(n8656), .B0(n3151), .Y(n8654) );
  NAND4X1 U5903 ( .A(n8591), .B(n8498), .C(n8657), .D(n8658), .Y(n8653) );
  AOI21X1 U5904 ( .A0(n7777), .A1(n3333), .B0(n7778), .Y(n7753) );
  AOI21X1 U5905 ( .A0(n7779), .A1(n7780), .B0(n3334), .Y(n7778) );
  NAND4X1 U5906 ( .A(n7715), .B(n7622), .C(n7781), .D(n7782), .Y(n7777) );
  AOI21X1 U5907 ( .A0(n11573), .A1(n2548), .B0(n11574), .Y(n11549) );
  AOI21X1 U5908 ( .A0(n11575), .A1(n11576), .B0(n2549), .Y(n11574) );
  NAND4X1 U5909 ( .A(n11511), .B(n11418), .C(n11577), .D(n11578), .Y(n11573)
         );
  AOI21X1 U5910 ( .A0(n10697), .A1(n2730), .B0(n10698), .Y(n10673) );
  AOI21X1 U5911 ( .A0(n10699), .A1(n10700), .B0(n2731), .Y(n10698) );
  NAND4X1 U5912 ( .A(n10635), .B(n10542), .C(n10701), .D(n10702), .Y(n10697)
         );
  AOI21X1 U5913 ( .A0(n9821), .A1(n2912), .B0(n9822), .Y(n9797) );
  AOI21X1 U5914 ( .A0(n9823), .A1(n9824), .B0(n2913), .Y(n9822) );
  NAND4X1 U5915 ( .A(n9759), .B(n9666), .C(n9825), .D(n9826), .Y(n9821) );
  AOI21X1 U5916 ( .A0(n8945), .A1(n3092), .B0(n8946), .Y(n8921) );
  AOI21X1 U5917 ( .A0(n8947), .A1(n8948), .B0(n3093), .Y(n8946) );
  NAND4X1 U5918 ( .A(n8883), .B(n8790), .C(n8949), .D(n8950), .Y(n8945) );
  AOI21X1 U5919 ( .A0(n8069), .A1(n3272), .B0(n8070), .Y(n8045) );
  AOI21X1 U5920 ( .A0(n8071), .A1(n8072), .B0(n3273), .Y(n8070) );
  NAND4X1 U5921 ( .A(n8007), .B(n7914), .C(n8073), .D(n8074), .Y(n8069) );
  CLKINVX3 U5922 ( .A(n17162), .Y(n5378) );
  CLKINVX3 U5923 ( .A(n14012), .Y(n6149) );
  CLKINVX3 U5924 ( .A(n15272), .Y(n5850) );
  CLKINVX3 U5925 ( .A(n18422), .Y(n5024) );
  CLKINVX3 U5926 ( .A(n15587), .Y(n5766) );
  CLKINVX3 U5927 ( .A(n16847), .Y(n5462) );
  CLKINVX3 U5928 ( .A(n18737), .Y(n4908) );
  CLKINVX3 U5929 ( .A(n14957), .Y(n5926) );
  CLKINVX3 U5930 ( .A(n16532), .Y(n5538) );
  CLKINVX3 U5931 ( .A(n18107), .Y(n5108) );
  CLKINVX3 U5932 ( .A(n14642), .Y(n6002) );
  CLKINVX3 U5933 ( .A(n16217), .Y(n5614) );
  CLKINVX3 U5934 ( .A(n17792), .Y(n5216) );
  CLKINVX3 U5935 ( .A(n14327), .Y(n6078) );
  CLKINVX3 U5936 ( .A(n15902), .Y(n5690) );
  CLKINVX3 U5937 ( .A(n17477), .Y(n5294) );
  NAND4BXL U5938 ( .AN(n17173), .B(n17004), .C(n17155), .D(n17164), .Y(n17171)
         );
  NAND4BXL U5939 ( .AN(n14023), .B(n13854), .C(n14005), .D(n14014), .Y(n14021)
         );
  NAND4BXL U5940 ( .AN(n18433), .B(n18264), .C(n18415), .D(n18424), .Y(n18431)
         );
  NAND4BXL U5941 ( .AN(n15283), .B(n15114), .C(n15265), .D(n15274), .Y(n15281)
         );
  NAND4BXL U5942 ( .AN(n15598), .B(n15429), .C(n15580), .D(n15589), .Y(n15596)
         );
  NAND4BXL U5943 ( .AN(n18748), .B(n18579), .C(n18730), .D(n18739), .Y(n18746)
         );
  NAND4BXL U5944 ( .AN(n16858), .B(n16689), .C(n16840), .D(n16849), .Y(n16856)
         );
  NAND4BXL U5945 ( .AN(n14968), .B(n14799), .C(n14950), .D(n14959), .Y(n14966)
         );
  NAND4BXL U5946 ( .AN(n16543), .B(n16374), .C(n16525), .D(n16534), .Y(n16541)
         );
  NAND4BXL U5947 ( .AN(n18118), .B(n17949), .C(n18100), .D(n18109), .Y(n18116)
         );
  NAND4BXL U5948 ( .AN(n14653), .B(n14484), .C(n14635), .D(n14644), .Y(n14651)
         );
  NAND4BXL U5949 ( .AN(n16228), .B(n16059), .C(n16210), .D(n16219), .Y(n16226)
         );
  NAND4BXL U5950 ( .AN(n17803), .B(n17634), .C(n17785), .D(n17794), .Y(n17801)
         );
  NAND4BXL U5951 ( .AN(n14338), .B(n14169), .C(n14320), .D(n14329), .Y(n14336)
         );
  NAND4BXL U5952 ( .AN(n15913), .B(n15744), .C(n15895), .D(n15904), .Y(n15911)
         );
  NAND4BXL U5953 ( .AN(n17488), .B(n17319), .C(n17470), .D(n17479), .Y(n17486)
         );
  CLKINVX3 U5954 ( .A(n3459), .Y(n3452) );
  CLKINVX3 U5955 ( .A(top_core_EC_ss_in[85]), .Y(n2851) );
  CLKINVX3 U5956 ( .A(top_core_EC_ss_in[117]), .Y(n2609) );
  CLKINVX3 U5957 ( .A(top_core_EC_ss_in[37]), .Y(n3211) );
  CLKINVX3 U5958 ( .A(top_core_EC_ss_in[69]), .Y(n2973) );
  CLKINVX3 U5959 ( .A(top_core_EC_ss_in[109]), .Y(n2670) );
  CLKINVX3 U5960 ( .A(top_core_EC_ss_in[45]), .Y(n3150) );
  CLKINVX3 U5961 ( .A(top_core_EC_ss_in[21]), .Y(n3333) );
  CLKINVX3 U5962 ( .A(top_core_EC_ss_in[61]), .Y(n3031) );
  CLKINVX3 U5963 ( .A(top_core_EC_ss_in[125]), .Y(n2548) );
  CLKINVX3 U5964 ( .A(top_core_EC_ss_in[101]), .Y(n2730) );
  CLKINVX3 U5965 ( .A(top_core_EC_ss_in[13]), .Y(n3391) );
  CLKINVX3 U5966 ( .A(top_core_EC_ss_in[77]), .Y(n2912) );
  CLKINVX3 U5967 ( .A(top_core_EC_ss_in[53]), .Y(n3092) );
  CLKINVX3 U5968 ( .A(top_core_EC_ss_in[93]), .Y(n2791) );
  CLKINVX3 U5969 ( .A(top_core_EC_ss_in[29]), .Y(n3272) );
  CLKINVX3 U5970 ( .A(n2874), .Y(n2871) );
  CLKINVX3 U5971 ( .A(n3478), .Y(n3472) );
  CLKINVX3 U5972 ( .A(n2632), .Y(n2629) );
  CLKINVX3 U5973 ( .A(n3235), .Y(n3231) );
  CLKINVX3 U5974 ( .A(n3174), .Y(n3170) );
  CLKINVX3 U5975 ( .A(n2571), .Y(n2568) );
  CLKINVX3 U5976 ( .A(n2935), .Y(n2932) );
  CLKINVX3 U5977 ( .A(n2693), .Y(n2690) );
  CLKINVX3 U5978 ( .A(n3054), .Y(n3051) );
  CLKINVX3 U5979 ( .A(n3414), .Y(n3411) );
  CLKINVX3 U5980 ( .A(n2814), .Y(n2811) );
  CLKINVX3 U5981 ( .A(n2996), .Y(n2993) );
  CLKINVX3 U5982 ( .A(n3357), .Y(n3353) );
  CLKINVX3 U5983 ( .A(n2754), .Y(n2750) );
  CLKINVX3 U5984 ( .A(n3115), .Y(n3112) );
  CLKINVX3 U5985 ( .A(n3295), .Y(n3292) );
  CLKINVX3 U5986 ( .A(n2858), .Y(n2853) );
  CLKINVX3 U5987 ( .A(top_core_EC_ss_in[5]), .Y(n3454) );
  CLKINVX3 U5988 ( .A(n2616), .Y(n2611) );
  CLKINVX3 U5989 ( .A(n3218), .Y(n3213) );
  CLKINVX3 U5990 ( .A(n2677), .Y(n2672) );
  CLKINVX3 U5991 ( .A(n3038), .Y(n3033) );
  CLKINVX3 U5992 ( .A(n3398), .Y(n3393) );
  CLKINVX3 U5993 ( .A(n2798), .Y(n2793) );
  CLKINVX3 U5994 ( .A(n2980), .Y(n2975) );
  CLKINVX3 U5995 ( .A(n3157), .Y(n3152) );
  CLKINVX3 U5996 ( .A(n3340), .Y(n3335) );
  CLKINVX3 U5997 ( .A(n2555), .Y(n2550) );
  CLKINVX3 U5998 ( .A(n2737), .Y(n2732) );
  CLKINVX3 U5999 ( .A(n2919), .Y(n2914) );
  CLKINVX3 U6000 ( .A(n3099), .Y(n3094) );
  CLKINVX3 U6001 ( .A(n3279), .Y(n3274) );
  INVX1 U6002 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n93), .Y(n6110) );
  INVX1 U6003 ( .A(n9909), .Y(n5323) );
  INVX1 U6004 ( .A(n11077), .Y(n4969) );
  INVX1 U6005 ( .A(n8157), .Y(n5795) );
  INVX1 U6006 ( .A(n10785), .Y(n5053) );
  INVX1 U6007 ( .A(n9033), .Y(n5559) );
  INVX1 U6008 ( .A(n7281), .Y(n6023) );
  INVX1 U6009 ( .A(n10201), .Y(n5239) );
  INVX1 U6010 ( .A(n9325), .Y(n5483) );
  INVX1 U6011 ( .A(n8449), .Y(n5711) );
  INVX1 U6012 ( .A(n7573), .Y(n5947) );
  INVX1 U6013 ( .A(n11369), .Y(n4853) );
  INVX1 U6014 ( .A(n10493), .Y(n5161) );
  INVX1 U6015 ( .A(n9617), .Y(n5407) );
  INVX1 U6016 ( .A(n8741), .Y(n5635) );
  INVX1 U6017 ( .A(n7865), .Y(n5871) );
  AND2X2 U6018 ( .A(n2892), .B(n2886), .Y(n433) );
  AND2X2 U6019 ( .A(n3493), .B(n3491), .Y(n434) );
  AND2X2 U6020 ( .A(n2651), .B(n2645), .Y(n435) );
  AND2X2 U6021 ( .A(n3252), .B(n3248), .Y(n436) );
  AND2X2 U6022 ( .A(n3191), .B(n3185), .Y(n437) );
  AND2X2 U6023 ( .A(n2953), .B(n2947), .Y(n438) );
  AND2X2 U6024 ( .A(n2589), .B(n2583), .Y(n439) );
  AND2X2 U6025 ( .A(n3313), .B(n3309), .Y(n440) );
  AND2X2 U6026 ( .A(n3014), .B(n3010), .Y(n441) );
  AND2X2 U6027 ( .A(n2710), .B(n2705), .Y(n442) );
  AND2X2 U6028 ( .A(n3374), .B(n3368), .Y(n443) );
  AND2X2 U6029 ( .A(n3073), .B(n3065), .Y(n444) );
  AND2X2 U6030 ( .A(n2771), .B(n2765), .Y(n445) );
  AND2X2 U6031 ( .A(n3432), .B(n3427), .Y(n446) );
  AND2X2 U6032 ( .A(n3133), .B(n3127), .Y(n447) );
  AND2X2 U6033 ( .A(n2832), .B(n2825), .Y(n448) );
  CLKINVX3 U6034 ( .A(n3476), .Y(n3473) );
  CLKINVX3 U6035 ( .A(n2873), .Y(n2872) );
  CLKINVX3 U6036 ( .A(n2631), .Y(n2630) );
  CLKINVX3 U6037 ( .A(n3233), .Y(n3232) );
  CLKINVX3 U6038 ( .A(n3172), .Y(n3171) );
  CLKINVX3 U6039 ( .A(n2938), .Y(n2933) );
  CLKINVX3 U6040 ( .A(n2570), .Y(n2569) );
  CLKINVX3 U6041 ( .A(n2999), .Y(n2994) );
  CLKINVX3 U6042 ( .A(n2696), .Y(n2691) );
  CLKINVX3 U6043 ( .A(n3355), .Y(n3354) );
  CLKINVX3 U6044 ( .A(n3053), .Y(n3052) );
  CLKINVX3 U6045 ( .A(n2752), .Y(n2751) );
  CLKINVX3 U6046 ( .A(n3417), .Y(n3412) );
  CLKINVX3 U6047 ( .A(n3114), .Y(n3113) );
  CLKINVX3 U6048 ( .A(n3298), .Y(n3293) );
  CLKINVX3 U6049 ( .A(n2817), .Y(n2812) );
  CLKINVX3 U6050 ( .A(n3491), .Y(n3483) );
  CLKINVX3 U6051 ( .A(n2885), .Y(n2882) );
  CLKINVX3 U6052 ( .A(n2646), .Y(n2640) );
  CLKINVX3 U6053 ( .A(n3251), .Y(n3242) );
  CLKINVX3 U6054 ( .A(n3190), .Y(n3181) );
  CLKINVX3 U6055 ( .A(n2588), .Y(n2579) );
  CLKINVX3 U6056 ( .A(n2949), .Y(n2943) );
  CLKINVX3 U6057 ( .A(n3013), .Y(n3004) );
  CLKINVX3 U6058 ( .A(n2709), .Y(n2701) );
  CLKINVX3 U6059 ( .A(n3373), .Y(n3364) );
  CLKINVX3 U6060 ( .A(n3068), .Y(n3062) );
  CLKINVX3 U6061 ( .A(n2770), .Y(n2761) );
  CLKINVX3 U6062 ( .A(n3428), .Y(n3422) );
  CLKINVX3 U6063 ( .A(n3132), .Y(n3123) );
  CLKINVX3 U6064 ( .A(n3312), .Y(n3303) );
  CLKINVX3 U6065 ( .A(n2828), .Y(n2822) );
  OAI21XL U6066 ( .A0(n5353), .A1(n997), .B0(n2898), .Y(n17071) );
  OAI21XL U6067 ( .A0(n6121), .A1(n1136), .B0(n3501), .Y(n13921) );
  OAI21XL U6068 ( .A0(n4999), .A1(n941), .B0(n2655), .Y(n18331) );
  OAI21XL U6069 ( .A0(n5825), .A1(n1081), .B0(n3258), .Y(n15181) );
  OAI21XL U6070 ( .A0(n5741), .A1(n1067), .B0(n3197), .Y(n15496) );
  OAI21XL U6071 ( .A0(n4883), .A1(n927), .B0(n2594), .Y(n18646) );
  OAI21XL U6072 ( .A0(n5437), .A1(n1011), .B0(n2959), .Y(n16756) );
  OAI21XL U6073 ( .A0(n5901), .A1(n1095), .B0(n3321), .Y(n14866) );
  OAI21XL U6074 ( .A0(n5513), .A1(n1025), .B0(n3022), .Y(n16441) );
  OAI21XL U6075 ( .A0(n5083), .A1(n955), .B0(n2716), .Y(n18016) );
  OAI21XL U6076 ( .A0(n5977), .A1(n1109), .B0(n3382), .Y(n14551) );
  OAI21XL U6077 ( .A0(n5589), .A1(n1039), .B0(n3077), .Y(n16126) );
  OAI21XL U6078 ( .A0(n5191), .A1(n969), .B0(n2775), .Y(n17701) );
  OAI21XL U6079 ( .A0(n6053), .A1(n1123), .B0(n3438), .Y(n14236) );
  OAI21XL U6080 ( .A0(n5665), .A1(n1053), .B0(n3141), .Y(n15811) );
  OAI21XL U6081 ( .A0(n5269), .A1(n983), .B0(n2841), .Y(n17386) );
  CLKINVX3 U6082 ( .A(n3459), .Y(n3453) );
  CLKINVX3 U6083 ( .A(n2858), .Y(n2852) );
  CLKINVX3 U6084 ( .A(n2616), .Y(n2610) );
  CLKINVX3 U6085 ( .A(n3218), .Y(n3212) );
  CLKINVX3 U6086 ( .A(n2980), .Y(n2974) );
  CLKINVX3 U6087 ( .A(n3157), .Y(n3151) );
  CLKINVX3 U6088 ( .A(n2677), .Y(n2671) );
  CLKINVX3 U6089 ( .A(n3340), .Y(n3334) );
  CLKINVX3 U6090 ( .A(n2555), .Y(n2549) );
  CLKINVX3 U6091 ( .A(n3038), .Y(n3032) );
  CLKINVX3 U6092 ( .A(n2737), .Y(n2731) );
  CLKINVX3 U6093 ( .A(n2919), .Y(n2913) );
  CLKINVX3 U6094 ( .A(n3398), .Y(n3392) );
  CLKINVX3 U6095 ( .A(n3099), .Y(n3093) );
  CLKINVX3 U6096 ( .A(n3279), .Y(n3273) );
  CLKINVX3 U6097 ( .A(n2798), .Y(n2792) );
  CLKINVX3 U6098 ( .A(n238), .Y(n3628) );
  CLKINVX3 U6099 ( .A(n617), .Y(n3636) );
  CLKINVX3 U6100 ( .A(n2234), .Y(n2227) );
  CLKINVX3 U6101 ( .A(n2234), .Y(n2226) );
  CLKINVX3 U6102 ( .A(n2233), .Y(n2225) );
  CLKINVX3 U6103 ( .A(n2230), .Y(n2224) );
  CLKINVX3 U6104 ( .A(n2235), .Y(n2223) );
  CLKINVX3 U6105 ( .A(n2233), .Y(n2222) );
  NAND4BXL U6106 ( .AN(n13849), .B(n14005), .C(n14114), .D(n14115), .Y(n14110)
         );
  AOI222X1 U6107 ( .A0(n466), .A1(n1136), .B0(n6151), .B1(n1142), .C0(n1133), 
        .C1(n418), .Y(n14115) );
  AOI2BB2X1 U6108 ( .B0(n6149), .B1(n3493), .A0N(n14073), .A1N(n402), .Y(
        n14114) );
  NAND4BXL U6109 ( .AN(n16999), .B(n17155), .C(n17264), .D(n17265), .Y(n17260)
         );
  AOI222X1 U6110 ( .A0(n465), .A1(n997), .B0(n5380), .B1(n1003), .C0(n994), 
        .C1(n417), .Y(n17265) );
  AOI2BB2X1 U6111 ( .B0(n5378), .B1(n2892), .A0N(n17223), .A1N(n401), .Y(
        n17264) );
  NAND4BXL U6112 ( .AN(n18259), .B(n18415), .C(n18524), .D(n18525), .Y(n18520)
         );
  AOI222X1 U6113 ( .A0(n467), .A1(n941), .B0(n5026), .B1(n947), .C0(n938), 
        .C1(n419), .Y(n18525) );
  AOI2BB2X1 U6114 ( .B0(n5024), .B1(n2660), .A0N(n18483), .A1N(n403), .Y(
        n18524) );
  NAND4BXL U6115 ( .AN(n15109), .B(n15265), .C(n15374), .D(n15375), .Y(n15370)
         );
  AOI222X1 U6116 ( .A0(n468), .A1(n1081), .B0(n5852), .B1(n1087), .C0(n1078), 
        .C1(n420), .Y(n15375) );
  AOI2BB2X1 U6117 ( .B0(n5850), .B1(n3252), .A0N(n15333), .A1N(n404), .Y(
        n15374) );
  NAND4BXL U6118 ( .AN(n15424), .B(n15580), .C(n15689), .D(n15690), .Y(n15685)
         );
  AOI222X1 U6119 ( .A0(n469), .A1(n1067), .B0(n5768), .B1(n1073), .C0(n1064), 
        .C1(n426), .Y(n15690) );
  AOI2BB2X1 U6120 ( .B0(n5766), .B1(n3191), .A0N(n15648), .A1N(n410), .Y(
        n15689) );
  NAND4BXL U6121 ( .AN(n18574), .B(n18730), .C(n18839), .D(n18840), .Y(n18835)
         );
  AOI222X1 U6122 ( .A0(n471), .A1(n927), .B0(n4910), .B1(n933), .C0(n924), 
        .C1(n428), .Y(n18840) );
  AOI2BB2X1 U6123 ( .B0(n4908), .B1(n2589), .A0N(n18798), .A1N(n412), .Y(
        n18839) );
  NAND4BXL U6124 ( .AN(n16684), .B(n16840), .C(n16949), .D(n16950), .Y(n16945)
         );
  AOI222X1 U6125 ( .A0(n470), .A1(n1011), .B0(n5464), .B1(n1017), .C0(n1008), 
        .C1(n430), .Y(n16950) );
  AOI2BB2X1 U6126 ( .B0(n5462), .B1(n2953), .A0N(n16908), .A1N(n414), .Y(
        n16949) );
  NAND4BXL U6127 ( .AN(n14794), .B(n14950), .C(n15059), .D(n15060), .Y(n15055)
         );
  AOI222X1 U6128 ( .A0(n472), .A1(n1095), .B0(n5928), .B1(n1101), .C0(n1092), 
        .C1(n432), .Y(n15060) );
  AOI2BB2X1 U6129 ( .B0(n5926), .B1(n3313), .A0N(n15018), .A1N(n416), .Y(
        n15059) );
  NAND4BXL U6130 ( .AN(n16369), .B(n16525), .C(n16634), .D(n16635), .Y(n16630)
         );
  AOI222X1 U6131 ( .A0(n473), .A1(n1025), .B0(n5540), .B1(n1031), .C0(n1022), 
        .C1(n425), .Y(n16635) );
  AOI2BB2X1 U6132 ( .B0(n5538), .B1(n3014), .A0N(n16593), .A1N(n409), .Y(
        n16634) );
  NAND4BXL U6133 ( .AN(n17944), .B(n18100), .C(n18209), .D(n18210), .Y(n18205)
         );
  AOI222X1 U6134 ( .A0(n474), .A1(n955), .B0(n5110), .B1(n961), .C0(n952), 
        .C1(n421), .Y(n18210) );
  AOI2BB2X1 U6135 ( .B0(n5108), .B1(n2710), .A0N(n18168), .A1N(n405), .Y(
        n18209) );
  NAND4BXL U6136 ( .AN(n14479), .B(n14635), .C(n14744), .D(n14745), .Y(n14740)
         );
  AOI222X1 U6137 ( .A0(n475), .A1(n1109), .B0(n6004), .B1(n1115), .C0(n1106), 
        .C1(n427), .Y(n14745) );
  AOI2BB2X1 U6138 ( .B0(n6002), .B1(n3374), .A0N(n14703), .A1N(n411), .Y(
        n14744) );
  NAND4BXL U6139 ( .AN(n16054), .B(n16210), .C(n16319), .D(n16320), .Y(n16315)
         );
  AOI222X1 U6140 ( .A0(n476), .A1(n1039), .B0(n5616), .B1(n1045), .C0(n1036), 
        .C1(n422), .Y(n16320) );
  AOI2BB2X1 U6141 ( .B0(n5614), .B1(n3082), .A0N(n16278), .A1N(n406), .Y(
        n16319) );
  NAND4BXL U6142 ( .AN(n17629), .B(n17785), .C(n17894), .D(n17895), .Y(n17890)
         );
  AOI222X1 U6143 ( .A0(n477), .A1(n969), .B0(n5218), .B1(n975), .C0(n966), 
        .C1(n429), .Y(n17895) );
  AOI2BB2X1 U6144 ( .B0(n5216), .B1(n2771), .A0N(n17853), .A1N(n413), .Y(
        n17894) );
  NAND4BXL U6145 ( .AN(n14164), .B(n14320), .C(n14429), .D(n14430), .Y(n14425)
         );
  AOI222X1 U6146 ( .A0(n478), .A1(n1123), .B0(n6080), .B1(n1129), .C0(n1120), 
        .C1(n423), .Y(n14430) );
  AOI2BB2X1 U6147 ( .B0(n6078), .B1(n3432), .A0N(n14388), .A1N(n407), .Y(
        n14429) );
  NAND4BXL U6148 ( .AN(n15739), .B(n15895), .C(n16004), .D(n16005), .Y(n16000)
         );
  AOI222X1 U6149 ( .A0(n479), .A1(n1053), .B0(n5692), .B1(n1059), .C0(n1050), 
        .C1(n431), .Y(n16005) );
  AOI2BB2X1 U6150 ( .B0(n5690), .B1(n3133), .A0N(n15963), .A1N(n415), .Y(
        n16004) );
  NAND4BXL U6151 ( .AN(n17314), .B(n17470), .C(n17579), .D(n17580), .Y(n17575)
         );
  AOI222X1 U6152 ( .A0(n480), .A1(n983), .B0(n5296), .B1(n989), .C0(n980), 
        .C1(n424), .Y(n17580) );
  AOI2BB2X1 U6153 ( .B0(n5294), .B1(n2832), .A0N(n17538), .A1N(n408), .Y(
        n17579) );
  CLKINVX3 U6154 ( .A(n767), .Y(n2347) );
  CLKINVX3 U6155 ( .A(n767), .Y(n2348) );
  CLKINVX3 U6156 ( .A(n767), .Y(n2349) );
  CLKINVX3 U6157 ( .A(n2354), .Y(n2350) );
  INVXL U6158 ( .A(n9896), .Y(n5347) );
  INVXL U6159 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .Y(n6143) );
  INVXL U6160 ( .A(n11064), .Y(n4993) );
  INVXL U6161 ( .A(n8144), .Y(n5819) );
  INVXL U6162 ( .A(n10772), .Y(n5077) );
  INVXL U6163 ( .A(n9020), .Y(n5583) );
  INVXL U6164 ( .A(n7268), .Y(n6047) );
  INVXL U6165 ( .A(n10188), .Y(n5263) );
  INVXL U6166 ( .A(n9312), .Y(n5507) );
  INVXL U6167 ( .A(n8436), .Y(n5735) );
  INVXL U6168 ( .A(n7560), .Y(n5971) );
  INVXL U6169 ( .A(n11356), .Y(n4877) );
  INVXL U6170 ( .A(n10480), .Y(n5185) );
  INVXL U6171 ( .A(n9604), .Y(n5431) );
  INVXL U6172 ( .A(n8728), .Y(n5659) );
  INVXL U6173 ( .A(n7852), .Y(n5895) );
  BUFX3 U6174 ( .A(n602), .Y(n1174) );
  BUFX3 U6175 ( .A(n603), .Y(n1214) );
  BUFX3 U6176 ( .A(n609), .Y(n1179) );
  BUFX3 U6177 ( .A(n604), .Y(n1220) );
  BUFX3 U6178 ( .A(n6164), .Y(n1139) );
  INVXL U6179 ( .A(n14), .Y(n6164) );
  BUFX3 U6180 ( .A(n5374), .Y(n996) );
  INVXL U6181 ( .A(n15), .Y(n5374) );
  BUFX3 U6182 ( .A(n5020), .Y(n940) );
  INVXL U6183 ( .A(n16), .Y(n5020) );
  BUFX3 U6184 ( .A(n5846), .Y(n1080) );
  INVXL U6185 ( .A(n17), .Y(n5846) );
  BUFX3 U6186 ( .A(n5104), .Y(n954) );
  INVXL U6187 ( .A(n18), .Y(n5104) );
  BUFX3 U6188 ( .A(n5610), .Y(n1038) );
  INVXL U6189 ( .A(n19), .Y(n5610) );
  BUFX3 U6190 ( .A(n6074), .Y(n1122) );
  INVXL U6191 ( .A(n20), .Y(n6074) );
  BUFX3 U6192 ( .A(n5290), .Y(n982) );
  INVXL U6193 ( .A(n21), .Y(n5290) );
  BUFX3 U6194 ( .A(n5534), .Y(n1024) );
  INVXL U6195 ( .A(n22), .Y(n5534) );
  BUFX3 U6196 ( .A(n5762), .Y(n1066) );
  INVXL U6197 ( .A(n23), .Y(n5762) );
  BUFX3 U6198 ( .A(n5998), .Y(n1108) );
  INVXL U6199 ( .A(n24), .Y(n5998) );
  BUFX3 U6200 ( .A(n4904), .Y(n926) );
  INVXL U6201 ( .A(n25), .Y(n4904) );
  BUFX3 U6202 ( .A(n5212), .Y(n968) );
  INVXL U6203 ( .A(n26), .Y(n5212) );
  BUFX3 U6204 ( .A(n5458), .Y(n1010) );
  INVXL U6205 ( .A(n27), .Y(n5458) );
  BUFX3 U6206 ( .A(n5686), .Y(n1052) );
  INVXL U6207 ( .A(n28), .Y(n5686) );
  BUFX3 U6208 ( .A(n5922), .Y(n1094) );
  INVXL U6209 ( .A(n29), .Y(n5922) );
  XOR2X1 U6210 ( .A(top_core_EC_mc_n614), .B(top_core_EC_mc_n849), .Y(
        top_core_EC_mc_n848) );
  XOR2X1 U6211 ( .A(top_core_EC_mc_n593), .B(top_core_EC_mc_n702), .Y(
        top_core_EC_mc_n701) );
  XOR2X1 U6212 ( .A(top_core_EC_mc_n6), .B(top_core_EC_mc_n7), .Y(
        top_core_EC_mc_n5) );
  XOR2X1 U6213 ( .A(top_core_EC_mc_n607), .B(top_core_EC_mc_n776), .Y(
        top_core_EC_mc_n775) );
  XOR2X1 U6214 ( .A(top_core_EC_mc_n600), .B(top_core_EC_mc_n709), .Y(
        top_core_EC_mc_n708) );
  BUFX3 U6215 ( .A(n613), .Y(n1223) );
  BUFX3 U6216 ( .A(n614), .Y(n1217) );
  BUFX3 U6217 ( .A(n601), .Y(n1182) );
  BUFX3 U6218 ( .A(n615), .Y(n1177) );
  BUFX3 U6219 ( .A(n6140), .Y(n1135) );
  INVXL U6220 ( .A(n91), .Y(n6140) );
  BUFX3 U6221 ( .A(n5344), .Y(n993) );
  INVXL U6222 ( .A(n90), .Y(n5344) );
  BUFX3 U6223 ( .A(n4990), .Y(n937) );
  INVXL U6224 ( .A(n92), .Y(n4990) );
  BUFX3 U6225 ( .A(n5816), .Y(n1077) );
  INVXL U6226 ( .A(n93), .Y(n5816) );
  BUFX3 U6227 ( .A(n5074), .Y(n951) );
  INVXL U6228 ( .A(n94), .Y(n5074) );
  BUFX3 U6229 ( .A(n5580), .Y(n1035) );
  INVXL U6230 ( .A(n96), .Y(n5580) );
  BUFX3 U6231 ( .A(n6044), .Y(n1119) );
  INVXL U6232 ( .A(n95), .Y(n6044) );
  BUFX3 U6233 ( .A(n5260), .Y(n979) );
  INVXL U6234 ( .A(n97), .Y(n5260) );
  BUFX3 U6235 ( .A(n5504), .Y(n1021) );
  INVXL U6236 ( .A(n98), .Y(n5504) );
  BUFX3 U6237 ( .A(n5732), .Y(n1063) );
  INVXL U6238 ( .A(n99), .Y(n5732) );
  BUFX3 U6239 ( .A(n5968), .Y(n1105) );
  INVXL U6240 ( .A(n100), .Y(n5968) );
  BUFX3 U6241 ( .A(n4874), .Y(n923) );
  INVXL U6242 ( .A(n101), .Y(n4874) );
  BUFX3 U6243 ( .A(n5182), .Y(n965) );
  INVXL U6244 ( .A(n102), .Y(n5182) );
  BUFX3 U6245 ( .A(n5428), .Y(n1007) );
  INVXL U6246 ( .A(n103), .Y(n5428) );
  BUFX3 U6247 ( .A(n5656), .Y(n1049) );
  INVXL U6248 ( .A(n104), .Y(n5656) );
  BUFX3 U6249 ( .A(n5892), .Y(n1091) );
  INVXL U6250 ( .A(n105), .Y(n5892) );
  INVX1 U6251 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n178), .Y(n6109) );
  INVX1 U6252 ( .A(n9992), .Y(n5322) );
  INVX1 U6253 ( .A(n11160), .Y(n4968) );
  INVX1 U6254 ( .A(n8240), .Y(n5794) );
  INVX1 U6255 ( .A(n10868), .Y(n5052) );
  INVX1 U6256 ( .A(n7364), .Y(n6022) );
  INVX1 U6257 ( .A(n9116), .Y(n5558) );
  INVX1 U6258 ( .A(n10284), .Y(n5238) );
  INVX1 U6259 ( .A(n9408), .Y(n5482) );
  INVX1 U6260 ( .A(n8532), .Y(n5710) );
  INVX1 U6261 ( .A(n7656), .Y(n5946) );
  INVX1 U6262 ( .A(n11452), .Y(n4852) );
  INVX1 U6263 ( .A(n10576), .Y(n5160) );
  INVX1 U6264 ( .A(n9700), .Y(n5406) );
  INVX1 U6265 ( .A(n8824), .Y(n5634) );
  INVX1 U6266 ( .A(n7948), .Y(n5870) );
  BUFX3 U6267 ( .A(n6150), .Y(n1136) );
  INVXL U6268 ( .A(n58), .Y(n6150) );
  BUFX3 U6269 ( .A(n5379), .Y(n997) );
  INVXL U6270 ( .A(n57), .Y(n5379) );
  BUFX3 U6271 ( .A(n5025), .Y(n941) );
  INVXL U6272 ( .A(n59), .Y(n5025) );
  BUFX3 U6273 ( .A(n5851), .Y(n1081) );
  INVXL U6274 ( .A(n60), .Y(n5851) );
  BUFX3 U6275 ( .A(n5767), .Y(n1067) );
  INVXL U6276 ( .A(n61), .Y(n5767) );
  BUFX3 U6277 ( .A(n4909), .Y(n927) );
  INVXL U6278 ( .A(n63), .Y(n4909) );
  BUFX3 U6279 ( .A(n5463), .Y(n1011) );
  INVXL U6280 ( .A(n62), .Y(n5463) );
  BUFX3 U6281 ( .A(n5927), .Y(n1095) );
  INVXL U6282 ( .A(n64), .Y(n5927) );
  BUFX3 U6283 ( .A(n5539), .Y(n1025) );
  INVXL U6284 ( .A(n65), .Y(n5539) );
  BUFX3 U6285 ( .A(n5109), .Y(n955) );
  INVXL U6286 ( .A(n66), .Y(n5109) );
  BUFX3 U6287 ( .A(n6003), .Y(n1109) );
  INVXL U6288 ( .A(n67), .Y(n6003) );
  BUFX3 U6289 ( .A(n5615), .Y(n1039) );
  INVXL U6290 ( .A(n68), .Y(n5615) );
  BUFX3 U6291 ( .A(n5217), .Y(n969) );
  INVXL U6292 ( .A(n69), .Y(n5217) );
  BUFX3 U6293 ( .A(n6079), .Y(n1123) );
  INVXL U6294 ( .A(n70), .Y(n6079) );
  BUFX3 U6295 ( .A(n5691), .Y(n1053) );
  INVXL U6296 ( .A(n71), .Y(n5691) );
  BUFX3 U6297 ( .A(n5295), .Y(n983) );
  INVXL U6298 ( .A(n72), .Y(n5295) );
  XNOR2X1 U6299 ( .A(n3989), .B(n2367), .Y(top_core_EC_n1020) );
  INVX1 U6300 ( .A(n17230), .Y(n5327) );
  INVX1 U6301 ( .A(n14080), .Y(n6111) );
  INVX1 U6302 ( .A(n15340), .Y(n5799) );
  INVX1 U6303 ( .A(n18490), .Y(n4973) );
  INVX1 U6304 ( .A(n15655), .Y(n5715) );
  INVX1 U6305 ( .A(n16915), .Y(n5411) );
  INVX1 U6306 ( .A(n18805), .Y(n4857) );
  INVX1 U6307 ( .A(n15025), .Y(n5875) );
  INVX1 U6308 ( .A(n16600), .Y(n5487) );
  INVX1 U6309 ( .A(n18175), .Y(n5057) );
  INVX1 U6310 ( .A(n14710), .Y(n5951) );
  INVX1 U6311 ( .A(n16285), .Y(n5563) );
  INVX1 U6312 ( .A(n17860), .Y(n5165) );
  INVX1 U6313 ( .A(n14395), .Y(n6027) );
  INVX1 U6314 ( .A(n15970), .Y(n5639) );
  INVX1 U6315 ( .A(n17545), .Y(n5243) );
  AND2X2 U6316 ( .A(n3481), .B(n3497), .Y(n449) );
  AND2X2 U6317 ( .A(n2880), .B(n2894), .Y(n450) );
  AND2X2 U6318 ( .A(n2638), .B(n2654), .Y(n451) );
  AND2X2 U6319 ( .A(n3240), .B(n3254), .Y(n452) );
  AND2X2 U6320 ( .A(n3179), .B(n3193), .Y(n453) );
  AND2X2 U6321 ( .A(n2577), .B(n2593), .Y(n454) );
  AND2X2 U6322 ( .A(n2941), .B(n2955), .Y(n455) );
  AND2X2 U6323 ( .A(n3301), .B(n3318), .Y(n456) );
  AND2X2 U6324 ( .A(n3002), .B(n3020), .Y(n457) );
  AND2X2 U6325 ( .A(n2699), .B(n2715), .Y(n458) );
  AND2X2 U6326 ( .A(n3362), .B(n3380), .Y(n459) );
  AND2X2 U6327 ( .A(n3060), .B(n3076), .Y(n460) );
  AND2X2 U6328 ( .A(n2759), .B(n2777), .Y(n461) );
  AND2X2 U6329 ( .A(n3420), .B(n3437), .Y(n462) );
  AND2X2 U6330 ( .A(n3121), .B(n3139), .Y(n463) );
  AND2X2 U6331 ( .A(n2820), .B(n2836), .Y(n464) );
  INVX1 U6332 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n91), .Y(n6133) );
  INVX1 U6333 ( .A(n9907), .Y(n5337) );
  INVX1 U6334 ( .A(n11075), .Y(n4983) );
  INVX1 U6335 ( .A(n8155), .Y(n5809) );
  INVX1 U6336 ( .A(n10783), .Y(n5067) );
  INVX1 U6337 ( .A(n9031), .Y(n5573) );
  INVX1 U6338 ( .A(n7279), .Y(n6037) );
  INVX1 U6339 ( .A(n10199), .Y(n5253) );
  INVX1 U6340 ( .A(n9323), .Y(n5497) );
  INVX1 U6341 ( .A(n8447), .Y(n5725) );
  INVX1 U6342 ( .A(n7571), .Y(n5961) );
  INVX1 U6343 ( .A(n11367), .Y(n4867) );
  INVX1 U6344 ( .A(n10491), .Y(n5175) );
  INVX1 U6345 ( .A(n9615), .Y(n5421) );
  INVX1 U6346 ( .A(n8739), .Y(n5649) );
  INVX1 U6347 ( .A(n7863), .Y(n5885) );
  AOI31X1 U6348 ( .A0(n13854), .A1(n6153), .A2(n13855), .B0(n3454), .Y(n13853)
         );
  AOI21X1 U6349 ( .A0(n6130), .A1(n3481), .B0(n6148), .Y(n13855) );
  INVX1 U6350 ( .A(n13856), .Y(n6148) );
  AOI31X1 U6351 ( .A0(n17004), .A1(n5382), .A2(n17005), .B0(n2853), .Y(n17003)
         );
  AOI21X1 U6352 ( .A0(n5362), .A1(n2880), .B0(n5377), .Y(n17005) );
  INVX1 U6353 ( .A(n17006), .Y(n5377) );
  AOI31X1 U6354 ( .A0(n18264), .A1(n5028), .A2(n18265), .B0(n2611), .Y(n18263)
         );
  AOI21X1 U6355 ( .A0(n5008), .A1(n2638), .B0(n5023), .Y(n18265) );
  INVX1 U6356 ( .A(n18266), .Y(n5023) );
  AOI31X1 U6357 ( .A0(n15114), .A1(n5854), .A2(n15115), .B0(n3213), .Y(n15113)
         );
  AOI21X1 U6358 ( .A0(n5834), .A1(n3240), .B0(n5849), .Y(n15115) );
  INVX1 U6359 ( .A(n15116), .Y(n5849) );
  AOI31X1 U6360 ( .A0(n15429), .A1(n5770), .A2(n15430), .B0(n3152), .Y(n15428)
         );
  AOI21X1 U6361 ( .A0(n5750), .A1(n3179), .B0(n5765), .Y(n15430) );
  INVX1 U6362 ( .A(n15431), .Y(n5765) );
  AOI31X1 U6363 ( .A0(n18579), .A1(n4912), .A2(n18580), .B0(n2550), .Y(n18578)
         );
  AOI21X1 U6364 ( .A0(n4892), .A1(n2577), .B0(n4907), .Y(n18580) );
  INVX1 U6365 ( .A(n18581), .Y(n4907) );
  AOI31X1 U6366 ( .A0(n16689), .A1(n5466), .A2(n16690), .B0(n2914), .Y(n16688)
         );
  AOI21X1 U6367 ( .A0(n5446), .A1(n2941), .B0(n5461), .Y(n16690) );
  INVX1 U6368 ( .A(n16691), .Y(n5461) );
  AOI31X1 U6369 ( .A0(n14799), .A1(n5930), .A2(n14800), .B0(n3274), .Y(n14798)
         );
  AOI21X1 U6370 ( .A0(n5910), .A1(n3301), .B0(n5925), .Y(n14800) );
  INVX1 U6371 ( .A(n14801), .Y(n5925) );
  AOI31X1 U6372 ( .A0(n16374), .A1(n5542), .A2(n16375), .B0(n2975), .Y(n16373)
         );
  AOI21X1 U6373 ( .A0(n5522), .A1(n3002), .B0(n5537), .Y(n16375) );
  INVX1 U6374 ( .A(n16376), .Y(n5537) );
  AOI31X1 U6375 ( .A0(n17949), .A1(n5112), .A2(n17950), .B0(n2672), .Y(n17948)
         );
  AOI21X1 U6376 ( .A0(n5092), .A1(n2699), .B0(n5107), .Y(n17950) );
  INVX1 U6377 ( .A(n17951), .Y(n5107) );
  AOI31X1 U6378 ( .A0(n14484), .A1(n6006), .A2(n14485), .B0(n3335), .Y(n14483)
         );
  AOI21X1 U6379 ( .A0(n5986), .A1(n3362), .B0(n6001), .Y(n14485) );
  INVX1 U6380 ( .A(n14486), .Y(n6001) );
  AOI31X1 U6381 ( .A0(n16059), .A1(n5618), .A2(n16060), .B0(n3033), .Y(n16058)
         );
  AOI21X1 U6382 ( .A0(n5598), .A1(n3060), .B0(n5613), .Y(n16060) );
  INVX1 U6383 ( .A(n16061), .Y(n5613) );
  AOI31X1 U6384 ( .A0(n17634), .A1(n5220), .A2(n17635), .B0(n2732), .Y(n17633)
         );
  AOI21X1 U6385 ( .A0(n5200), .A1(n2759), .B0(n5215), .Y(n17635) );
  INVX1 U6386 ( .A(n17636), .Y(n5215) );
  AOI31X1 U6387 ( .A0(n14169), .A1(n6082), .A2(n14170), .B0(n3393), .Y(n14168)
         );
  AOI21X1 U6388 ( .A0(n6062), .A1(n3420), .B0(n6077), .Y(n14170) );
  INVX1 U6389 ( .A(n14171), .Y(n6077) );
  AOI31X1 U6390 ( .A0(n15744), .A1(n5694), .A2(n15745), .B0(n3094), .Y(n15743)
         );
  AOI21X1 U6391 ( .A0(n5674), .A1(n3121), .B0(n5689), .Y(n15745) );
  INVX1 U6392 ( .A(n15746), .Y(n5689) );
  AOI31X1 U6393 ( .A0(n17319), .A1(n5298), .A2(n17320), .B0(n2793), .Y(n17318)
         );
  AOI21X1 U6394 ( .A0(n5278), .A1(n2820), .B0(n5293), .Y(n17320) );
  INVX1 U6395 ( .A(n17321), .Y(n5293) );
  AND2X2 U6396 ( .A(n2885), .B(n2897), .Y(n465) );
  AND2X2 U6397 ( .A(n3484), .B(n3496), .Y(n466) );
  AND2X2 U6398 ( .A(n2649), .B(n2657), .Y(n467) );
  AND2X2 U6399 ( .A(n3244), .B(n3257), .Y(n468) );
  AND2X2 U6400 ( .A(n3185), .B(n3196), .Y(n469) );
  AND2X2 U6401 ( .A(n2952), .B(n2958), .Y(n470) );
  AND2X2 U6402 ( .A(n2583), .B(n2596), .Y(n471) );
  AND2X2 U6403 ( .A(n3305), .B(n3322), .Y(n472) );
  AND2X2 U6404 ( .A(n3006), .B(n3023), .Y(n473) );
  AND2X2 U6405 ( .A(n2705), .B(n2715), .Y(n474) );
  AND2X2 U6406 ( .A(n3368), .B(n3383), .Y(n475) );
  AND2X2 U6407 ( .A(n3071), .B(n3079), .Y(n476) );
  AND2X2 U6408 ( .A(n2765), .B(n2782), .Y(n477) );
  AND2X2 U6409 ( .A(n3431), .B(n3437), .Y(n478) );
  AND2X2 U6410 ( .A(n3127), .B(n3142), .Y(n479) );
  AND2X2 U6411 ( .A(n2831), .B(n2840), .Y(n480) );
  AND2X2 U6412 ( .A(n2892), .B(n2891), .Y(n481) );
  AND2X2 U6413 ( .A(n3493), .B(n3486), .Y(n482) );
  AND2X2 U6414 ( .A(n2651), .B(n2642), .Y(n483) );
  AND2X2 U6415 ( .A(n3252), .B(n3245), .Y(n484) );
  AND2X2 U6416 ( .A(n2710), .B(n2704), .Y(n485) );
  AND2X2 U6417 ( .A(n3073), .B(n3064), .Y(n486) );
  AND2X2 U6418 ( .A(n3432), .B(n3424), .Y(n487) );
  AND2X2 U6419 ( .A(n2832), .B(n2824), .Y(n488) );
  AND2X2 U6420 ( .A(n3014), .B(n3007), .Y(n489) );
  AND2X2 U6421 ( .A(n3191), .B(n3184), .Y(n490) );
  AND2X2 U6422 ( .A(n3374), .B(n3367), .Y(n491) );
  AND2X2 U6423 ( .A(n2589), .B(n2582), .Y(n492) );
  AND2X2 U6424 ( .A(n2771), .B(n2764), .Y(n493) );
  AND2X2 U6425 ( .A(n2953), .B(n2945), .Y(n494) );
  AND2X2 U6426 ( .A(n3133), .B(n3126), .Y(n495) );
  AND2X2 U6427 ( .A(n3313), .B(n3306), .Y(n496) );
  CLKINVX3 U6428 ( .A(n2652), .Y(n2651) );
  CLKINVX3 U6429 ( .A(n3074), .Y(n3073) );
  CLKINVX3 U6430 ( .A(n3019), .Y(n3016) );
  CLKINVX3 U6431 ( .A(n3379), .Y(n3376) );
  CLKINVX3 U6432 ( .A(n2591), .Y(n2590) );
  CLKINVX3 U6433 ( .A(n2778), .Y(n2773) );
  CLKINVX3 U6434 ( .A(n3138), .Y(n3135) );
  CLKINVX3 U6435 ( .A(n2838), .Y(n2834) );
  INVX1 U6436 ( .A(n10062), .Y(n5345) );
  INVX1 U6437 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n248), .Y(n6141) );
  INVX1 U6438 ( .A(n11230), .Y(n4991) );
  INVX1 U6439 ( .A(n8310), .Y(n5817) );
  INVX1 U6440 ( .A(n10938), .Y(n5075) );
  INVX1 U6441 ( .A(n7434), .Y(n6045) );
  INVX1 U6442 ( .A(n9186), .Y(n5581) );
  INVX1 U6443 ( .A(n10354), .Y(n5261) );
  INVX1 U6444 ( .A(n9478), .Y(n5505) );
  INVX1 U6445 ( .A(n8602), .Y(n5733) );
  INVX1 U6446 ( .A(n7726), .Y(n5969) );
  INVX1 U6447 ( .A(n11522), .Y(n4875) );
  INVX1 U6448 ( .A(n10646), .Y(n5183) );
  INVX1 U6449 ( .A(n9770), .Y(n5429) );
  INVX1 U6450 ( .A(n8894), .Y(n5657) );
  INVX1 U6451 ( .A(n8018), .Y(n5893) );
  AND2X2 U6452 ( .A(n3488), .B(n3496), .Y(n497) );
  AND2X2 U6453 ( .A(n2885), .B(n2901), .Y(n498) );
  AND2X2 U6454 ( .A(n3187), .B(n3200), .Y(n499) );
  AND2X2 U6455 ( .A(n3250), .B(n3261), .Y(n500) );
  AND2X2 U6456 ( .A(n2644), .B(n2664), .Y(n501) );
  AND2X2 U6457 ( .A(n2585), .B(n2603), .Y(n502) );
  AND2X2 U6458 ( .A(n2946), .B(n2962), .Y(n503) );
  AND2X2 U6459 ( .A(n3311), .B(n3327), .Y(n504) );
  AND2X2 U6460 ( .A(n3012), .B(n3019), .Y(n505) );
  AND2X2 U6461 ( .A(n2707), .B(n2719), .Y(n506) );
  AND2X2 U6462 ( .A(n3370), .B(n3379), .Y(n507) );
  AND2X2 U6463 ( .A(n3066), .B(n3086), .Y(n508) );
  AND2X2 U6464 ( .A(n2767), .B(n2785), .Y(n509) );
  AND2X2 U6465 ( .A(n3426), .B(n3441), .Y(n510) );
  AND2X2 U6466 ( .A(n3129), .B(n3138), .Y(n511) );
  AND2X2 U6467 ( .A(n2826), .B(n2845), .Y(n512) );
  AND2X2 U6468 ( .A(n2880), .B(n2894), .Y(n513) );
  AND2X2 U6469 ( .A(n3481), .B(n3497), .Y(n514) );
  AND2X2 U6470 ( .A(n2638), .B(n2662), .Y(n515) );
  AND2X2 U6471 ( .A(n3240), .B(n3254), .Y(n516) );
  AND2X2 U6472 ( .A(n3179), .B(n3193), .Y(n517) );
  AND2X2 U6473 ( .A(n2577), .B(n2601), .Y(n518) );
  AND2X2 U6474 ( .A(n2941), .B(n2955), .Y(n519) );
  AND2X2 U6475 ( .A(n3301), .B(n3318), .Y(n520) );
  AND2X2 U6476 ( .A(n3002), .B(n3018), .Y(n521) );
  AND2X2 U6477 ( .A(n2699), .B(n2722), .Y(n522) );
  AND2X2 U6478 ( .A(n3362), .B(n3378), .Y(n523) );
  AND2X2 U6479 ( .A(n3060), .B(n3084), .Y(n524) );
  AND2X2 U6480 ( .A(n2759), .B(n2777), .Y(n525) );
  AND2X2 U6481 ( .A(n3420), .B(n3444), .Y(n526) );
  AND2X2 U6482 ( .A(n3121), .B(n3137), .Y(n527) );
  AND2X2 U6483 ( .A(n2820), .B(n2838), .Y(n528) );
  AND2X2 U6484 ( .A(n2892), .B(n2891), .Y(n529) );
  AND2X2 U6485 ( .A(n3493), .B(n3486), .Y(n530) );
  AND2X2 U6486 ( .A(n2651), .B(n2648), .Y(n531) );
  AND2X2 U6487 ( .A(n3252), .B(n3243), .Y(n532) );
  AND2X2 U6488 ( .A(n2710), .B(n2706), .Y(n533) );
  AND2X2 U6489 ( .A(n3073), .B(n3070), .Y(n534) );
  AND2X2 U6490 ( .A(n3432), .B(n3430), .Y(n535) );
  AND2X2 U6491 ( .A(n2832), .B(n2830), .Y(n536) );
  AND2X2 U6492 ( .A(n3014), .B(n3005), .Y(n537) );
  AND2X2 U6493 ( .A(n3191), .B(n3186), .Y(n538) );
  AND2X2 U6494 ( .A(n3374), .B(n3369), .Y(n539) );
  AND2X2 U6495 ( .A(n2589), .B(n2584), .Y(n540) );
  AND2X2 U6496 ( .A(n2771), .B(n2766), .Y(n541) );
  AND2X2 U6497 ( .A(n2953), .B(n2951), .Y(n542) );
  AND2X2 U6498 ( .A(n3133), .B(n3128), .Y(n543) );
  AND2X2 U6499 ( .A(n3313), .B(n3304), .Y(n544) );
  INVXL U6500 ( .A(n9988), .Y(n5351) );
  INVXL U6501 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n174), .Y(n6147) );
  INVXL U6502 ( .A(n11156), .Y(n4997) );
  INVXL U6503 ( .A(n8236), .Y(n5823) );
  INVXL U6504 ( .A(n10864), .Y(n5081) );
  INVXL U6505 ( .A(n9112), .Y(n5587) );
  INVXL U6506 ( .A(n7360), .Y(n6051) );
  INVXL U6507 ( .A(n10280), .Y(n5267) );
  INVXL U6508 ( .A(n9404), .Y(n5511) );
  INVXL U6509 ( .A(n8528), .Y(n5739) );
  INVXL U6510 ( .A(n7652), .Y(n5975) );
  INVXL U6511 ( .A(n11448), .Y(n4881) );
  INVXL U6512 ( .A(n10572), .Y(n5189) );
  INVXL U6513 ( .A(n9696), .Y(n5435) );
  INVXL U6514 ( .A(n8820), .Y(n5663) );
  INVXL U6515 ( .A(n7944), .Y(n5899) );
  INVX1 U6516 ( .A(top_core_EC_n1021), .Y(n6307) );
  INVX1 U6517 ( .A(n2510), .Y(n2438) );
  INVX1 U6518 ( .A(n2511), .Y(n2435) );
  INVX1 U6519 ( .A(n2513), .Y(n2429) );
  INVX1 U6520 ( .A(n2512), .Y(n2434) );
  INVX1 U6521 ( .A(n2511), .Y(n2436) );
  INVX1 U6522 ( .A(n2513), .Y(n2430) );
  INVX1 U6523 ( .A(n2510), .Y(n2440) );
  INVX1 U6524 ( .A(n2510), .Y(n2439) );
  INVX1 U6525 ( .A(n2513), .Y(n2431) );
  INVX1 U6526 ( .A(n2512), .Y(n2432) );
  INVX1 U6527 ( .A(n2512), .Y(n2433) );
  INVX1 U6528 ( .A(n2511), .Y(n2437) );
  INVX1 U6529 ( .A(n2504), .Y(n2463) );
  INVX1 U6530 ( .A(n2367), .Y(n2441) );
  INVX1 U6531 ( .A(n2509), .Y(n2446) );
  INVX1 U6532 ( .A(n2507), .Y(n2454) );
  INVX1 U6533 ( .A(n2394), .Y(n2443) );
  INVX1 U6534 ( .A(n2369), .Y(n2445) );
  INVX1 U6535 ( .A(n2503), .Y(n2464) );
  INVX1 U6536 ( .A(n2501), .Y(n2472) );
  INVX1 U6537 ( .A(n2504), .Y(n2462) );
  INVX1 U6538 ( .A(n2509), .Y(n2447) );
  INVX1 U6539 ( .A(n2393), .Y(n2442) );
  INVX1 U6540 ( .A(n2509), .Y(n2448) );
  INVX1 U6541 ( .A(n2503), .Y(n2465) );
  INVX1 U6542 ( .A(n2372), .Y(n2444) );
  INVX1 U6543 ( .A(n2508), .Y(n2449) );
  INVX1 U6544 ( .A(n2508), .Y(n2450) );
  INVX1 U6545 ( .A(n2508), .Y(n2451) );
  INVX1 U6546 ( .A(n2507), .Y(n2452) );
  INVX1 U6547 ( .A(n2507), .Y(n2453) );
  INVX1 U6548 ( .A(n2506), .Y(n2455) );
  INVX1 U6549 ( .A(n2506), .Y(n2456) );
  INVX1 U6550 ( .A(n2506), .Y(n2457) );
  INVX1 U6551 ( .A(n2505), .Y(n2458) );
  INVX1 U6552 ( .A(n2505), .Y(n2459) );
  INVX1 U6553 ( .A(n2505), .Y(n2460) );
  INVX1 U6554 ( .A(n2504), .Y(n2461) );
  INVX1 U6555 ( .A(n2500), .Y(n2475) );
  INVX1 U6556 ( .A(n2500), .Y(n2474) );
  INVX1 U6557 ( .A(n2500), .Y(n2473) );
  INVX1 U6558 ( .A(n2501), .Y(n2471) );
  INVX1 U6559 ( .A(n2501), .Y(n2470) );
  INVX1 U6560 ( .A(n2502), .Y(n2469) );
  INVX1 U6561 ( .A(n2502), .Y(n2468) );
  INVX1 U6562 ( .A(n2502), .Y(n2467) );
  INVX1 U6563 ( .A(n2503), .Y(n2466) );
  INVX1 U6564 ( .A(n2499), .Y(n2476) );
  INVX1 U6565 ( .A(n2499), .Y(n2477) );
  INVX1 U6566 ( .A(n2499), .Y(n2478) );
  INVX1 U6567 ( .A(n2498), .Y(n2479) );
  INVX1 U6568 ( .A(n2498), .Y(n2480) );
  INVX1 U6569 ( .A(n2498), .Y(n2481) );
  INVX1 U6570 ( .A(n2497), .Y(n2482) );
  INVX1 U6571 ( .A(n2497), .Y(n2483) );
  INVX1 U6572 ( .A(n2497), .Y(n2484) );
  INVX1 U6573 ( .A(n3625), .Y(n3619) );
  INVX1 U6574 ( .A(n3624), .Y(n3620) );
  INVX1 U6575 ( .A(n3624), .Y(n3614) );
  INVX1 U6576 ( .A(n3627), .Y(n3615) );
  INVX1 U6577 ( .A(n3624), .Y(n3621) );
  INVX1 U6578 ( .A(n3625), .Y(n3618) );
  INVX1 U6579 ( .A(n3591), .Y(n3617) );
  INVX1 U6580 ( .A(n3601), .Y(n3622) );
  INVX1 U6581 ( .A(n3600), .Y(n3623) );
  INVX1 U6582 ( .A(n3625), .Y(n3616) );
  INVX1 U6583 ( .A(top_core_KE_n2182), .Y(n2345) );
  INVX1 U6584 ( .A(top_core_KE_n2182), .Y(n2346) );
  NOR2X2 U6585 ( .A(n3452), .B(n3447), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n93) );
  NOR2X2 U6586 ( .A(n2851), .B(n2846), .Y(n9909) );
  NOR2X2 U6587 ( .A(n2609), .B(n2604), .Y(n11077) );
  NOR2X2 U6588 ( .A(n3211), .B(n3206), .Y(n8157) );
  NOR2X2 U6589 ( .A(n2670), .B(n2665), .Y(n10785) );
  NOR2X2 U6590 ( .A(n3031), .B(n3026), .Y(n9033) );
  NOR2X2 U6591 ( .A(n3391), .B(n3386), .Y(n7281) );
  NOR2X2 U6592 ( .A(n2791), .B(n2786), .Y(n10201) );
  NOR2X2 U6593 ( .A(n2973), .B(n2968), .Y(n9325) );
  NOR2X2 U6594 ( .A(n3150), .B(n3145), .Y(n8449) );
  NOR2X2 U6595 ( .A(n3333), .B(n3328), .Y(n7573) );
  NOR2X2 U6596 ( .A(n2548), .B(n2543), .Y(n11369) );
  NOR2X2 U6597 ( .A(n2730), .B(n2725), .Y(n10493) );
  NOR2X2 U6598 ( .A(n2912), .B(n2907), .Y(n9617) );
  NOR2X2 U6599 ( .A(n3092), .B(n3087), .Y(n8741) );
  NOR2X2 U6600 ( .A(n3272), .B(n3267), .Y(n7865) );
  NAND2X2 U6601 ( .A(n5363), .B(n2877), .Y(n17073) );
  NAND2X2 U6602 ( .A(n6131), .B(n3477), .Y(n13923) );
  NAND2X2 U6603 ( .A(n5009), .B(n2635), .Y(n18333) );
  NAND2X2 U6604 ( .A(n5835), .B(n3237), .Y(n15183) );
  NAND2X2 U6605 ( .A(n5751), .B(n3176), .Y(n15498) );
  NAND2X2 U6606 ( .A(n5447), .B(n2937), .Y(n16758) );
  NAND2X2 U6607 ( .A(n4893), .B(n2574), .Y(n18648) );
  NAND2X2 U6608 ( .A(n5911), .B(n3297), .Y(n14868) );
  NAND2X2 U6609 ( .A(n5523), .B(n2998), .Y(n16443) );
  NAND2X2 U6610 ( .A(n5093), .B(n2695), .Y(n18018) );
  NAND2X2 U6611 ( .A(n5987), .B(n3359), .Y(n14553) );
  NAND2X2 U6612 ( .A(n5599), .B(n3057), .Y(n16128) );
  NAND2X2 U6613 ( .A(n5201), .B(n2756), .Y(n17703) );
  NAND2X2 U6614 ( .A(n6063), .B(n3416), .Y(n14238) );
  NAND2X2 U6615 ( .A(n5675), .B(n3118), .Y(n15813) );
  NAND2X2 U6616 ( .A(n5279), .B(n2816), .Y(n17388) );
  NOR3X1 U6617 ( .A(n3989), .B(n2512), .C(n4058), .Y(top_core_EC_n1022) );
  NOR2X2 U6618 ( .A(n2851), .B(n2846), .Y(n17051) );
  NOR2X2 U6619 ( .A(n3452), .B(n3447), .Y(n13901) );
  NOR2X2 U6620 ( .A(n2609), .B(n2604), .Y(n18311) );
  NOR2X2 U6621 ( .A(n3211), .B(n3206), .Y(n15161) );
  NOR2X2 U6622 ( .A(n3150), .B(n3145), .Y(n15476) );
  NOR2X2 U6623 ( .A(n2548), .B(n2543), .Y(n18626) );
  NOR2X2 U6624 ( .A(n2912), .B(n2907), .Y(n16736) );
  NOR2X2 U6625 ( .A(n3272), .B(n3267), .Y(n14846) );
  NOR2X2 U6626 ( .A(n2973), .B(n2968), .Y(n16421) );
  NOR2X2 U6627 ( .A(n2670), .B(n2665), .Y(n17996) );
  NOR2X2 U6628 ( .A(n3333), .B(n3328), .Y(n14531) );
  NOR2X2 U6629 ( .A(n3031), .B(n3026), .Y(n16106) );
  NOR2X2 U6630 ( .A(n2730), .B(n2725), .Y(n17681) );
  NOR2X2 U6631 ( .A(n3391), .B(n3386), .Y(n14216) );
  NOR2X2 U6632 ( .A(n3092), .B(n3087), .Y(n15791) );
  NOR2X2 U6633 ( .A(n2791), .B(n2786), .Y(n17366) );
  AOI22X1 U6634 ( .A0(n2871), .A1(n2898), .B0(n2873), .B1(n481), .Y(n17074) );
  AOI22X1 U6635 ( .A0(n3472), .A1(n3495), .B0(n3475), .B1(n482), .Y(n13924) );
  AOI22X1 U6636 ( .A0(n2629), .A1(n2655), .B0(n2631), .B1(n483), .Y(n18334) );
  AOI22X1 U6637 ( .A0(n3231), .A1(n3258), .B0(n3234), .B1(n484), .Y(n15184) );
  AOI22X1 U6638 ( .A0(n3170), .A1(n3197), .B0(n3173), .B1(n490), .Y(n15499) );
  AOI22X1 U6639 ( .A0(n2568), .A1(n2594), .B0(n2570), .B1(n492), .Y(n18649) );
  AOI22X1 U6640 ( .A0(n2932), .A1(n2959), .B0(n2934), .B1(n494), .Y(n16759) );
  AOI22X1 U6641 ( .A0(n3292), .A1(n3316), .B0(n3294), .B1(n496), .Y(n14869) );
  AOI22X1 U6642 ( .A0(n2993), .A1(n3017), .B0(n2995), .B1(n489), .Y(n16444) );
  AOI22X1 U6643 ( .A0(n2690), .A1(n2712), .B0(n2692), .B1(n485), .Y(n18019) );
  AOI22X1 U6644 ( .A0(n3353), .A1(n3377), .B0(n3356), .B1(n491), .Y(n14554) );
  AOI22X1 U6645 ( .A0(n3051), .A1(n3077), .B0(n3053), .B1(n486), .Y(n16129) );
  AOI22X1 U6646 ( .A0(n2750), .A1(n2775), .B0(n2753), .B1(n493), .Y(n17704) );
  AOI22X1 U6647 ( .A0(n3411), .A1(n3434), .B0(n3413), .B1(n487), .Y(n14239) );
  AOI22X1 U6648 ( .A0(n3112), .A1(n3136), .B0(n3114), .B1(n495), .Y(n15814) );
  AOI22X1 U6649 ( .A0(n2811), .A1(n2836), .B0(n2813), .B1(n488), .Y(n17389) );
  NOR2X1 U6650 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n128), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n86) );
  NOR2X1 U6651 ( .A(n9970), .B(n9943), .Y(n9903) );
  NOR2X1 U6652 ( .A(n11138), .B(n11111), .Y(n11071) );
  NOR2X1 U6653 ( .A(n8218), .B(n8191), .Y(n8151) );
  NOR2X1 U6654 ( .A(n10846), .B(n10819), .Y(n10779) );
  NOR2X1 U6655 ( .A(n9094), .B(n9067), .Y(n9027) );
  NOR2X1 U6656 ( .A(n7342), .B(n7315), .Y(n7275) );
  NOR2X1 U6657 ( .A(n10262), .B(n10235), .Y(n10195) );
  NOR2X1 U6658 ( .A(n9386), .B(n9359), .Y(n9319) );
  NOR2X1 U6659 ( .A(n8510), .B(n8483), .Y(n8443) );
  NOR2X1 U6660 ( .A(n7634), .B(n7607), .Y(n7567) );
  NOR2X1 U6661 ( .A(n11430), .B(n11403), .Y(n11363) );
  NOR2X1 U6662 ( .A(n10554), .B(n10527), .Y(n10487) );
  NOR2X1 U6663 ( .A(n9678), .B(n9651), .Y(n9611) );
  NOR2X1 U6664 ( .A(n8802), .B(n8775), .Y(n8735) );
  NOR2X1 U6665 ( .A(n7926), .B(n7899), .Y(n7859) );
  NOR2X1 U6666 ( .A(n9943), .B(n513), .Y(n9926) );
  NOR2X1 U6667 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n128), .B(n514), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n111) );
  NOR2X1 U6668 ( .A(n11111), .B(n515), .Y(n11094) );
  NOR2X1 U6669 ( .A(n8191), .B(n516), .Y(n8174) );
  NOR2X1 U6670 ( .A(n10819), .B(n522), .Y(n10802) );
  NOR2X1 U6671 ( .A(n7315), .B(n526), .Y(n7298) );
  NOR2X1 U6672 ( .A(n9067), .B(n524), .Y(n9050) );
  NOR2X1 U6673 ( .A(n10235), .B(n528), .Y(n10218) );
  NOR2X1 U6674 ( .A(n9359), .B(n521), .Y(n9342) );
  NOR2X1 U6675 ( .A(n8483), .B(n517), .Y(n8466) );
  NOR2X1 U6676 ( .A(n7607), .B(n523), .Y(n7590) );
  NOR2X1 U6677 ( .A(n11403), .B(n518), .Y(n11386) );
  NOR2X1 U6678 ( .A(n10527), .B(n525), .Y(n10510) );
  NOR2X1 U6679 ( .A(n9651), .B(n519), .Y(n9634) );
  NOR2X1 U6680 ( .A(n8775), .B(n527), .Y(n8758) );
  NOR2X1 U6681 ( .A(n7899), .B(n520), .Y(n7882) );
  NAND2X1 U6682 ( .A(n686), .B(n1151), .Y(n13384) );
  NAND2X1 U6683 ( .A(n688), .B(n1191), .Y(n12754) );
  NAND2X1 U6684 ( .A(n687), .B(n1200), .Y(n13069) );
  NOR2X1 U6685 ( .A(n17208), .B(n17061), .Y(n17098) );
  NOR2X1 U6686 ( .A(n14058), .B(n13911), .Y(n13948) );
  NOR2X1 U6687 ( .A(n18468), .B(n18321), .Y(n18358) );
  NOR2X1 U6688 ( .A(n15318), .B(n15171), .Y(n15208) );
  NOR2X1 U6689 ( .A(n15633), .B(n15486), .Y(n15523) );
  NOR2X1 U6690 ( .A(n18783), .B(n18636), .Y(n18673) );
  NOR2X1 U6691 ( .A(n16893), .B(n16746), .Y(n16783) );
  NOR2X1 U6692 ( .A(n15003), .B(n14856), .Y(n14893) );
  NOR2X1 U6693 ( .A(n16578), .B(n16431), .Y(n16468) );
  NOR2X1 U6694 ( .A(n18153), .B(n18006), .Y(n18043) );
  NOR2X1 U6695 ( .A(n14688), .B(n14541), .Y(n14578) );
  NOR2X1 U6696 ( .A(n16263), .B(n16116), .Y(n16153) );
  NOR2X1 U6697 ( .A(n17838), .B(n17691), .Y(n17728) );
  NOR2X1 U6698 ( .A(n14373), .B(n14226), .Y(n14263) );
  NOR2X1 U6699 ( .A(n15948), .B(n15801), .Y(n15838) );
  NOR2X1 U6700 ( .A(n17523), .B(n17376), .Y(n17413) );
  NOR2X1 U6701 ( .A(n17061), .B(n164), .Y(n17037) );
  NOR2X1 U6702 ( .A(n13911), .B(n165), .Y(n13887) );
  NOR2X1 U6703 ( .A(n18321), .B(n166), .Y(n18297) );
  NOR2X1 U6704 ( .A(n15171), .B(n167), .Y(n15147) );
  NOR2X1 U6705 ( .A(n15486), .B(n168), .Y(n15462) );
  NOR2X1 U6706 ( .A(n18636), .B(n169), .Y(n18612) );
  NOR2X1 U6707 ( .A(n16746), .B(n170), .Y(n16722) );
  NOR2X1 U6708 ( .A(n14856), .B(n171), .Y(n14832) );
  NOR2X1 U6709 ( .A(n16431), .B(n172), .Y(n16407) );
  NOR2X1 U6710 ( .A(n18006), .B(n173), .Y(n17982) );
  NOR2X1 U6711 ( .A(n14541), .B(n174), .Y(n14517) );
  NOR2X1 U6712 ( .A(n16116), .B(n175), .Y(n16092) );
  NOR2X1 U6713 ( .A(n17691), .B(n176), .Y(n17667) );
  NOR2X1 U6714 ( .A(n14226), .B(n177), .Y(n14202) );
  NOR2X1 U6715 ( .A(n15801), .B(n178), .Y(n15777) );
  NOR2X1 U6716 ( .A(n17376), .B(n179), .Y(n17352) );
  NOR2X1 U6717 ( .A(n9944), .B(n2883), .Y(n10064) );
  NOR2X1 U6718 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n129), .B(n3485), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n250) );
  NOR2X1 U6719 ( .A(n11112), .B(n2641), .Y(n11232) );
  NOR2X1 U6720 ( .A(n8192), .B(n3251), .Y(n8312) );
  NOR2X1 U6721 ( .A(n10820), .B(n2707), .Y(n10940) );
  NOR2X1 U6722 ( .A(n7316), .B(n3423), .Y(n7436) );
  NOR2X1 U6723 ( .A(n9068), .B(n3063), .Y(n9188) );
  NOR2X1 U6724 ( .A(n10236), .B(n2823), .Y(n10356) );
  NOR2X1 U6725 ( .A(n9360), .B(n3013), .Y(n9480) );
  NOR2X1 U6726 ( .A(n8484), .B(n3187), .Y(n8604) );
  NOR2X1 U6727 ( .A(n7608), .B(n3370), .Y(n7728) );
  NOR2X1 U6728 ( .A(n11404), .B(n2585), .Y(n11524) );
  NOR2X1 U6729 ( .A(n10528), .B(n2767), .Y(n10648) );
  NOR2X1 U6730 ( .A(n9652), .B(n2944), .Y(n9772) );
  NOR2X1 U6731 ( .A(n8776), .B(n3129), .Y(n8896) );
  NOR2X1 U6732 ( .A(n7900), .B(n3312), .Y(n8020) );
  NOR2X1 U6733 ( .A(n9900), .B(n9944), .Y(n10004) );
  NOR2X1 U6734 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n129), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n190) );
  NOR2X1 U6735 ( .A(n11068), .B(n11112), .Y(n11172) );
  NOR2X1 U6736 ( .A(n8148), .B(n8192), .Y(n8252) );
  NOR2X1 U6737 ( .A(n10776), .B(n10820), .Y(n10880) );
  NOR2X1 U6738 ( .A(n9024), .B(n9068), .Y(n9128) );
  NOR2X1 U6739 ( .A(n7272), .B(n7316), .Y(n7376) );
  NOR2X1 U6740 ( .A(n10192), .B(n10236), .Y(n10296) );
  NOR2X1 U6741 ( .A(n9316), .B(n9360), .Y(n9420) );
  NOR2X1 U6742 ( .A(n8440), .B(n8484), .Y(n8544) );
  NOR2X1 U6743 ( .A(n7564), .B(n7608), .Y(n7668) );
  NOR2X1 U6744 ( .A(n11360), .B(n11404), .Y(n11464) );
  NOR2X1 U6745 ( .A(n10484), .B(n10528), .Y(n10588) );
  NOR2X1 U6746 ( .A(n9608), .B(n9652), .Y(n9712) );
  NOR2X1 U6747 ( .A(n8732), .B(n8776), .Y(n8836) );
  NOR2X1 U6748 ( .A(n7856), .B(n7900), .Y(n7960) );
  AOI22X1 U6749 ( .A0(n2880), .A1(n2876), .B0(n2871), .B1(n529), .Y(n17093) );
  AOI22X1 U6750 ( .A0(n2638), .A1(n2634), .B0(n2629), .B1(n531), .Y(n18353) );
  AOI22X1 U6751 ( .A0(n3240), .A1(n3235), .B0(n3231), .B1(n532), .Y(n15203) );
  AOI22X1 U6752 ( .A0(n3179), .A1(n3174), .B0(n3170), .B1(n538), .Y(n15518) );
  AOI22X1 U6753 ( .A0(n2941), .A1(n2937), .B0(n2932), .B1(n542), .Y(n16778) );
  AOI22X1 U6754 ( .A0(n2577), .A1(n2573), .B0(n2568), .B1(n540), .Y(n18668) );
  AOI22X1 U6755 ( .A0(n3301), .A1(n3296), .B0(n3292), .B1(n544), .Y(n14888) );
  AOI22X1 U6756 ( .A0(n3002), .A1(n2998), .B0(n2993), .B1(n537), .Y(n16463) );
  AOI22X1 U6757 ( .A0(n2699), .A1(n2695), .B0(n2690), .B1(n533), .Y(n18038) );
  AOI22X1 U6758 ( .A0(n3362), .A1(n3357), .B0(n3353), .B1(n539), .Y(n14573) );
  AOI22X1 U6759 ( .A0(n3060), .A1(n3056), .B0(n3051), .B1(n534), .Y(n16148) );
  AOI22X1 U6760 ( .A0(n2759), .A1(n2754), .B0(n2750), .B1(n541), .Y(n17723) );
  AOI22X1 U6761 ( .A0(n3420), .A1(n3416), .B0(n3411), .B1(n535), .Y(n14258) );
  AOI22X1 U6762 ( .A0(n3121), .A1(n3117), .B0(n3112), .B1(n543), .Y(n15833) );
  AOI22X1 U6763 ( .A0(n2820), .A1(n2815), .B0(n2811), .B1(n536), .Y(n17408) );
  NOR2X1 U6764 ( .A(n14058), .B(n3485), .Y(n13849) );
  NOR2X1 U6765 ( .A(n17208), .B(n2886), .Y(n16999) );
  NOR2X1 U6766 ( .A(n18468), .B(n2648), .Y(n18259) );
  NOR2X1 U6767 ( .A(n15318), .B(n3244), .Y(n15109) );
  NOR2X1 U6768 ( .A(n15633), .B(n3182), .Y(n15424) );
  NOR2X1 U6769 ( .A(n18783), .B(n2580), .Y(n18574) );
  NOR2X1 U6770 ( .A(n16893), .B(n2945), .Y(n16684) );
  NOR2X1 U6771 ( .A(n15003), .B(n3305), .Y(n14794) );
  NOR2X1 U6772 ( .A(n16578), .B(n3006), .Y(n16369) );
  NOR2X1 U6773 ( .A(n18153), .B(n2702), .Y(n17944) );
  NOR2X1 U6774 ( .A(n14688), .B(n3365), .Y(n14479) );
  NOR2X1 U6775 ( .A(n16263), .B(n3064), .Y(n16054) );
  NOR2X1 U6776 ( .A(n17838), .B(n2762), .Y(n17629) );
  NOR2X1 U6777 ( .A(n14373), .B(n3430), .Y(n14164) );
  NOR2X1 U6778 ( .A(n15948), .B(n3124), .Y(n15739) );
  NOR2X1 U6779 ( .A(n17523), .B(n2824), .Y(n17314) );
  NOR2X1 U6780 ( .A(n1152), .B(n6544), .Y(n13443) );
  NOR2X1 U6781 ( .A(n1192), .B(n6839), .Y(n12813) );
  NOR2X1 U6782 ( .A(n1201), .B(n6885), .Y(n13128) );
  NAND2X1 U6783 ( .A(n6919), .B(n613), .Y(n11787) );
  NAND2X1 U6784 ( .A(n6873), .B(n614), .Y(top_core_KE_sb1_n215) );
  NAND2X1 U6785 ( .A(n6579), .B(n615), .Y(n12103) );
  NAND2X1 U6786 ( .A(n6554), .B(n1174), .Y(n13363) );
  NAND2X1 U6787 ( .A(n6849), .B(n1214), .Y(n12733) );
  NAND2X1 U6788 ( .A(n6602), .B(n1179), .Y(n13678) );
  NAND2X1 U6789 ( .A(n6895), .B(n1220), .Y(n13048) );
  NAND2X1 U6790 ( .A(n2846), .B(n2857), .Y(n9990) );
  NAND2X1 U6791 ( .A(n3447), .B(n3458), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n176) );
  NAND2X1 U6792 ( .A(n2604), .B(n2615), .Y(n11158) );
  NAND2X1 U6793 ( .A(n3206), .B(n3217), .Y(n8238) );
  NAND2X1 U6794 ( .A(n2665), .B(n2676), .Y(n10866) );
  NAND2X1 U6795 ( .A(n3026), .B(n3037), .Y(n9114) );
  NAND2X1 U6796 ( .A(n3386), .B(n3397), .Y(n7362) );
  NAND2X1 U6797 ( .A(n2786), .B(n2797), .Y(n10282) );
  NAND2X1 U6798 ( .A(n2968), .B(n2979), .Y(n9406) );
  NAND2X1 U6799 ( .A(n3145), .B(n3156), .Y(n8530) );
  NAND2X1 U6800 ( .A(n3328), .B(n3339), .Y(n7654) );
  NAND2X1 U6801 ( .A(n2543), .B(n2554), .Y(n11450) );
  NAND2X1 U6802 ( .A(n2725), .B(n2736), .Y(n10574) );
  NAND2X1 U6803 ( .A(n2907), .B(n2918), .Y(n9698) );
  NAND2X1 U6804 ( .A(n3087), .B(n3098), .Y(n8822) );
  NAND2X1 U6805 ( .A(n3267), .B(n3278), .Y(n7946) );
  AND2X2 U6806 ( .A(n2171), .B(n2290), .Y(top_core_KE_n2182) );
  NAND2X1 U6807 ( .A(n1152), .B(n1173), .Y(n13334) );
  NAND2X1 U6808 ( .A(n1192), .B(n1213), .Y(n12704) );
  NAND2X1 U6809 ( .A(n1201), .B(n1219), .Y(n13019) );
  NAND2X1 U6810 ( .A(n3478), .B(n3469), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n98) );
  NAND2X1 U6811 ( .A(n2874), .B(n2870), .Y(n9914) );
  NAND2X1 U6812 ( .A(n2632), .B(n2628), .Y(n11082) );
  NAND2X1 U6813 ( .A(n3238), .B(n3230), .Y(n8162) );
  NAND2X1 U6814 ( .A(n2696), .B(n2688), .Y(n10790) );
  NAND2X1 U6815 ( .A(n3054), .B(n3050), .Y(n9038) );
  NAND2X1 U6816 ( .A(n3417), .B(n3410), .Y(n7286) );
  NAND2X1 U6817 ( .A(n2817), .B(n2810), .Y(n10206) );
  NAND2X1 U6818 ( .A(n2999), .B(n2992), .Y(n9330) );
  NAND2X1 U6819 ( .A(n3177), .B(n3169), .Y(n8454) );
  NAND2X1 U6820 ( .A(n3360), .B(n3352), .Y(n7578) );
  NAND2X1 U6821 ( .A(n2571), .B(n2567), .Y(n11374) );
  NAND2X1 U6822 ( .A(n2757), .B(n2748), .Y(n10498) );
  NAND2X1 U6823 ( .A(n2938), .B(n2931), .Y(n9622) );
  NAND2X1 U6824 ( .A(n3115), .B(n3111), .Y(n8746) );
  NAND2X1 U6825 ( .A(n3298), .B(n3291), .Y(n7870) );
  NOR2XL U6826 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n70), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n186) );
  NOR2XL U6827 ( .A(n8139), .B(n8136), .Y(n8248) );
  NAND2X1 U6828 ( .A(n6131), .B(n3473), .Y(n13864) );
  NAND2X1 U6829 ( .A(n5363), .B(n2872), .Y(n17014) );
  NAND2X1 U6830 ( .A(n5009), .B(n2630), .Y(n18274) );
  NAND2X1 U6831 ( .A(n5835), .B(n3232), .Y(n15124) );
  NAND2X1 U6832 ( .A(n5751), .B(n3171), .Y(n15439) );
  NAND2X1 U6833 ( .A(n4893), .B(n2569), .Y(n18589) );
  NAND2X1 U6834 ( .A(n5447), .B(n2933), .Y(n16699) );
  NAND2X1 U6835 ( .A(n5911), .B(n3293), .Y(n14809) );
  NAND2X1 U6836 ( .A(n5523), .B(n2994), .Y(n16384) );
  NAND2X1 U6837 ( .A(n5093), .B(n2691), .Y(n17959) );
  NAND2X1 U6838 ( .A(n5987), .B(n3354), .Y(n14494) );
  NAND2X1 U6839 ( .A(n5599), .B(n3052), .Y(n16069) );
  NAND2X1 U6840 ( .A(n5201), .B(n2751), .Y(n17644) );
  NAND2X1 U6841 ( .A(n6063), .B(n3412), .Y(n14179) );
  NAND2X1 U6842 ( .A(n5675), .B(n3113), .Y(n15754) );
  NAND2X1 U6843 ( .A(n5279), .B(n2812), .Y(n17329) );
  OAI22X1 U6844 ( .A0(top_core_EC_mc_n2), .A1(n2413), .B0(n2367), .B1(
        top_core_EC_mc_n3), .Y(top_core_EC_mix_out_9_) );
  XOR2X1 U6845 ( .A(top_core_EC_mc_n4), .B(top_core_EC_mc_n5), .Y(
        top_core_EC_mc_n3) );
  XNOR2X1 U6846 ( .A(top_core_EC_mc_mix_in_4_10_), .B(top_core_EC_mc_n6), .Y(
        top_core_EC_mc_n2) );
  XNOR2X1 U6847 ( .A(top_core_EC_mc_mix_in_4_10_), .B(top_core_EC_mc_n8), .Y(
        top_core_EC_mc_n4) );
  OAI22X1 U6848 ( .A0(top_core_EC_mc_n772), .A1(n2416), .B0(n2377), .B1(
        top_core_EC_mc_n773), .Y(top_core_EC_mix_out_11_) );
  XOR2X1 U6849 ( .A(top_core_EC_mc_n774), .B(top_core_EC_mc_n775), .Y(
        top_core_EC_mc_n773) );
  XNOR2X1 U6850 ( .A(top_core_EC_mc_mix_in_2_11_), .B(top_core_EC_mc_n776), 
        .Y(top_core_EC_mc_n772) );
  XNOR2X1 U6851 ( .A(top_core_EC_mc_mix_in_2_11_), .B(top_core_EC_mc_n498), 
        .Y(top_core_EC_mc_n774) );
  OAI22X1 U6852 ( .A0(top_core_EC_mc_n705), .A1(n2466), .B0(n2377), .B1(
        top_core_EC_mc_n706), .Y(top_core_EC_mix_out_12_) );
  XOR2X1 U6853 ( .A(top_core_EC_mc_n707), .B(top_core_EC_mc_n708), .Y(
        top_core_EC_mc_n706) );
  XNOR2X1 U6854 ( .A(top_core_EC_mc_mix_in_8[14]), .B(top_core_EC_mc_n709), 
        .Y(top_core_EC_mc_n705) );
  XNOR2X1 U6855 ( .A(top_core_EC_mc_mix_in_8[14]), .B(top_core_EC_mc_n433), 
        .Y(top_core_EC_mc_n707) );
  OAI22X1 U6856 ( .A0(top_core_EC_mc_n671), .A1(n2472), .B0(n2378), .B1(
        top_core_EC_mc_n672), .Y(top_core_EC_mix_out_17_) );
  XOR2X1 U6857 ( .A(top_core_EC_mc_n618), .B(top_core_EC_mc_n673), .Y(
        top_core_EC_mc_n672) );
  XNOR2X1 U6858 ( .A(top_core_EC_mc_mix_in_4_26_), .B(top_core_EC_mc_n674), 
        .Y(top_core_EC_mc_n671) );
  XOR2X1 U6859 ( .A(top_core_EC_mc_n657), .B(top_core_EC_mc_n674), .Y(
        top_core_EC_mc_n673) );
  OAI22X1 U6860 ( .A0(top_core_EC_mc_n659), .A1(n2471), .B0(n2378), .B1(
        top_core_EC_mc_n660), .Y(top_core_EC_mix_out_19_) );
  XOR2X1 U6861 ( .A(top_core_EC_mc_n604), .B(top_core_EC_mc_n661), .Y(
        top_core_EC_mc_n660) );
  XNOR2X1 U6862 ( .A(top_core_EC_mc_mix_in_2_27_), .B(top_core_EC_mc_n662), 
        .Y(top_core_EC_mc_n659) );
  XOR2X1 U6863 ( .A(top_core_EC_mc_n497), .B(top_core_EC_mc_n662), .Y(
        top_core_EC_mc_n661) );
  OAI22X1 U6864 ( .A0(top_core_EC_mc_n646), .A1(n2417), .B0(n2378), .B1(
        top_core_EC_mc_n647), .Y(top_core_EC_mix_out_20_) );
  XOR2X1 U6865 ( .A(top_core_EC_mc_n597), .B(top_core_EC_mc_n648), .Y(
        top_core_EC_mc_n647) );
  XNOR2X1 U6866 ( .A(top_core_EC_mc_mix_in_8[30]), .B(top_core_EC_mc_n649), 
        .Y(top_core_EC_mc_n646) );
  XOR2X1 U6867 ( .A(top_core_EC_mc_n432), .B(top_core_EC_mc_n649), .Y(
        top_core_EC_mc_n648) );
  OAI22X1 U6868 ( .A0(top_core_EC_mc_n616), .A1(n2477), .B0(n2378), .B1(
        top_core_EC_mc_n617), .Y(top_core_EC_mix_out_25_) );
  XOR2X1 U6869 ( .A(top_core_EC_mc_n618), .B(top_core_EC_mc_n619), .Y(
        top_core_EC_mc_n617) );
  XNOR2X1 U6870 ( .A(top_core_EC_mc_mix_in_4_26_), .B(top_core_EC_mc_n620), 
        .Y(top_core_EC_mc_n616) );
  XOR2X1 U6871 ( .A(top_core_EC_mc_n7), .B(top_core_EC_mc_n620), .Y(
        top_core_EC_mc_n619) );
  OAI22X1 U6872 ( .A0(top_core_EC_mc_n602), .A1(n2478), .B0(n2379), .B1(
        top_core_EC_mc_n603), .Y(top_core_EC_mix_out_27_) );
  XOR2X1 U6873 ( .A(top_core_EC_mc_n604), .B(top_core_EC_mc_n605), .Y(
        top_core_EC_mc_n603) );
  XNOR2X1 U6874 ( .A(top_core_EC_mc_mix_in_2_27_), .B(top_core_EC_mc_n606), 
        .Y(top_core_EC_mc_n602) );
  XOR2X1 U6875 ( .A(top_core_EC_mc_n606), .B(top_core_EC_mc_n607), .Y(
        top_core_EC_mc_n605) );
  OAI22X1 U6876 ( .A0(top_core_EC_mc_n595), .A1(n2478), .B0(n2379), .B1(
        top_core_EC_mc_n596), .Y(top_core_EC_mix_out_28_) );
  XOR2X1 U6877 ( .A(top_core_EC_mc_n597), .B(top_core_EC_mc_n598), .Y(
        top_core_EC_mc_n596) );
  XNOR2X1 U6878 ( .A(top_core_EC_mc_mix_in_8[30]), .B(top_core_EC_mc_n599), 
        .Y(top_core_EC_mc_n595) );
  XOR2X1 U6879 ( .A(top_core_EC_mc_n599), .B(top_core_EC_mc_n600), .Y(
        top_core_EC_mc_n598) );
  OAI22X1 U6880 ( .A0(top_core_EC_mc_n482), .A1(n2483), .B0(n2380), .B1(
        top_core_EC_mc_n483), .Y(top_core_EC_mix_out_41_) );
  XOR2X1 U6881 ( .A(top_core_EC_mc_n484), .B(top_core_EC_mc_n485), .Y(
        top_core_EC_mc_n483) );
  XNOR2X1 U6882 ( .A(top_core_EC_mc_mix_in_4_42_), .B(top_core_EC_mc_n486), 
        .Y(top_core_EC_mc_n482) );
  XNOR2X1 U6883 ( .A(top_core_EC_mc_mix_in_4_42_), .B(top_core_EC_mc_n441), 
        .Y(top_core_EC_mc_n484) );
  OAI22X1 U6884 ( .A0(top_core_EC_mc_n472), .A1(n2484), .B0(n2380), .B1(
        top_core_EC_mc_n473), .Y(top_core_EC_mix_out_43_) );
  XOR2X1 U6885 ( .A(top_core_EC_mc_n474), .B(top_core_EC_mc_n475), .Y(
        top_core_EC_mc_n473) );
  XNOR2X1 U6886 ( .A(top_core_EC_mc_mix_in_2_43_), .B(top_core_EC_mc_n476), 
        .Y(top_core_EC_mc_n472) );
  XNOR2X1 U6887 ( .A(top_core_EC_mc_mix_in_2_43_), .B(top_core_EC_mc_n416), 
        .Y(top_core_EC_mc_n474) );
  OAI22X1 U6888 ( .A0(top_core_EC_mc_n467), .A1(n2484), .B0(n2380), .B1(
        top_core_EC_mc_n468), .Y(top_core_EC_mix_out_44_) );
  XOR2X1 U6889 ( .A(top_core_EC_mc_n469), .B(top_core_EC_mc_n470), .Y(
        top_core_EC_mc_n468) );
  XNOR2X1 U6890 ( .A(top_core_EC_mc_mix_in_8[46]), .B(top_core_EC_mc_n471), 
        .Y(top_core_EC_mc_n467) );
  XNOR2X1 U6891 ( .A(top_core_EC_mc_mix_in_8[46]), .B(top_core_EC_mc_n408), 
        .Y(top_core_EC_mc_n469) );
  NAND2X1 U6892 ( .A(n3447), .B(n3453), .Y(n13847) );
  NAND2X1 U6893 ( .A(n2846), .B(n2852), .Y(n16997) );
  NAND2X1 U6894 ( .A(n2604), .B(n2610), .Y(n18257) );
  NAND2X1 U6895 ( .A(n3206), .B(n3212), .Y(n15107) );
  NAND2X1 U6896 ( .A(n3145), .B(n3151), .Y(n15422) );
  NAND2X1 U6897 ( .A(n2543), .B(n2549), .Y(n18572) );
  NAND2X1 U6898 ( .A(n2907), .B(n2913), .Y(n16682) );
  NAND2X1 U6899 ( .A(n3267), .B(n3273), .Y(n14792) );
  NAND2X1 U6900 ( .A(n2968), .B(n2974), .Y(n16367) );
  NAND2X1 U6901 ( .A(n2665), .B(n2671), .Y(n17942) );
  NAND2X1 U6902 ( .A(n3328), .B(n3334), .Y(n14477) );
  NAND2X1 U6903 ( .A(n3026), .B(n3032), .Y(n16052) );
  NAND2X1 U6904 ( .A(n2725), .B(n2731), .Y(n17627) );
  NAND2X1 U6905 ( .A(n3386), .B(n3392), .Y(n14162) );
  NAND2X1 U6906 ( .A(n3087), .B(n3093), .Y(n15737) );
  NAND2X1 U6907 ( .A(n2786), .B(n2792), .Y(n17312) );
  NAND2X1 U6908 ( .A(n633), .B(n2872), .Y(n17162) );
  NAND2X1 U6909 ( .A(n634), .B(n3473), .Y(n14012) );
  NAND2X1 U6910 ( .A(n635), .B(n2630), .Y(n18422) );
  NAND2X1 U6911 ( .A(n636), .B(n3232), .Y(n15272) );
  NAND2X1 U6912 ( .A(n637), .B(n3171), .Y(n15587) );
  NAND2X1 U6913 ( .A(n639), .B(n2933), .Y(n16847) );
  NAND2X1 U6914 ( .A(n638), .B(n2569), .Y(n18737) );
  NAND2X1 U6915 ( .A(n641), .B(n2994), .Y(n16532) );
  NAND2X1 U6916 ( .A(n642), .B(n2691), .Y(n18107) );
  NAND2X1 U6917 ( .A(n643), .B(n3354), .Y(n14642) );
  NAND2X1 U6918 ( .A(n644), .B(n3052), .Y(n16217) );
  NAND2X1 U6919 ( .A(n645), .B(n2751), .Y(n17792) );
  NAND2X1 U6920 ( .A(n646), .B(n3412), .Y(n14327) );
  NAND2X1 U6921 ( .A(n647), .B(n3113), .Y(n15902) );
  NAND2X1 U6922 ( .A(n648), .B(n2812), .Y(n17477) );
  NAND2X1 U6923 ( .A(n640), .B(n3293), .Y(n14957) );
  NAND2X1 U6924 ( .A(n634), .B(n6118), .Y(n13881) );
  NAND2X1 U6925 ( .A(n633), .B(n5335), .Y(n17031) );
  NAND2X1 U6926 ( .A(n635), .B(n4981), .Y(n18291) );
  NAND2X1 U6927 ( .A(n636), .B(n5807), .Y(n15141) );
  NAND2X1 U6928 ( .A(n637), .B(n5723), .Y(n15456) );
  NAND2X1 U6929 ( .A(n639), .B(n5419), .Y(n16716) );
  NAND2X1 U6930 ( .A(n638), .B(n4865), .Y(n18606) );
  NAND2X1 U6931 ( .A(n640), .B(n5883), .Y(n14826) );
  NAND2X1 U6932 ( .A(n641), .B(n5495), .Y(n16401) );
  NAND2X1 U6933 ( .A(n642), .B(n5065), .Y(n17976) );
  NAND2X1 U6934 ( .A(n643), .B(n5959), .Y(n14511) );
  NAND2X1 U6935 ( .A(n644), .B(n5571), .Y(n16086) );
  NAND2X1 U6936 ( .A(n645), .B(n5173), .Y(n17661) );
  NAND2X1 U6937 ( .A(n646), .B(n6035), .Y(n14196) );
  NAND2X1 U6938 ( .A(n647), .B(n5647), .Y(n15771) );
  NAND2X1 U6939 ( .A(n648), .B(n5251), .Y(n17346) );
  NAND2X1 U6940 ( .A(n15), .B(n9887), .Y(n9906) );
  NAND2X1 U6941 ( .A(n14), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n69), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n89) );
  NAND2X1 U6942 ( .A(n17), .B(n8135), .Y(n8154) );
  NAND2X1 U6943 ( .A(n16), .B(n11055), .Y(n11074) );
  NAND2X1 U6944 ( .A(n18), .B(n10763), .Y(n10782) );
  NAND2X1 U6945 ( .A(n20), .B(n7259), .Y(n7278) );
  NAND2X1 U6946 ( .A(n19), .B(n9011), .Y(n9030) );
  NAND2X1 U6947 ( .A(n21), .B(n10179), .Y(n10198) );
  NAND2X1 U6948 ( .A(n22), .B(n9303), .Y(n9322) );
  NAND2X1 U6949 ( .A(n23), .B(n8427), .Y(n8446) );
  NAND2X1 U6950 ( .A(n24), .B(n7551), .Y(n7570) );
  NAND2X1 U6951 ( .A(n25), .B(n11347), .Y(n11366) );
  NAND2X1 U6952 ( .A(n26), .B(n10471), .Y(n10490) );
  NAND2X1 U6953 ( .A(n27), .B(n9595), .Y(n9614) );
  NAND2X1 U6954 ( .A(n28), .B(n8719), .Y(n8738) );
  NAND2X1 U6955 ( .A(n29), .B(n7843), .Y(n7862) );
  XNOR2X1 U6956 ( .A(top_core_EC_mc_n850), .B(top_core_EC_mc_n851), .Y(
        top_core_EC_mc_n585) );
  XNOR2X1 U6957 ( .A(top_core_EC_mc_mix_in_8[18]), .B(
        top_core_EC_mc_mix_in_8[10]), .Y(top_core_EC_mc_n850) );
  XOR2X1 U6958 ( .A(top_core_EC_mc_mix_in_8[2]), .B(
        top_core_EC_mc_mix_in_8[26]), .Y(top_core_EC_mc_n851) );
  XNOR2X1 U6959 ( .A(top_core_EC_mc_n703), .B(top_core_EC_mc_n704), .Y(
        top_core_EC_mc_n344) );
  XNOR2X1 U6960 ( .A(top_core_EC_mc_mix_in_8[21]), .B(
        top_core_EC_mc_mix_in_8[13]), .Y(top_core_EC_mc_n703) );
  XOR2X1 U6961 ( .A(top_core_EC_mc_mix_in_8[5]), .B(
        top_core_EC_mc_mix_in_8[29]), .Y(top_core_EC_mc_n704) );
  XNOR2X1 U6962 ( .A(top_core_EC_mc_n696), .B(top_core_EC_mc_n697), .Y(
        top_core_EC_mc_n255) );
  XNOR2X1 U6963 ( .A(top_core_EC_mc_mix_in_8[22]), .B(
        top_core_EC_mc_mix_in_8[14]), .Y(top_core_EC_mc_n696) );
  XOR2X1 U6964 ( .A(top_core_EC_mc_mix_in_8[6]), .B(
        top_core_EC_mc_mix_in_8[30]), .Y(top_core_EC_mc_n697) );
  AOI31X1 U6965 ( .A0(n2893), .A1(n2867), .A2(n17008), .B0(n17189), .Y(n17180)
         );
  AOI31X1 U6966 ( .A0(n3494), .A1(n3468), .A2(n13858), .B0(n14039), .Y(n14030)
         );
  AOI31X1 U6967 ( .A0(n2650), .A1(n2625), .A2(n18268), .B0(n18449), .Y(n18440)
         );
  AOI31X1 U6968 ( .A0(n3253), .A1(n3227), .A2(n15118), .B0(n15299), .Y(n15290)
         );
  AOI31X1 U6969 ( .A0(n3192), .A1(n3166), .A2(n15433), .B0(n15614), .Y(n15605)
         );
  AOI31X1 U6970 ( .A0(n2954), .A1(n2928), .A2(n16693), .B0(n16874), .Y(n16865)
         );
  AOI31X1 U6971 ( .A0(n2600), .A1(n2564), .A2(n18583), .B0(n18764), .Y(n18755)
         );
  AOI31X1 U6972 ( .A0(n3314), .A1(n3288), .A2(n14803), .B0(n14984), .Y(n14975)
         );
  AOI31X1 U6973 ( .A0(n3015), .A1(n2989), .A2(n16378), .B0(n16559), .Y(n16550)
         );
  AOI31X1 U6974 ( .A0(n2711), .A1(n2686), .A2(n17953), .B0(n18134), .Y(n18125)
         );
  AOI31X1 U6975 ( .A0(n3375), .A1(n3349), .A2(n14488), .B0(n14669), .Y(n14660)
         );
  AOI31X1 U6976 ( .A0(n3072), .A1(n3047), .A2(n16063), .B0(n16244), .Y(n16235)
         );
  AOI31X1 U6977 ( .A0(n2772), .A1(n2746), .A2(n17638), .B0(n17819), .Y(n17810)
         );
  AOI31X1 U6978 ( .A0(n3433), .A1(n3407), .A2(n14173), .B0(n14354), .Y(n14345)
         );
  AOI31X1 U6979 ( .A0(n3134), .A1(n3108), .A2(n15748), .B0(n15929), .Y(n15920)
         );
  AOI31X1 U6980 ( .A0(n2833), .A1(n2807), .A2(n17323), .B0(n17504), .Y(n17495)
         );
  AOI22X1 U6981 ( .A0(n2871), .A1(n513), .B0(n2873), .B1(n481), .Y(n10041) );
  AOI22X1 U6982 ( .A0(n3472), .A1(n514), .B0(n3475), .B1(n482), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n227) );
  AOI22X1 U6983 ( .A0(n2629), .A1(n515), .B0(n2631), .B1(n483), .Y(n11209) );
  AOI22X1 U6984 ( .A0(n3231), .A1(n516), .B0(n3234), .B1(n484), .Y(n8289) );
  AOI22X1 U6985 ( .A0(n2690), .A1(n522), .B0(n2692), .B1(n485), .Y(n10917) );
  AOI22X1 U6986 ( .A0(n3051), .A1(n524), .B0(n3053), .B1(n486), .Y(n9165) );
  AOI22X1 U6987 ( .A0(n3411), .A1(n526), .B0(n3413), .B1(n487), .Y(n7413) );
  AOI22X1 U6988 ( .A0(n2811), .A1(n528), .B0(n2813), .B1(n488), .Y(n10333) );
  AOI22X1 U6989 ( .A0(n2993), .A1(n521), .B0(n2995), .B1(n489), .Y(n9457) );
  AOI22X1 U6990 ( .A0(n3170), .A1(n517), .B0(n3173), .B1(n490), .Y(n8581) );
  AOI22X1 U6991 ( .A0(n3353), .A1(n523), .B0(n3356), .B1(n491), .Y(n7705) );
  AOI22X1 U6992 ( .A0(n2568), .A1(n518), .B0(n2570), .B1(n492), .Y(n11501) );
  AOI22X1 U6993 ( .A0(n2750), .A1(n525), .B0(n2753), .B1(n493), .Y(n10625) );
  AOI22X1 U6994 ( .A0(n2932), .A1(n519), .B0(n2934), .B1(n494), .Y(n9749) );
  AOI22X1 U6995 ( .A0(n3112), .A1(n527), .B0(n3114), .B1(n495), .Y(n8873) );
  AOI22X1 U6996 ( .A0(n3292), .A1(n520), .B0(n3294), .B1(n496), .Y(n7997) );
  NOR4BX1 U6997 ( .AN(n17293), .B(n17294), .C(n5380), .D(n17037), .Y(n17291)
         );
  OAI221XL U6998 ( .A0(n1002), .A1(n17208), .B0(n2899), .B1(n30), .C0(n17295), 
        .Y(n17294) );
  AOI22X1 U6999 ( .A0(n401), .A1(n997), .B0(n5362), .B1(n2884), .Y(n17295) );
  NOR4BX1 U7000 ( .AN(n14143), .B(n14144), .C(n6151), .D(n13887), .Y(n14141)
         );
  OAI221XL U7001 ( .A0(n1141), .A1(n14058), .B0(n3499), .B1(n31), .C0(n14145), 
        .Y(n14144) );
  AOI22X1 U7002 ( .A0(n402), .A1(n1136), .B0(n6130), .B1(n3489), .Y(n14145) );
  NOR4BX1 U7003 ( .AN(n15403), .B(n15404), .C(n5852), .D(n15147), .Y(n15401)
         );
  OAI221XL U7004 ( .A0(n1086), .A1(n15318), .B0(n3259), .B1(n33), .C0(n15405), 
        .Y(n15404) );
  AOI22X1 U7005 ( .A0(n404), .A1(n1081), .B0(n5834), .B1(n3243), .Y(n15405) );
  NOR4BX1 U7006 ( .AN(n18553), .B(n18554), .C(n5026), .D(n18297), .Y(n18551)
         );
  OAI221XL U7007 ( .A0(n946), .A1(n18468), .B0(n2656), .B1(n32), .C0(n18555), 
        .Y(n18554) );
  AOI22X1 U7008 ( .A0(n403), .A1(n941), .B0(n5008), .B1(n2641), .Y(n18555) );
  NOR4BX1 U7009 ( .AN(n15718), .B(n15719), .C(n5768), .D(n15462), .Y(n15716)
         );
  OAI221XL U7010 ( .A0(n1072), .A1(n15633), .B0(n3198), .B1(n34), .C0(n15720), 
        .Y(n15719) );
  AOI22X1 U7011 ( .A0(n410), .A1(n1067), .B0(n5750), .B1(n3190), .Y(n15720) );
  NOR4BX1 U7012 ( .AN(n16978), .B(n16979), .C(n5464), .D(n16722), .Y(n16976)
         );
  OAI221XL U7013 ( .A0(n1016), .A1(n16893), .B0(n2960), .B1(n36), .C0(n16980), 
        .Y(n16979) );
  AOI22X1 U7014 ( .A0(n414), .A1(n1011), .B0(n5446), .B1(n2951), .Y(n16980) );
  NOR4BX1 U7015 ( .AN(n18868), .B(n18869), .C(n4910), .D(n18612), .Y(n18866)
         );
  OAI221XL U7016 ( .A0(n932), .A1(n18783), .B0(n2595), .B1(n35), .C0(n18870), 
        .Y(n18869) );
  AOI22X1 U7017 ( .A0(n412), .A1(n927), .B0(n4892), .B1(n2588), .Y(n18870) );
  NOR4BX1 U7018 ( .AN(n15088), .B(n15089), .C(n5928), .D(n14832), .Y(n15086)
         );
  OAI221XL U7019 ( .A0(n1100), .A1(n15003), .B0(n3322), .B1(n37), .C0(n15090), 
        .Y(n15089) );
  AOI22X1 U7020 ( .A0(n416), .A1(n1095), .B0(n5910), .B1(n3304), .Y(n15090) );
  NOR4BX1 U7021 ( .AN(n16663), .B(n16664), .C(n5540), .D(n16407), .Y(n16661)
         );
  OAI221XL U7022 ( .A0(n1030), .A1(n16578), .B0(n3020), .B1(n38), .C0(n16665), 
        .Y(n16664) );
  AOI22X1 U7023 ( .A0(n409), .A1(n1025), .B0(n5522), .B1(n3005), .Y(n16665) );
  NOR4BX1 U7024 ( .AN(n18238), .B(n18239), .C(n5110), .D(n17982), .Y(n18236)
         );
  OAI221XL U7025 ( .A0(n960), .A1(n18153), .B0(n2717), .B1(n39), .C0(n18240), 
        .Y(n18239) );
  AOI22X1 U7026 ( .A0(n405), .A1(n955), .B0(n5092), .B1(n2709), .Y(n18240) );
  NOR4BX1 U7027 ( .AN(n14773), .B(n14774), .C(n6004), .D(n14517), .Y(n14771)
         );
  OAI221XL U7028 ( .A0(n1114), .A1(n14688), .B0(n3380), .B1(n40), .C0(n14775), 
        .Y(n14774) );
  AOI22X1 U7029 ( .A0(n411), .A1(n1109), .B0(n5986), .B1(n3373), .Y(n14775) );
  NOR4BX1 U7030 ( .AN(n16348), .B(n16349), .C(n5616), .D(n16092), .Y(n16346)
         );
  OAI221XL U7031 ( .A0(n1044), .A1(n16263), .B0(n3078), .B1(n41), .C0(n16350), 
        .Y(n16349) );
  AOI22X1 U7032 ( .A0(n406), .A1(n1039), .B0(n5598), .B1(n3066), .Y(n16350) );
  NOR4BX1 U7033 ( .AN(n17923), .B(n17924), .C(n5218), .D(n17667), .Y(n17921)
         );
  OAI221XL U7034 ( .A0(n974), .A1(n17838), .B0(n2776), .B1(n42), .C0(n17925), 
        .Y(n17924) );
  AOI22X1 U7035 ( .A0(n413), .A1(n969), .B0(n5200), .B1(n2770), .Y(n17925) );
  NOR4BX1 U7036 ( .AN(n14458), .B(n14459), .C(n6080), .D(n14202), .Y(n14456)
         );
  OAI221XL U7037 ( .A0(n1128), .A1(n14373), .B0(n3439), .B1(n43), .C0(n14460), 
        .Y(n14459) );
  AOI22X1 U7038 ( .A0(n407), .A1(n1123), .B0(n6062), .B1(n3423), .Y(n14460) );
  NOR4BX1 U7039 ( .AN(n16033), .B(n16034), .C(n5692), .D(n15777), .Y(n16031)
         );
  OAI221XL U7040 ( .A0(n1058), .A1(n15948), .B0(n3139), .B1(n44), .C0(n16035), 
        .Y(n16034) );
  AOI22X1 U7041 ( .A0(n415), .A1(n1053), .B0(n5674), .B1(n3132), .Y(n16035) );
  NOR4BX1 U7042 ( .AN(n17608), .B(n17609), .C(n5296), .D(n17352), .Y(n17606)
         );
  OAI221XL U7043 ( .A0(n988), .A1(n17523), .B0(n2842), .B1(n45), .C0(n17610), 
        .Y(n17609) );
  AOI22X1 U7044 ( .A0(n408), .A1(n983), .B0(n5278), .B1(n2826), .Y(n17610) );
  NOR4X1 U7045 ( .A(n5340), .B(n10033), .C(n10034), .D(n10004), .Y(n10028) );
  AOI21XL U7046 ( .A0(n9888), .A1(n9896), .B0(n9913), .Y(n10034) );
  NOR4X1 U7047 ( .A(n6136), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n219), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n220), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n190), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n214) );
  AOI21XL U7048 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n70), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n220) );
  NOR4X1 U7049 ( .A(n4986), .B(n11201), .C(n11202), .D(n11172), .Y(n11196) );
  AOI21XL U7050 ( .A0(n11056), .A1(n11064), .B0(n11081), .Y(n11202) );
  NOR4X1 U7051 ( .A(n5812), .B(n8281), .C(n8282), .D(n8252), .Y(n8276) );
  AOI21XL U7052 ( .A0(n8136), .A1(n8144), .B0(n8161), .Y(n8282) );
  NOR4X1 U7053 ( .A(n5070), .B(n10909), .C(n10910), .D(n10880), .Y(n10904) );
  AOI21XL U7054 ( .A0(n10764), .A1(n10772), .B0(n10789), .Y(n10910) );
  NOR4X1 U7055 ( .A(n5576), .B(n9157), .C(n9158), .D(n9128), .Y(n9152) );
  AOI21XL U7056 ( .A0(n9012), .A1(n9020), .B0(n9037), .Y(n9158) );
  NOR4X1 U7057 ( .A(n6040), .B(n7405), .C(n7406), .D(n7376), .Y(n7400) );
  AOI21XL U7058 ( .A0(n7260), .A1(n7268), .B0(n7285), .Y(n7406) );
  NOR4X1 U7059 ( .A(n5256), .B(n10325), .C(n10326), .D(n10296), .Y(n10320) );
  AOI21XL U7060 ( .A0(n10180), .A1(n10188), .B0(n10205), .Y(n10326) );
  NOR4X1 U7061 ( .A(n5500), .B(n9449), .C(n9450), .D(n9420), .Y(n9444) );
  AOI21XL U7062 ( .A0(n9304), .A1(n9312), .B0(n9329), .Y(n9450) );
  NOR4X1 U7063 ( .A(n5728), .B(n8573), .C(n8574), .D(n8544), .Y(n8568) );
  AOI21XL U7064 ( .A0(n8428), .A1(n8436), .B0(n8453), .Y(n8574) );
  NOR4X1 U7065 ( .A(n5964), .B(n7697), .C(n7698), .D(n7668), .Y(n7692) );
  AOI21XL U7066 ( .A0(n7552), .A1(n7560), .B0(n7577), .Y(n7698) );
  NOR4X1 U7067 ( .A(n4870), .B(n11493), .C(n11494), .D(n11464), .Y(n11488) );
  AOI21XL U7068 ( .A0(n11348), .A1(n11356), .B0(n11373), .Y(n11494) );
  NOR4X1 U7069 ( .A(n5178), .B(n10617), .C(n10618), .D(n10588), .Y(n10612) );
  AOI21XL U7070 ( .A0(n10472), .A1(n10480), .B0(n10497), .Y(n10618) );
  NOR4X1 U7071 ( .A(n5424), .B(n9741), .C(n9742), .D(n9712), .Y(n9736) );
  AOI21XL U7072 ( .A0(n9596), .A1(n9604), .B0(n9621), .Y(n9742) );
  NOR4X1 U7073 ( .A(n5652), .B(n8865), .C(n8866), .D(n8836), .Y(n8860) );
  AOI21XL U7074 ( .A0(n8720), .A1(n8728), .B0(n8745), .Y(n8866) );
  NOR4X1 U7075 ( .A(n5888), .B(n7989), .C(n7990), .D(n7960), .Y(n7984) );
  AOI21XL U7076 ( .A0(n7844), .A1(n7852), .B0(n7869), .Y(n7990) );
  NAND2X1 U7077 ( .A(n6549), .B(n13238), .Y(n13333) );
  NAND2X1 U7078 ( .A(n6844), .B(n12608), .Y(n12703) );
  NAND2X1 U7079 ( .A(n6890), .B(n12923), .Y(n13018) );
  NAND2X1 U7080 ( .A(n2846), .B(n2852), .Y(n9992) );
  NAND2X1 U7081 ( .A(n3447), .B(n3453), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n178) );
  NAND2X1 U7082 ( .A(n2604), .B(n2610), .Y(n11160) );
  NAND2X1 U7083 ( .A(n3206), .B(n3212), .Y(n8240) );
  NAND2X1 U7084 ( .A(n2665), .B(n2671), .Y(n10868) );
  NAND2X1 U7085 ( .A(n3026), .B(n3032), .Y(n9116) );
  NAND2X1 U7086 ( .A(n3386), .B(n3392), .Y(n7364) );
  NAND2X1 U7087 ( .A(n2786), .B(n2792), .Y(n10284) );
  NAND2X1 U7088 ( .A(n2968), .B(n2974), .Y(n9408) );
  NAND2X1 U7089 ( .A(n3145), .B(n3151), .Y(n8532) );
  NAND2X1 U7090 ( .A(n3328), .B(n3334), .Y(n7656) );
  NAND2X1 U7091 ( .A(n2543), .B(n2549), .Y(n11452) );
  NAND2X1 U7092 ( .A(n2725), .B(n2731), .Y(n10576) );
  NAND2X1 U7093 ( .A(n2907), .B(n2913), .Y(n9700) );
  NAND2X1 U7094 ( .A(n3087), .B(n3093), .Y(n8824) );
  NAND2X1 U7095 ( .A(n3267), .B(n3273), .Y(n7948) );
  NAND2X1 U7096 ( .A(n3447), .B(n3458), .Y(n13937) );
  NAND2X1 U7097 ( .A(n2846), .B(n2857), .Y(n17087) );
  NAND2X1 U7098 ( .A(n2604), .B(n2615), .Y(n18347) );
  NAND2X1 U7099 ( .A(n3206), .B(n3217), .Y(n15197) );
  NAND2X1 U7100 ( .A(n3145), .B(n3156), .Y(n15512) );
  NAND2X1 U7101 ( .A(n2543), .B(n2554), .Y(n18662) );
  NAND2X1 U7102 ( .A(n2907), .B(n2918), .Y(n16772) );
  NAND2X1 U7103 ( .A(n3267), .B(n3278), .Y(n14882) );
  NAND2X1 U7104 ( .A(n2968), .B(n2979), .Y(n16457) );
  NAND2X1 U7105 ( .A(n2665), .B(n2676), .Y(n18032) );
  NAND2X1 U7106 ( .A(n3328), .B(n3339), .Y(n14567) );
  NAND2X1 U7107 ( .A(n3026), .B(n3037), .Y(n16142) );
  NAND2X1 U7108 ( .A(n2725), .B(n2736), .Y(n17717) );
  NAND2X1 U7109 ( .A(n3386), .B(n3397), .Y(n14252) );
  NAND2X1 U7110 ( .A(n3087), .B(n3098), .Y(n15827) );
  NAND2X1 U7111 ( .A(n2786), .B(n2797), .Y(n17402) );
  AOI31X1 U7112 ( .A0(n3468), .A1(n6167), .A2(n1142), .B0(n13849), .Y(n13844)
         );
  AOI31X1 U7113 ( .A0(n2867), .A1(n5385), .A2(n1003), .B0(n16999), .Y(n16994)
         );
  AOI31X1 U7114 ( .A0(n2625), .A1(n5031), .A2(n947), .B0(n18259), .Y(n18254)
         );
  AOI31X1 U7115 ( .A0(n3227), .A1(n5857), .A2(n1087), .B0(n15109), .Y(n15104)
         );
  AOI31X1 U7116 ( .A0(n3166), .A1(n5773), .A2(n1073), .B0(n15424), .Y(n15419)
         );
  AOI31X1 U7117 ( .A0(n2564), .A1(n4915), .A2(n933), .B0(n18574), .Y(n18569)
         );
  AOI31X1 U7118 ( .A0(n2928), .A1(n5469), .A2(n1017), .B0(n16684), .Y(n16679)
         );
  AOI31X1 U7119 ( .A0(n3288), .A1(n5933), .A2(n1101), .B0(n14794), .Y(n14789)
         );
  AOI31X1 U7120 ( .A0(n2989), .A1(n5545), .A2(n1031), .B0(n16369), .Y(n16364)
         );
  AOI31X1 U7121 ( .A0(n2686), .A1(n5115), .A2(n961), .B0(n17944), .Y(n17939)
         );
  AOI31X1 U7122 ( .A0(n3349), .A1(n6009), .A2(n1115), .B0(n14479), .Y(n14474)
         );
  AOI31X1 U7123 ( .A0(n3047), .A1(n5621), .A2(n1045), .B0(n16054), .Y(n16049)
         );
  AOI31X1 U7124 ( .A0(n2746), .A1(n5223), .A2(n975), .B0(n17629), .Y(n17624)
         );
  AOI31X1 U7125 ( .A0(n3407), .A1(n6085), .A2(n1129), .B0(n14164), .Y(n14159)
         );
  AOI31X1 U7126 ( .A0(n3108), .A1(n5697), .A2(n1059), .B0(n15739), .Y(n15734)
         );
  AOI31X1 U7127 ( .A0(n2807), .A1(n5301), .A2(n989), .B0(n17314), .Y(n17309)
         );
  NOR2XL U7128 ( .A(n165), .B(n3493), .Y(n14085) );
  NOR2XL U7129 ( .A(n164), .B(n2892), .Y(n17235) );
  NOR2XL U7130 ( .A(n166), .B(n2651), .Y(n18495) );
  NOR2XL U7131 ( .A(n167), .B(n3252), .Y(n15345) );
  NOR2XL U7132 ( .A(n169), .B(n2589), .Y(n18810) );
  NOR2XL U7133 ( .A(n168), .B(n3191), .Y(n15660) );
  NOR2XL U7134 ( .A(n170), .B(n2953), .Y(n16920) );
  NOR2XL U7135 ( .A(n171), .B(n3313), .Y(n15030) );
  NOR2XL U7136 ( .A(n172), .B(n3014), .Y(n16605) );
  NOR2XL U7137 ( .A(n173), .B(n2710), .Y(n18180) );
  NOR2XL U7138 ( .A(n174), .B(n3374), .Y(n14715) );
  NOR2XL U7139 ( .A(n175), .B(n3073), .Y(n16290) );
  NOR2XL U7140 ( .A(n176), .B(n2771), .Y(n17865) );
  NOR2XL U7141 ( .A(n177), .B(n3432), .Y(n14400) );
  NOR2XL U7142 ( .A(n178), .B(n3133), .Y(n15975) );
  NOR2XL U7143 ( .A(n179), .B(n2832), .Y(n17550) );
  NOR2X1 U7144 ( .A(n586), .B(n5384), .Y(n9998) );
  NOR2X1 U7145 ( .A(n585), .B(n6169), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n184) );
  NOR2X1 U7146 ( .A(n588), .B(n5856), .Y(n8246) );
  NOR2X1 U7147 ( .A(n587), .B(n5030), .Y(n11166) );
  NOR2X1 U7148 ( .A(n589), .B(n5114), .Y(n10874) );
  NOR2X1 U7149 ( .A(n591), .B(n6084), .Y(n7370) );
  NOR2X1 U7150 ( .A(n590), .B(n5620), .Y(n9122) );
  NOR2X1 U7151 ( .A(n592), .B(n5300), .Y(n10290) );
  NOR2X1 U7152 ( .A(n593), .B(n5544), .Y(n9414) );
  NOR2X1 U7153 ( .A(n594), .B(n5772), .Y(n8538) );
  NOR2X1 U7154 ( .A(n595), .B(n6008), .Y(n7662) );
  NOR2X1 U7155 ( .A(n596), .B(n4914), .Y(n11458) );
  NOR2X1 U7156 ( .A(n597), .B(n5222), .Y(n10582) );
  NOR2X1 U7157 ( .A(n598), .B(n5468), .Y(n9706) );
  NOR2X1 U7158 ( .A(n599), .B(n5696), .Y(n8830) );
  NOR2X1 U7159 ( .A(n600), .B(n5932), .Y(n7954) );
  NAND2X1 U7160 ( .A(n3493), .B(n634), .Y(n13856) );
  NAND2X1 U7161 ( .A(n2892), .B(n633), .Y(n17006) );
  NAND2X1 U7162 ( .A(n2661), .B(n635), .Y(n18266) );
  NAND2X1 U7163 ( .A(n3252), .B(n636), .Y(n15116) );
  NAND2X1 U7164 ( .A(n3191), .B(n637), .Y(n15431) );
  NAND2X1 U7165 ( .A(n2589), .B(n638), .Y(n18581) );
  NAND2X1 U7166 ( .A(n2953), .B(n639), .Y(n16691) );
  NAND2X1 U7167 ( .A(n3313), .B(n640), .Y(n14801) );
  NAND2X1 U7168 ( .A(n3014), .B(n641), .Y(n16376) );
  NAND2X1 U7169 ( .A(n2710), .B(n642), .Y(n17951) );
  NAND2X1 U7170 ( .A(n3374), .B(n643), .Y(n14486) );
  NAND2X1 U7171 ( .A(n3083), .B(n644), .Y(n16061) );
  NAND2X1 U7172 ( .A(n2771), .B(n645), .Y(n17636) );
  NAND2X1 U7173 ( .A(n3432), .B(n646), .Y(n14171) );
  NAND2X1 U7174 ( .A(n3133), .B(n647), .Y(n15746) );
  NAND2X1 U7175 ( .A(n2832), .B(n648), .Y(n17321) );
  NAND2X1 U7176 ( .A(n465), .B(n5363), .Y(n17036) );
  NAND2X1 U7177 ( .A(n466), .B(n6131), .Y(n13886) );
  NAND2X1 U7178 ( .A(n468), .B(n5835), .Y(n15146) );
  NAND2X1 U7179 ( .A(n467), .B(n5009), .Y(n18296) );
  NAND2X1 U7180 ( .A(n469), .B(n5751), .Y(n15461) );
  NAND2X1 U7181 ( .A(n470), .B(n5447), .Y(n16721) );
  NAND2X1 U7182 ( .A(n471), .B(n4893), .Y(n18611) );
  NAND2X1 U7183 ( .A(n472), .B(n5911), .Y(n14831) );
  NAND2X1 U7184 ( .A(n473), .B(n5523), .Y(n16406) );
  NAND2X1 U7185 ( .A(n474), .B(n5093), .Y(n17981) );
  NAND2X1 U7186 ( .A(n475), .B(n5987), .Y(n14516) );
  NAND2X1 U7187 ( .A(n476), .B(n5599), .Y(n16091) );
  NAND2X1 U7188 ( .A(n477), .B(n5201), .Y(n17666) );
  NAND2X1 U7189 ( .A(n478), .B(n6063), .Y(n14201) );
  NAND2X1 U7190 ( .A(n479), .B(n5675), .Y(n15776) );
  NAND2X1 U7191 ( .A(n480), .B(n5279), .Y(n17351) );
  NAND2X1 U7192 ( .A(n2851), .B(n2849), .Y(n17056) );
  NAND2X1 U7193 ( .A(n3452), .B(n3449), .Y(n13906) );
  NAND2X1 U7194 ( .A(n2609), .B(n2607), .Y(n18316) );
  NAND2X1 U7195 ( .A(n3211), .B(n3209), .Y(n15166) );
  NAND2X1 U7196 ( .A(n3150), .B(n3148), .Y(n15481) );
  NAND2X1 U7197 ( .A(n2912), .B(n2910), .Y(n16741) );
  NAND2X1 U7198 ( .A(n2548), .B(n2546), .Y(n18631) );
  NAND2X1 U7199 ( .A(n3272), .B(n3270), .Y(n14851) );
  NAND2X1 U7200 ( .A(n2973), .B(n2971), .Y(n16426) );
  NAND2X1 U7201 ( .A(n2670), .B(n2668), .Y(n18001) );
  NAND2X1 U7202 ( .A(n3333), .B(n3331), .Y(n14536) );
  NAND2X1 U7203 ( .A(n3031), .B(n3029), .Y(n16111) );
  NAND2X1 U7204 ( .A(n2730), .B(n2728), .Y(n17686) );
  NAND2X1 U7205 ( .A(n3391), .B(n3389), .Y(n14221) );
  NAND2X1 U7206 ( .A(n3092), .B(n3090), .Y(n15796) );
  NAND2X1 U7207 ( .A(n2791), .B(n2789), .Y(n17371) );
  NOR4X1 U7208 ( .A(n13871), .B(n13872), .C(n13873), .D(n13874), .Y(n13838) );
  OAI21XL U7209 ( .A0(n3481), .A1(n13881), .B0(n13882), .Y(n13872) );
  AOI31X1 U7210 ( .A0(n13875), .A1(n13876), .A2(n13877), .B0(n3463), .Y(n13874) );
  AOI31X1 U7211 ( .A0(n13878), .A1(n13879), .A2(n13856), .B0(n13880), .Y(
        n13873) );
  NOR4X1 U7212 ( .A(n17021), .B(n17022), .C(n17023), .D(n17024), .Y(n16988) );
  OAI21XL U7213 ( .A0(n2880), .A1(n17031), .B0(n17032), .Y(n17022) );
  AOI31X1 U7214 ( .A0(n17025), .A1(n17026), .A2(n17027), .B0(n2861), .Y(n17024) );
  AOI31X1 U7215 ( .A0(n17028), .A1(n17029), .A2(n17006), .B0(n17030), .Y(
        n17023) );
  NOR4X1 U7216 ( .A(n18281), .B(n18282), .C(n18283), .D(n18284), .Y(n18248) );
  OAI21XL U7217 ( .A0(n2638), .A1(n18291), .B0(n18292), .Y(n18282) );
  AOI31X1 U7218 ( .A0(n18285), .A1(n18286), .A2(n18287), .B0(n2612), .Y(n18284) );
  AOI31X1 U7219 ( .A0(n18288), .A1(n18289), .A2(n18266), .B0(n18290), .Y(
        n18283) );
  NOR4X1 U7220 ( .A(n15131), .B(n15132), .C(n15133), .D(n15134), .Y(n15098) );
  OAI21XL U7221 ( .A0(n3240), .A1(n15141), .B0(n15142), .Y(n15132) );
  AOI31X1 U7222 ( .A0(n15135), .A1(n15136), .A2(n15137), .B0(n3221), .Y(n15134) );
  AOI31X1 U7223 ( .A0(n15138), .A1(n15139), .A2(n15116), .B0(n15140), .Y(
        n15133) );
  NOR4X1 U7224 ( .A(n15446), .B(n15447), .C(n15448), .D(n15449), .Y(n15413) );
  OAI21XL U7225 ( .A0(n3179), .A1(n15456), .B0(n15457), .Y(n15447) );
  AOI31X1 U7226 ( .A0(n15450), .A1(n15451), .A2(n15452), .B0(n3153), .Y(n15449) );
  AOI31X1 U7227 ( .A0(n15453), .A1(n15454), .A2(n15431), .B0(n15455), .Y(
        n15448) );
  NOR4X1 U7228 ( .A(n18596), .B(n18597), .C(n18598), .D(n18599), .Y(n18563) );
  OAI21XL U7229 ( .A0(n2577), .A1(n18606), .B0(n18607), .Y(n18597) );
  AOI31X1 U7230 ( .A0(n18600), .A1(n18601), .A2(n18602), .B0(n2556), .Y(n18599) );
  AOI31X1 U7231 ( .A0(n18603), .A1(n18604), .A2(n18581), .B0(n18605), .Y(
        n18598) );
  NOR4X1 U7232 ( .A(n16706), .B(n16707), .C(n16708), .D(n16709), .Y(n16673) );
  OAI21XL U7233 ( .A0(n2941), .A1(n16716), .B0(n16717), .Y(n16707) );
  AOI31X1 U7234 ( .A0(n16710), .A1(n16711), .A2(n16712), .B0(n2915), .Y(n16709) );
  AOI31X1 U7235 ( .A0(n16713), .A1(n16714), .A2(n16691), .B0(n16715), .Y(
        n16708) );
  NOR4X1 U7236 ( .A(n14816), .B(n14817), .C(n14818), .D(n14819), .Y(n14783) );
  OAI21XL U7237 ( .A0(n3301), .A1(n14826), .B0(n14827), .Y(n14817) );
  AOI31X1 U7238 ( .A0(n14820), .A1(n14821), .A2(n14822), .B0(n3275), .Y(n14819) );
  AOI31X1 U7239 ( .A0(n14823), .A1(n14824), .A2(n14801), .B0(n14825), .Y(
        n14818) );
  NOR4X1 U7240 ( .A(n16391), .B(n16392), .C(n16393), .D(n16394), .Y(n16358) );
  OAI21XL U7241 ( .A0(n3002), .A1(n16401), .B0(n16402), .Y(n16392) );
  AOI31X1 U7242 ( .A0(n16395), .A1(n16396), .A2(n16397), .B0(n2976), .Y(n16394) );
  AOI31X1 U7243 ( .A0(n16398), .A1(n16399), .A2(n16376), .B0(n16400), .Y(
        n16393) );
  NOR4X1 U7244 ( .A(n17966), .B(n17967), .C(n17968), .D(n17969), .Y(n17933) );
  OAI21XL U7245 ( .A0(n2699), .A1(n17976), .B0(n17977), .Y(n17967) );
  AOI31X1 U7246 ( .A0(n17970), .A1(n17971), .A2(n17972), .B0(n2680), .Y(n17969) );
  AOI31X1 U7247 ( .A0(n17973), .A1(n17974), .A2(n17951), .B0(n17975), .Y(
        n17968) );
  NOR4X1 U7248 ( .A(n14501), .B(n14502), .C(n14503), .D(n14504), .Y(n14468) );
  OAI21XL U7249 ( .A0(n3362), .A1(n14511), .B0(n14512), .Y(n14502) );
  AOI31X1 U7250 ( .A0(n14505), .A1(n14506), .A2(n14507), .B0(n3336), .Y(n14504) );
  AOI31X1 U7251 ( .A0(n14508), .A1(n14509), .A2(n14486), .B0(n14510), .Y(
        n14503) );
  NOR4X1 U7252 ( .A(n16076), .B(n16077), .C(n16078), .D(n16079), .Y(n16043) );
  OAI21XL U7253 ( .A0(n3060), .A1(n16086), .B0(n16087), .Y(n16077) );
  AOI31X1 U7254 ( .A0(n16080), .A1(n16081), .A2(n16082), .B0(n3034), .Y(n16079) );
  AOI31X1 U7255 ( .A0(n16083), .A1(n16084), .A2(n16061), .B0(n16085), .Y(
        n16078) );
  NOR4X1 U7256 ( .A(n17651), .B(n17652), .C(n17653), .D(n17654), .Y(n17618) );
  OAI21XL U7257 ( .A0(n2759), .A1(n17661), .B0(n17662), .Y(n17652) );
  AOI31X1 U7258 ( .A0(n17655), .A1(n17656), .A2(n17657), .B0(n2740), .Y(n17654) );
  AOI31X1 U7259 ( .A0(n17658), .A1(n17659), .A2(n17636), .B0(n17660), .Y(
        n17653) );
  NOR4X1 U7260 ( .A(n14186), .B(n14187), .C(n14188), .D(n14189), .Y(n14153) );
  OAI21XL U7261 ( .A0(n3420), .A1(n14196), .B0(n14197), .Y(n14187) );
  AOI31X1 U7262 ( .A0(n14190), .A1(n14191), .A2(n14192), .B0(n3394), .Y(n14189) );
  AOI31X1 U7263 ( .A0(n14193), .A1(n14194), .A2(n14171), .B0(n14195), .Y(
        n14188) );
  NOR4X1 U7264 ( .A(n15761), .B(n15762), .C(n15763), .D(n15764), .Y(n15728) );
  OAI21XL U7265 ( .A0(n3121), .A1(n15771), .B0(n15772), .Y(n15762) );
  AOI31X1 U7266 ( .A0(n15765), .A1(n15766), .A2(n15767), .B0(n3102), .Y(n15764) );
  AOI31X1 U7267 ( .A0(n15768), .A1(n15769), .A2(n15746), .B0(n15770), .Y(
        n15763) );
  NOR4X1 U7268 ( .A(n17336), .B(n17337), .C(n17338), .D(n17339), .Y(n17303) );
  OAI21XL U7269 ( .A0(n2820), .A1(n17346), .B0(n17347), .Y(n17337) );
  AOI31X1 U7270 ( .A0(n17340), .A1(n17341), .A2(n17342), .B0(n2794), .Y(n17339) );
  AOI31X1 U7271 ( .A0(n17343), .A1(n17344), .A2(n17321), .B0(n17345), .Y(
        n17338) );
  OAI21XL U7272 ( .A0(n465), .A1(n9943), .B0(n90), .Y(n9964) );
  OAI21XL U7273 ( .A0(n466), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n128), 
        .B0(n91), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n149) );
  OAI21XL U7274 ( .A0(n467), .A1(n11111), .B0(n92), .Y(n11132) );
  OAI21XL U7275 ( .A0(n468), .A1(n8191), .B0(n93), .Y(n8212) );
  OAI21XL U7276 ( .A0(n474), .A1(n10819), .B0(n94), .Y(n10840) );
  OAI21XL U7277 ( .A0(n476), .A1(n9067), .B0(n96), .Y(n9088) );
  OAI21XL U7278 ( .A0(n478), .A1(n7315), .B0(n95), .Y(n7336) );
  OAI21XL U7279 ( .A0(n480), .A1(n10235), .B0(n97), .Y(n10256) );
  OAI21XL U7280 ( .A0(n473), .A1(n9359), .B0(n98), .Y(n9380) );
  OAI21XL U7281 ( .A0(n469), .A1(n8483), .B0(n99), .Y(n8504) );
  OAI21XL U7282 ( .A0(n475), .A1(n7607), .B0(n100), .Y(n7628) );
  OAI21XL U7283 ( .A0(n471), .A1(n11403), .B0(n101), .Y(n11424) );
  OAI21XL U7284 ( .A0(n477), .A1(n10527), .B0(n102), .Y(n10548) );
  OAI21XL U7285 ( .A0(n470), .A1(n9651), .B0(n103), .Y(n9672) );
  OAI21XL U7286 ( .A0(n479), .A1(n8775), .B0(n104), .Y(n8796) );
  OAI21XL U7287 ( .A0(n472), .A1(n7899), .B0(n105), .Y(n7920) );
  NAND2X1 U7288 ( .A(n1148), .B(n1172), .Y(n13225) );
  NAND2X1 U7289 ( .A(n1197), .B(n1218), .Y(n12910) );
  NAND2X1 U7290 ( .A(n1188), .B(n1212), .Y(n12595) );
  NOR2X1 U7291 ( .A(n13286), .B(n692), .Y(n13312) );
  NOR2X1 U7292 ( .A(n12656), .B(n694), .Y(n12682) );
  NOR2X1 U7293 ( .A(n12971), .B(n696), .Y(n12997) );
  AOI31X1 U7294 ( .A0(n17198), .A1(n17199), .A2(n17200), .B0(n17056), .Y(
        n17197) );
  AOI222X1 U7295 ( .A0(n17093), .A1(n633), .B0(n994), .B1(n2896), .C0(n401), 
        .C1(n998), .Y(n17200) );
  AOI22X1 U7296 ( .A0(n5357), .A1(n2892), .B0(n5353), .B1(n1005), .Y(n17198)
         );
  AOI31X1 U7297 ( .A0(n14048), .A1(n14049), .A2(n14050), .B0(n13906), .Y(
        n14047) );
  AOI222X1 U7298 ( .A0(n13943), .A1(n634), .B0(n1133), .B1(n3502), .C0(n402), 
        .C1(n1137), .Y(n14050) );
  AOI22X1 U7299 ( .A0(n6125), .A1(n3493), .B0(n6121), .B1(n1144), .Y(n14048)
         );
  AOI31X1 U7300 ( .A0(n18458), .A1(n18459), .A2(n18460), .B0(n18316), .Y(
        n18457) );
  AOI222X1 U7301 ( .A0(n18353), .A1(n635), .B0(n938), .B1(n2653), .C0(n403), 
        .C1(n942), .Y(n18460) );
  AOI22X1 U7302 ( .A0(n5003), .A1(top_core_EC_ss_in[112]), .B0(n4999), .B1(
        n949), .Y(n18458) );
  AOI31X1 U7303 ( .A0(n15308), .A1(n15309), .A2(n15310), .B0(n15166), .Y(
        n15307) );
  AOI222X1 U7304 ( .A0(n15203), .A1(n636), .B0(n1078), .B1(n3256), .C0(n404), 
        .C1(n1082), .Y(n15310) );
  AOI22X1 U7305 ( .A0(n5829), .A1(n3252), .B0(n5825), .B1(n1089), .Y(n15308)
         );
  AOI31X1 U7306 ( .A0(n15623), .A1(n15624), .A2(n15625), .B0(n15481), .Y(
        n15622) );
  AOI222X1 U7307 ( .A0(n15518), .A1(n637), .B0(n1064), .B1(n3195), .C0(n410), 
        .C1(n1068), .Y(n15625) );
  AOI22X1 U7308 ( .A0(n5745), .A1(n3191), .B0(n5741), .B1(n1075), .Y(n15623)
         );
  AOI31X1 U7309 ( .A0(n16883), .A1(n16884), .A2(n16885), .B0(n16741), .Y(
        n16882) );
  AOI222X1 U7310 ( .A0(n16778), .A1(n639), .B0(n1008), .B1(n2957), .C0(n414), 
        .C1(n1012), .Y(n16885) );
  AOI22X1 U7311 ( .A0(n5441), .A1(n2953), .B0(n5437), .B1(n1019), .Y(n16883)
         );
  AOI31X1 U7312 ( .A0(n18773), .A1(n18774), .A2(n18775), .B0(n18631), .Y(
        n18772) );
  AOI222X1 U7313 ( .A0(n18668), .A1(n638), .B0(n924), .B1(n2592), .C0(n412), 
        .C1(n928), .Y(n18775) );
  AOI22X1 U7314 ( .A0(n4887), .A1(n2589), .B0(n4883), .B1(n935), .Y(n18773) );
  AOI31X1 U7315 ( .A0(n14993), .A1(n14994), .A2(n14995), .B0(n14851), .Y(
        n14992) );
  AOI222X1 U7316 ( .A0(n14888), .A1(n640), .B0(n1092), .B1(n3316), .C0(n416), 
        .C1(n1096), .Y(n14995) );
  AOI22X1 U7317 ( .A0(n5905), .A1(n3313), .B0(n5901), .B1(n1103), .Y(n14993)
         );
  AOI31X1 U7318 ( .A0(n16568), .A1(n16569), .A2(n16570), .B0(n16426), .Y(
        n16567) );
  AOI222X1 U7319 ( .A0(n16463), .A1(n641), .B0(n1022), .B1(n3023), .C0(n409), 
        .C1(n1026), .Y(n16570) );
  AOI22X1 U7320 ( .A0(n5517), .A1(n3014), .B0(n5513), .B1(n1033), .Y(n16568)
         );
  AOI31X1 U7321 ( .A0(n18143), .A1(n18144), .A2(n18145), .B0(n18001), .Y(
        n18142) );
  AOI222X1 U7322 ( .A0(n18038), .A1(n642), .B0(n952), .B1(n2718), .C0(n405), 
        .C1(n956), .Y(n18145) );
  AOI22X1 U7323 ( .A0(n5087), .A1(n2710), .B0(n5083), .B1(n963), .Y(n18143) );
  AOI31X1 U7324 ( .A0(n14678), .A1(n14679), .A2(n14680), .B0(n14536), .Y(
        n14677) );
  AOI222X1 U7325 ( .A0(n14573), .A1(n643), .B0(n1106), .B1(n3383), .C0(n411), 
        .C1(n1110), .Y(n14680) );
  AOI22X1 U7326 ( .A0(n5981), .A1(n3374), .B0(n5977), .B1(n1117), .Y(n14678)
         );
  AOI31X1 U7327 ( .A0(n16253), .A1(n16254), .A2(n16255), .B0(n16111), .Y(
        n16252) );
  AOI222X1 U7328 ( .A0(n16148), .A1(n644), .B0(n1036), .B1(n3075), .C0(n406), 
        .C1(n1040), .Y(n16255) );
  AOI22X1 U7329 ( .A0(n5593), .A1(top_core_EC_ss_in[56]), .B0(n5589), .B1(
        n1047), .Y(n16253) );
  AOI31X1 U7330 ( .A0(n17828), .A1(n17829), .A2(n17830), .B0(n17686), .Y(
        n17827) );
  AOI222X1 U7331 ( .A0(n17723), .A1(n645), .B0(n966), .B1(n2782), .C0(n413), 
        .C1(n970), .Y(n17830) );
  AOI22X1 U7332 ( .A0(n5195), .A1(n2771), .B0(n5191), .B1(n977), .Y(n17828) );
  AOI31X1 U7333 ( .A0(n14363), .A1(n14364), .A2(n14365), .B0(n14221), .Y(
        n14362) );
  AOI222X1 U7334 ( .A0(n14258), .A1(n646), .B0(n1120), .B1(n3440), .C0(n407), 
        .C1(n1124), .Y(n14365) );
  AOI22X1 U7335 ( .A0(n6057), .A1(n3432), .B0(n6053), .B1(n1131), .Y(n14363)
         );
  AOI31X1 U7336 ( .A0(n15938), .A1(n15939), .A2(n15940), .B0(n15796), .Y(
        n15937) );
  AOI222X1 U7337 ( .A0(n15833), .A1(n647), .B0(n1050), .B1(n3142), .C0(n415), 
        .C1(n1054), .Y(n15940) );
  AOI22X1 U7338 ( .A0(n5669), .A1(n3133), .B0(n5665), .B1(n1061), .Y(n15938)
         );
  AOI31X1 U7339 ( .A0(n17513), .A1(n17514), .A2(n17515), .B0(n17371), .Y(
        n17512) );
  AOI222X1 U7340 ( .A0(n17408), .A1(n648), .B0(n980), .B1(n2843), .C0(n408), 
        .C1(n984), .Y(n17515) );
  AOI22X1 U7341 ( .A0(n5273), .A1(n2832), .B0(n5269), .B1(n991), .Y(n17513) );
  NOR2X1 U7342 ( .A(n6165), .B(n6166), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n255) );
  NOR2X1 U7343 ( .A(n5847), .B(n5848), .Y(n8317) );
  NOR2X1 U7344 ( .A(n5375), .B(n5376), .Y(n10069) );
  NOR2X1 U7345 ( .A(n5021), .B(n5022), .Y(n11237) );
  NOR2X1 U7346 ( .A(n5611), .B(n5612), .Y(n9193) );
  NOR2X1 U7347 ( .A(n5105), .B(n5106), .Y(n10945) );
  NOR2X1 U7348 ( .A(n6075), .B(n6076), .Y(n7441) );
  NOR2X1 U7349 ( .A(n5291), .B(n5292), .Y(n10361) );
  NOR2X1 U7350 ( .A(n5535), .B(n5536), .Y(n9485) );
  NOR2X1 U7351 ( .A(n5763), .B(n5764), .Y(n8609) );
  NOR2X1 U7352 ( .A(n5999), .B(n6000), .Y(n7733) );
  NOR2X1 U7353 ( .A(n4905), .B(n4906), .Y(n11529) );
  NOR2X1 U7354 ( .A(n5213), .B(n5214), .Y(n10653) );
  NOR2X1 U7355 ( .A(n5459), .B(n5460), .Y(n9777) );
  NOR2X1 U7356 ( .A(n5687), .B(n5688), .Y(n8901) );
  NOR2X1 U7357 ( .A(n5923), .B(n5924), .Y(n8025) );
  NOR2XL U7358 ( .A(n31), .B(n3457), .Y(n13862) );
  NOR2XL U7359 ( .A(n34), .B(n3155), .Y(n15437) );
  NOR2XL U7360 ( .A(n35), .B(n2553), .Y(n18587) );
  NOR2XL U7361 ( .A(n30), .B(n2863), .Y(n17012) );
  NOR2XL U7362 ( .A(n36), .B(n2917), .Y(n16697) );
  NOR2XL U7363 ( .A(n32), .B(n2614), .Y(n18272) );
  NOR2XL U7364 ( .A(n33), .B(n3223), .Y(n15122) );
  NOR2XL U7365 ( .A(n37), .B(n3277), .Y(n14807) );
  NOR2XL U7366 ( .A(n38), .B(n2978), .Y(n16382) );
  NOR2XL U7367 ( .A(n39), .B(n2682), .Y(n17957) );
  NOR2XL U7368 ( .A(n40), .B(n3338), .Y(n14492) );
  NOR2XL U7369 ( .A(n41), .B(n3036), .Y(n16067) );
  NOR2XL U7370 ( .A(n42), .B(n2742), .Y(n17642) );
  NOR2XL U7371 ( .A(n43), .B(n3396), .Y(n14177) );
  NOR2XL U7372 ( .A(n44), .B(n3104), .Y(n15752) );
  NOR2XL U7373 ( .A(n45), .B(n2796), .Y(n17327) );
  NAND2X1 U7374 ( .A(n418), .B(n634), .Y(n13892) );
  NAND2X1 U7375 ( .A(n417), .B(n633), .Y(n17042) );
  NAND2X1 U7376 ( .A(n419), .B(n635), .Y(n18302) );
  NAND2X1 U7377 ( .A(n420), .B(n636), .Y(n15152) );
  NAND2X1 U7378 ( .A(n426), .B(n637), .Y(n15467) );
  NAND2X1 U7379 ( .A(n428), .B(n638), .Y(n18617) );
  NAND2X1 U7380 ( .A(n430), .B(n639), .Y(n16727) );
  NAND2X1 U7381 ( .A(n432), .B(n640), .Y(n14837) );
  NAND2X1 U7382 ( .A(n425), .B(n641), .Y(n16412) );
  NAND2X1 U7383 ( .A(n421), .B(n642), .Y(n17987) );
  NAND2X1 U7384 ( .A(n427), .B(n643), .Y(n14522) );
  NAND2X1 U7385 ( .A(n422), .B(n644), .Y(n16097) );
  NAND2X1 U7386 ( .A(n429), .B(n645), .Y(n17672) );
  NAND2X1 U7387 ( .A(n423), .B(n646), .Y(n14207) );
  NAND2X1 U7388 ( .A(n431), .B(n647), .Y(n15782) );
  NAND2X1 U7389 ( .A(n424), .B(n648), .Y(n17357) );
  NOR2X1 U7390 ( .A(n5375), .B(n5371), .Y(n9976) );
  NOR2X1 U7391 ( .A(n6165), .B(n6161), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n162) );
  NOR2X1 U7392 ( .A(n5021), .B(n5017), .Y(n11144) );
  NOR2X1 U7393 ( .A(n5847), .B(n5843), .Y(n8224) );
  NOR2X1 U7394 ( .A(n5105), .B(n5101), .Y(n10852) );
  NOR2X1 U7395 ( .A(n5611), .B(n5607), .Y(n9100) );
  NOR2X1 U7396 ( .A(n6075), .B(n6071), .Y(n7348) );
  NOR2X1 U7397 ( .A(n5291), .B(n5287), .Y(n10268) );
  NOR2X1 U7398 ( .A(n5535), .B(n5531), .Y(n9392) );
  NOR2X1 U7399 ( .A(n5763), .B(n5759), .Y(n8516) );
  NOR2X1 U7400 ( .A(n5999), .B(n5995), .Y(n7640) );
  NOR2X1 U7401 ( .A(n4905), .B(n4901), .Y(n11436) );
  NOR2X1 U7402 ( .A(n5213), .B(n5209), .Y(n10560) );
  NOR2X1 U7403 ( .A(n5459), .B(n5455), .Y(n9684) );
  NOR2X1 U7404 ( .A(n5687), .B(n5683), .Y(n8808) );
  NOR2X1 U7405 ( .A(n5923), .B(n5919), .Y(n7932) );
  CLKINVX3 U7406 ( .A(n3918), .Y(n3836) );
  CLKINVX3 U7407 ( .A(n3918), .Y(n3835) );
  CLKINVX3 U7408 ( .A(n3919), .Y(n3834) );
  CLKINVX3 U7409 ( .A(n3919), .Y(n3833) );
  CLKINVX3 U7410 ( .A(n3920), .Y(n3831) );
  CLKINVX3 U7411 ( .A(n3920), .Y(n3830) );
  CLKINVX3 U7412 ( .A(n3920), .Y(n3829) );
  CLKINVX3 U7413 ( .A(n3921), .Y(n3828) );
  CLKINVX3 U7414 ( .A(n3919), .Y(n3832) );
  CLKINVX3 U7415 ( .A(n3935), .Y(n3847) );
  CLKINVX3 U7416 ( .A(n3931), .Y(n3846) );
  CLKINVX3 U7417 ( .A(n3919), .Y(n3845) );
  CLKINVX3 U7418 ( .A(n3917), .Y(n3844) );
  CLKINVX3 U7419 ( .A(n3921), .Y(n3843) );
  CLKINVX3 U7420 ( .A(n3940), .Y(n3841) );
  CLKINVX3 U7421 ( .A(n3917), .Y(n3840) );
  CLKINVX3 U7422 ( .A(n3917), .Y(n3839) );
  CLKINVX3 U7423 ( .A(n3917), .Y(n3838) );
  CLKINVX3 U7424 ( .A(n3918), .Y(n3837) );
  CLKINVX3 U7425 ( .A(n3939), .Y(n3842) );
  CLKINVX3 U7426 ( .A(n3925), .Y(n3816) );
  CLKINVX3 U7427 ( .A(n3925), .Y(n3815) );
  CLKINVX3 U7428 ( .A(n3925), .Y(n3814) );
  CLKINVX3 U7429 ( .A(n3926), .Y(n3813) );
  CLKINVX3 U7430 ( .A(n3926), .Y(n3812) );
  CLKINVX3 U7431 ( .A(n3927), .Y(n3810) );
  CLKINVX3 U7432 ( .A(n3927), .Y(n3809) );
  CLKINVX3 U7433 ( .A(n3927), .Y(n3808) );
  CLKINVX3 U7434 ( .A(n3928), .Y(n3807) );
  CLKINVX3 U7435 ( .A(n3926), .Y(n3811) );
  CLKINVX3 U7436 ( .A(n3921), .Y(n3826) );
  CLKINVX3 U7437 ( .A(n3922), .Y(n3825) );
  CLKINVX3 U7438 ( .A(n3922), .Y(n3824) );
  CLKINVX3 U7439 ( .A(n3922), .Y(n3823) );
  CLKINVX3 U7440 ( .A(n3923), .Y(n3821) );
  CLKINVX3 U7441 ( .A(n3923), .Y(n3820) );
  CLKINVX3 U7442 ( .A(n3924), .Y(n3819) );
  CLKINVX3 U7443 ( .A(n3924), .Y(n3818) );
  CLKINVX3 U7444 ( .A(n3924), .Y(n3817) );
  CLKINVX3 U7445 ( .A(n3923), .Y(n3822) );
  CLKINVX3 U7446 ( .A(n3921), .Y(n3827) );
  CLKINVX3 U7447 ( .A(n3962), .Y(n3882) );
  CLKINVX3 U7448 ( .A(n3910), .Y(n3881) );
  CLKINVX3 U7449 ( .A(n3908), .Y(n3880) );
  CLKINVX3 U7450 ( .A(n3910), .Y(n3879) );
  CLKINVX3 U7451 ( .A(n3910), .Y(n3878) );
  CLKINVX3 U7452 ( .A(n3910), .Y(n3877) );
  CLKINVX3 U7453 ( .A(n3911), .Y(n3875) );
  CLKINVX3 U7454 ( .A(n3911), .Y(n3874) );
  CLKINVX3 U7455 ( .A(n3912), .Y(n3873) );
  CLKINVX3 U7456 ( .A(n3912), .Y(n3872) );
  CLKINVX3 U7457 ( .A(n3912), .Y(n3871) );
  CLKINVX3 U7458 ( .A(n3911), .Y(n3876) );
  CLKINVX3 U7459 ( .A(n3909), .Y(n3884) );
  CLKINVX3 U7460 ( .A(n3909), .Y(n3885) );
  CLKINVX3 U7461 ( .A(n3908), .Y(n3886) );
  CLKINVX3 U7462 ( .A(n3908), .Y(n3887) );
  CLKINVX3 U7463 ( .A(n3908), .Y(n3888) );
  CLKINVX3 U7464 ( .A(n3909), .Y(n3883) );
  CLKINVX3 U7465 ( .A(n3924), .Y(n3858) );
  CLKINVX3 U7466 ( .A(n3923), .Y(n3857) );
  CLKINVX3 U7467 ( .A(n3936), .Y(n3856) );
  CLKINVX3 U7468 ( .A(n3943), .Y(n3855) );
  CLKINVX3 U7469 ( .A(n3941), .Y(n3854) );
  CLKINVX3 U7470 ( .A(n3915), .Y(n3852) );
  CLKINVX3 U7471 ( .A(n3912), .Y(n3851) );
  CLKINVX3 U7472 ( .A(n3911), .Y(n3850) );
  CLKINVX3 U7473 ( .A(n3930), .Y(n3849) );
  CLKINVX3 U7474 ( .A(n3920), .Y(n3848) );
  CLKINVX3 U7475 ( .A(n3914), .Y(n3853) );
  CLKINVX3 U7476 ( .A(n3913), .Y(n3869) );
  CLKINVX3 U7477 ( .A(n3913), .Y(n3868) );
  CLKINVX3 U7478 ( .A(n3914), .Y(n3867) );
  CLKINVX3 U7479 ( .A(n3914), .Y(n3866) );
  CLKINVX3 U7480 ( .A(n3914), .Y(n3865) );
  CLKINVX3 U7481 ( .A(n3915), .Y(n3863) );
  CLKINVX3 U7482 ( .A(n3915), .Y(n3862) );
  CLKINVX3 U7483 ( .A(n3916), .Y(n3861) );
  CLKINVX3 U7484 ( .A(n3916), .Y(n3860) );
  CLKINVX3 U7485 ( .A(n3916), .Y(n3859) );
  CLKINVX3 U7486 ( .A(n3915), .Y(n3864) );
  CLKINVX3 U7487 ( .A(n3913), .Y(n3870) );
  CLKINVX3 U7488 ( .A(n3943), .Y(n3743) );
  CLKINVX3 U7489 ( .A(n3943), .Y(n3742) );
  CLKINVX3 U7490 ( .A(n3943), .Y(n3741) );
  CLKINVX3 U7491 ( .A(n3941), .Y(n3740) );
  CLKINVX3 U7492 ( .A(n3914), .Y(n3739) );
  CLKINVX3 U7493 ( .A(n3937), .Y(n3737) );
  CLKINVX3 U7494 ( .A(n3935), .Y(n3736) );
  CLKINVX3 U7495 ( .A(n3942), .Y(n3735) );
  CLKINVX3 U7496 ( .A(n3925), .Y(n3734) );
  CLKINVX3 U7497 ( .A(n3924), .Y(n3733) );
  CLKINVX3 U7498 ( .A(n3932), .Y(n3738) );
  CLKINVX3 U7499 ( .A(n3927), .Y(n3756) );
  CLKINVX3 U7500 ( .A(n3926), .Y(n3755) );
  CLKINVX3 U7501 ( .A(n3928), .Y(n3754) );
  CLKINVX3 U7502 ( .A(n3938), .Y(n3753) );
  CLKINVX3 U7503 ( .A(n3940), .Y(n3752) );
  CLKINVX3 U7504 ( .A(n3939), .Y(n3751) );
  CLKINVX3 U7505 ( .A(n3941), .Y(n3749) );
  CLKINVX3 U7506 ( .A(n3941), .Y(n3748) );
  CLKINVX3 U7507 ( .A(n3942), .Y(n3747) );
  CLKINVX3 U7508 ( .A(n3942), .Y(n3746) );
  CLKINVX3 U7509 ( .A(n3942), .Y(n3745) );
  CLKINVX3 U7510 ( .A(n3943), .Y(n3744) );
  CLKINVX3 U7511 ( .A(n3941), .Y(n3750) );
  CLKINVX3 U7512 ( .A(n3945), .Y(n3718) );
  CLKINVX3 U7513 ( .A(n3946), .Y(n3717) );
  CLKINVX3 U7514 ( .A(n3946), .Y(n3716) );
  CLKINVX3 U7515 ( .A(n3946), .Y(n3715) );
  CLKINVX3 U7516 ( .A(n3933), .Y(n3731) );
  CLKINVX3 U7517 ( .A(n3937), .Y(n3730) );
  CLKINVX3 U7518 ( .A(n3934), .Y(n3729) );
  CLKINVX3 U7519 ( .A(n3933), .Y(n3728) );
  CLKINVX3 U7520 ( .A(n3923), .Y(n3727) );
  CLKINVX3 U7521 ( .A(n3915), .Y(n3726) );
  CLKINVX3 U7522 ( .A(n3912), .Y(n3724) );
  CLKINVX3 U7523 ( .A(n3944), .Y(n3723) );
  CLKINVX3 U7524 ( .A(n3944), .Y(n3721) );
  CLKINVX3 U7525 ( .A(n3945), .Y(n3720) );
  CLKINVX3 U7526 ( .A(n3945), .Y(n3719) );
  CLKINVX3 U7527 ( .A(n3911), .Y(n3725) );
  CLKINVX3 U7528 ( .A(n3925), .Y(n3732) );
  CLKINVX3 U7529 ( .A(n3929), .Y(n3793) );
  CLKINVX3 U7530 ( .A(n3909), .Y(n3792) );
  CLKINVX3 U7531 ( .A(n3946), .Y(n3791) );
  CLKINVX3 U7532 ( .A(n3944), .Y(n3790) );
  CLKINVX3 U7533 ( .A(n3922), .Y(n3789) );
  CLKINVX3 U7534 ( .A(n3945), .Y(n3787) );
  CLKINVX3 U7535 ( .A(n3932), .Y(n3786) );
  CLKINVX3 U7536 ( .A(n3932), .Y(n3785) );
  CLKINVX3 U7537 ( .A(n3932), .Y(n3784) );
  CLKINVX3 U7538 ( .A(n3933), .Y(n3783) );
  CLKINVX3 U7539 ( .A(n3933), .Y(n3782) );
  CLKINVX3 U7540 ( .A(n3961), .Y(n3788) );
  CLKINVX3 U7541 ( .A(n3928), .Y(n3805) );
  CLKINVX3 U7542 ( .A(n3929), .Y(n3804) );
  CLKINVX3 U7543 ( .A(n3929), .Y(n3803) );
  CLKINVX3 U7544 ( .A(n3929), .Y(n3802) );
  CLKINVX3 U7545 ( .A(n3930), .Y(n3801) );
  CLKINVX3 U7546 ( .A(n3930), .Y(n3799) );
  CLKINVX3 U7547 ( .A(n3931), .Y(n3798) );
  CLKINVX3 U7548 ( .A(n3931), .Y(n3797) );
  CLKINVX3 U7549 ( .A(n3931), .Y(n3796) );
  CLKINVX3 U7550 ( .A(n3927), .Y(n3795) );
  CLKINVX3 U7551 ( .A(n3926), .Y(n3794) );
  CLKINVX3 U7552 ( .A(n3930), .Y(n3800) );
  CLKINVX3 U7553 ( .A(n3938), .Y(n3768) );
  CLKINVX3 U7554 ( .A(n3938), .Y(n3767) );
  CLKINVX3 U7555 ( .A(n3938), .Y(n3766) );
  CLKINVX3 U7556 ( .A(n3939), .Y(n3765) );
  CLKINVX3 U7557 ( .A(n3939), .Y(n3764) );
  CLKINVX3 U7558 ( .A(n3940), .Y(n3762) );
  CLKINVX3 U7559 ( .A(n3940), .Y(n3761) );
  CLKINVX3 U7560 ( .A(n3940), .Y(n3760) );
  CLKINVX3 U7561 ( .A(n3936), .Y(n3759) );
  CLKINVX3 U7562 ( .A(n3907), .Y(n3758) );
  CLKINVX3 U7563 ( .A(n3916), .Y(n3757) );
  CLKINVX3 U7564 ( .A(n3939), .Y(n3763) );
  CLKINVX3 U7565 ( .A(n3934), .Y(n3780) );
  CLKINVX3 U7566 ( .A(n3934), .Y(n3779) );
  CLKINVX3 U7567 ( .A(n3934), .Y(n3778) );
  CLKINVX3 U7568 ( .A(n3935), .Y(n3777) );
  CLKINVX3 U7569 ( .A(n3935), .Y(n3776) );
  CLKINVX3 U7570 ( .A(n3936), .Y(n3774) );
  CLKINVX3 U7571 ( .A(n3936), .Y(n3773) );
  CLKINVX3 U7572 ( .A(n3936), .Y(n3772) );
  CLKINVX3 U7573 ( .A(n3937), .Y(n3771) );
  CLKINVX3 U7574 ( .A(n3937), .Y(n3770) );
  CLKINVX3 U7575 ( .A(n3937), .Y(n3769) );
  CLKINVX3 U7576 ( .A(n3935), .Y(n3775) );
  CLKINVX3 U7577 ( .A(n3933), .Y(n3781) );
  CLKINVX3 U7578 ( .A(n3928), .Y(n3806) );
  CLKINVX3 U7579 ( .A(n3919), .Y(n3889) );
  CLKINVX3 U7580 ( .A(n3917), .Y(n3890) );
  CLKINVX3 U7581 ( .A(n3947), .Y(n3901) );
  CLKINVX3 U7582 ( .A(n3920), .Y(n3892) );
  CLKINVX3 U7583 ( .A(n3922), .Y(n3894) );
  CLKINVX3 U7584 ( .A(n3944), .Y(n3895) );
  CLKINVX3 U7585 ( .A(n3945), .Y(n3896) );
  CLKINVX3 U7586 ( .A(n3921), .Y(n3893) );
  CLKINVX3 U7587 ( .A(n3918), .Y(n3891) );
  CLKINVX3 U7588 ( .A(n3942), .Y(n3903) );
  CLKINVX3 U7589 ( .A(n3916), .Y(n3902) );
  CLKINVX3 U7590 ( .A(n3909), .Y(n3897) );
  CLKINVX3 U7591 ( .A(n3961), .Y(n3898) );
  CLKINVX3 U7592 ( .A(n3931), .Y(n3899) );
  CLKINVX3 U7593 ( .A(n3946), .Y(n3900) );
  CLKINVX3 U7594 ( .A(n13912), .Y(n6151) );
  CLKINVX3 U7595 ( .A(n17062), .Y(n5380) );
  CLKINVX3 U7596 ( .A(n18322), .Y(n5026) );
  CLKINVX3 U7597 ( .A(n15172), .Y(n5852) );
  CLKINVX3 U7598 ( .A(n15487), .Y(n5768) );
  CLKINVX3 U7599 ( .A(n18637), .Y(n4910) );
  CLKINVX3 U7600 ( .A(n16747), .Y(n5464) );
  CLKINVX3 U7601 ( .A(n14857), .Y(n5928) );
  CLKINVX3 U7602 ( .A(n16432), .Y(n5540) );
  CLKINVX3 U7603 ( .A(n18007), .Y(n5110) );
  CLKINVX3 U7604 ( .A(n14542), .Y(n6004) );
  CLKINVX3 U7605 ( .A(n16117), .Y(n5616) );
  CLKINVX3 U7606 ( .A(n17692), .Y(n5218) );
  CLKINVX3 U7607 ( .A(n14227), .Y(n6080) );
  CLKINVX3 U7608 ( .A(n15802), .Y(n5692) );
  CLKINVX3 U7609 ( .A(n17377), .Y(n5296) );
  CLKINVX3 U7610 ( .A(n9887), .Y(n5350) );
  CLKINVX3 U7611 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n69), .Y(n6146) );
  CLKINVX3 U7612 ( .A(n11055), .Y(n4996) );
  CLKINVX3 U7613 ( .A(n8135), .Y(n5822) );
  CLKINVX3 U7614 ( .A(n10763), .Y(n5080) );
  CLKINVX3 U7615 ( .A(n7259), .Y(n6050) );
  CLKINVX3 U7616 ( .A(n9011), .Y(n5586) );
  CLKINVX3 U7617 ( .A(n10179), .Y(n5266) );
  CLKINVX3 U7618 ( .A(n9303), .Y(n5510) );
  CLKINVX3 U7619 ( .A(n8427), .Y(n5738) );
  CLKINVX3 U7620 ( .A(n7551), .Y(n5974) );
  CLKINVX3 U7621 ( .A(n11347), .Y(n4880) );
  CLKINVX3 U7622 ( .A(n10471), .Y(n5188) );
  CLKINVX3 U7623 ( .A(n9595), .Y(n5434) );
  CLKINVX3 U7624 ( .A(n8719), .Y(n5662) );
  CLKINVX3 U7625 ( .A(n7843), .Y(n5898) );
  CLKINVX3 U7626 ( .A(n3944), .Y(n3722) );
  CLKINVX3 U7627 ( .A(n13293), .Y(n6549) );
  CLKINVX3 U7628 ( .A(n12663), .Y(n6844) );
  CLKINVX3 U7629 ( .A(n12978), .Y(n6890) );
  XOR2X1 U7630 ( .A(top_core_EC_mc_n651), .B(top_core_EC_mc_n601), .Y(
        top_core_EC_mc_n709) );
  XOR2X1 U7631 ( .A(top_core_EC_mc_n443), .B(top_core_EC_mc_n370), .Y(
        top_core_EC_mc_n486) );
  XOR2X1 U7632 ( .A(top_core_EC_mc_n639), .B(top_core_EC_mc_n578), .Y(
        top_core_EC_mc_n695) );
  XOR2X1 U7633 ( .A(top_core_EC_mc_n633), .B(top_core_EC_mc_n571), .Y(
        top_core_EC_mc_n688) );
  XOR2X1 U7634 ( .A(top_core_EC_mc_n621), .B(top_core_EC_mc_n9), .Y(
        top_core_EC_mc_n620) );
  XOR2X1 U7635 ( .A(top_core_EC_mc_n670), .B(top_core_EC_mc_n615), .Y(
        top_core_EC_mc_n849) );
  XOR2X1 U7636 ( .A(top_core_EC_mc_n664), .B(top_core_EC_mc_n608), .Y(
        top_core_EC_mc_n776) );
  XOR2X1 U7637 ( .A(top_core_EC_mc_n627), .B(top_core_EC_mc_n102), .Y(
        top_core_EC_mc_n626) );
  XOR2X1 U7638 ( .A(top_core_EC_mc_n451), .B(top_core_EC_mc_n378), .Y(
        top_core_EC_mc_n491) );
  XOR2X1 U7639 ( .A(top_core_EC_mc_n645), .B(top_core_EC_mc_n594), .Y(
        top_core_EC_mc_n702) );
  OAI22XL U7640 ( .A0(n1144), .A1(n165), .B0(n3506), .B1(n58), .Y(n14120) );
  OAI22XL U7641 ( .A0(n1005), .A1(n164), .B0(n2905), .B1(n57), .Y(n17270) );
  OAI22XL U7642 ( .A0(n949), .A1(n166), .B0(n2663), .B1(n59), .Y(n18530) );
  OAI22XL U7643 ( .A0(n1089), .A1(n167), .B0(n3265), .B1(n60), .Y(n15380) );
  OAI22XL U7644 ( .A0(n1075), .A1(n168), .B0(n3204), .B1(n61), .Y(n15695) );
  OAI22XL U7645 ( .A0(n935), .A1(n169), .B0(n2602), .B1(n63), .Y(n18845) );
  OAI22XL U7646 ( .A0(n1019), .A1(n170), .B0(n2966), .B1(n62), .Y(n16955) );
  OAI22XL U7647 ( .A0(n1103), .A1(n171), .B0(n3323), .B1(n64), .Y(n15065) );
  OAI22XL U7648 ( .A0(n1033), .A1(n172), .B0(n3024), .B1(n65), .Y(n16640) );
  OAI22XL U7649 ( .A0(n963), .A1(n173), .B0(n2723), .B1(n66), .Y(n18215) );
  OAI22XL U7650 ( .A0(n1117), .A1(n174), .B0(n3384), .B1(n67), .Y(n14750) );
  OAI22XL U7651 ( .A0(n1047), .A1(n175), .B0(n3085), .B1(n68), .Y(n16325) );
  OAI22XL U7652 ( .A0(n977), .A1(n176), .B0(n2781), .B1(n69), .Y(n17900) );
  OAI22XL U7653 ( .A0(n1131), .A1(n177), .B0(n3445), .B1(n70), .Y(n14435) );
  OAI22XL U7654 ( .A0(n1061), .A1(n178), .B0(n3143), .B1(n71), .Y(n16010) );
  OAI22XL U7655 ( .A0(n991), .A1(n179), .B0(n2837), .B1(n72), .Y(n17585) );
  NAND2XL U7656 ( .A(n9896), .B(n9887), .Y(n10040) );
  NAND2XL U7657 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n69), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n226) );
  NAND2XL U7658 ( .A(n11064), .B(n11055), .Y(n11208) );
  NAND2XL U7659 ( .A(n8144), .B(n8135), .Y(n8288) );
  NAND2XL U7660 ( .A(n10772), .B(n10763), .Y(n10916) );
  NAND2XL U7661 ( .A(n9020), .B(n9011), .Y(n9164) );
  NAND2XL U7662 ( .A(n7268), .B(n7259), .Y(n7412) );
  NAND2XL U7663 ( .A(n10188), .B(n10179), .Y(n10332) );
  NAND2XL U7664 ( .A(n9312), .B(n9303), .Y(n9456) );
  NAND2XL U7665 ( .A(n8436), .B(n8427), .Y(n8580) );
  NAND2XL U7666 ( .A(n7560), .B(n7551), .Y(n7704) );
  NAND2XL U7667 ( .A(n11356), .B(n11347), .Y(n11500) );
  NAND2XL U7668 ( .A(n10480), .B(n10471), .Y(n10624) );
  NAND2XL U7669 ( .A(n9604), .B(n9595), .Y(n9748) );
  NAND2XL U7670 ( .A(n8728), .B(n8719), .Y(n8872) );
  NAND2XL U7671 ( .A(n7852), .B(n7843), .Y(n7996) );
  NAND2X1 U7672 ( .A(n5363), .B(n5330), .Y(n17033) );
  NAND2X1 U7673 ( .A(n6131), .B(n6114), .Y(n13883) );
  NAND2X1 U7674 ( .A(n5009), .B(n4976), .Y(n18293) );
  NAND2X1 U7675 ( .A(n5835), .B(n5802), .Y(n15143) );
  NAND2X1 U7676 ( .A(n5751), .B(n5718), .Y(n15458) );
  NAND2X1 U7677 ( .A(n4893), .B(n4860), .Y(n18608) );
  NAND2X1 U7678 ( .A(n5447), .B(n5414), .Y(n16718) );
  NAND2X1 U7679 ( .A(n5911), .B(n5878), .Y(n14828) );
  NAND2X1 U7680 ( .A(n5523), .B(n5490), .Y(n16403) );
  NAND2X1 U7681 ( .A(n5093), .B(n5060), .Y(n17978) );
  NAND2X1 U7682 ( .A(n5987), .B(n5954), .Y(n14513) );
  NAND2X1 U7683 ( .A(n5599), .B(n5566), .Y(n16088) );
  NAND2X1 U7684 ( .A(n5201), .B(n5168), .Y(n17663) );
  NAND2X1 U7685 ( .A(n6063), .B(n6030), .Y(n14198) );
  NAND2X1 U7686 ( .A(n5675), .B(n5642), .Y(n15773) );
  NAND2X1 U7687 ( .A(n5279), .B(n5246), .Y(n17348) );
  XOR2X1 U7688 ( .A(top_core_EC_mc_mix_in_4_26_), .B(
        top_core_EC_mc_mix_in_4_10_), .Y(top_core_EC_mc_n614) );
  XOR2X1 U7689 ( .A(top_core_EC_mc_mix_in_8[30]), .B(
        top_core_EC_mc_mix_in_8[14]), .Y(top_core_EC_mc_n593) );
  XOR2X1 U7690 ( .A(top_core_EC_mc_mix_in_4_2_), .B(
        top_core_EC_mc_mix_in_4_18_), .Y(top_core_EC_mc_n584) );
  XOR2X1 U7691 ( .A(top_core_EC_mc_mix_in_4_50_), .B(
        top_core_EC_mc_mix_in_4_34_), .Y(top_core_EC_mc_n423) );
  XOR2X1 U7692 ( .A(top_core_EC_mc_mix_in_8[54]), .B(
        top_core_EC_mc_mix_in_8[38]), .Y(top_core_EC_mc_n399) );
  XOR2X1 U7693 ( .A(top_core_EC_mc_mix_in_8[6]), .B(
        top_core_EC_mc_mix_in_8[22]), .Y(top_core_EC_mc_n343) );
  CLKINVX3 U7694 ( .A(n9943), .Y(n5341) );
  CLKINVX3 U7695 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n128), .Y(n6137) );
  CLKINVX3 U7696 ( .A(n11111), .Y(n4987) );
  CLKINVX3 U7697 ( .A(n8191), .Y(n5813) );
  CLKINVX3 U7698 ( .A(n10819), .Y(n5071) );
  CLKINVX3 U7699 ( .A(n7315), .Y(n6041) );
  CLKINVX3 U7700 ( .A(n9067), .Y(n5577) );
  CLKINVX3 U7701 ( .A(n10235), .Y(n5257) );
  CLKINVX3 U7702 ( .A(n9359), .Y(n5501) );
  CLKINVX3 U7703 ( .A(n8483), .Y(n5729) );
  CLKINVX3 U7704 ( .A(n7607), .Y(n5965) );
  CLKINVX3 U7705 ( .A(n11403), .Y(n4871) );
  CLKINVX3 U7706 ( .A(n10527), .Y(n5179) );
  CLKINVX3 U7707 ( .A(n9651), .Y(n5425) );
  CLKINVX3 U7708 ( .A(n8775), .Y(n5653) );
  CLKINVX3 U7709 ( .A(n7899), .Y(n5889) );
  XOR2X1 U7710 ( .A(top_core_EC_mc_mix_in_4_3_), .B(
        top_core_EC_mc_mix_in_4_19_), .Y(top_core_EC_mc_n497) );
  XOR2X1 U7711 ( .A(top_core_EC_mc_mix_in_8[50]), .B(
        top_core_EC_mc_mix_in_8[34]), .Y(top_core_EC_mc_n440) );
  XOR2X1 U7712 ( .A(top_core_EC_mc_mix_in_4_51_), .B(
        top_core_EC_mc_mix_in_4_35_), .Y(top_core_EC_mc_n415) );
  XOR2X1 U7713 ( .A(top_core_EC_mc_mix_in_8[53]), .B(
        top_core_EC_mc_mix_in_8[37]), .Y(top_core_EC_mc_n407) );
  XOR2X1 U7714 ( .A(top_core_EC_mc_mix_in_4_27_), .B(
        top_core_EC_mc_mix_in_4_11_), .Y(top_core_EC_mc_n607) );
  XOR2X1 U7715 ( .A(top_core_EC_mc_mix_in_8[10]), .B(
        top_core_EC_mc_mix_in_8[26]), .Y(top_core_EC_mc_n7) );
  XOR2X1 U7716 ( .A(top_core_EC_mc_mix_in_8[29]), .B(
        top_core_EC_mc_mix_in_8[13]), .Y(top_core_EC_mc_n600) );
  XOR2X1 U7717 ( .A(top_core_EC_mc_n594), .B(top_core_EC_mc_n346), .Y(
        top_core_EC_mc_n592) );
  XOR2X1 U7718 ( .A(top_core_EC_mc_n578), .B(top_core_EC_mc_n257), .Y(
        top_core_EC_mc_n576) );
  XOR2X1 U7719 ( .A(top_core_EC_mc_n571), .B(top_core_EC_mc_n192), .Y(
        top_core_EC_mc_n569) );
  XOR2X1 U7720 ( .A(top_core_EC_mc_n336), .B(top_core_EC_mc_n337), .Y(
        top_core_EC_mc_n334) );
  XOR2X1 U7721 ( .A(top_core_EC_mc_n369), .B(top_core_EC_mc_n370), .Y(
        top_core_EC_mc_n367) );
  XOR2X1 U7722 ( .A(top_core_EC_mc_n601), .B(top_core_EC_mc_n435), .Y(
        top_core_EC_mc_n599) );
  XOR2X1 U7723 ( .A(top_core_EC_mc_n320), .B(top_core_EC_mc_n321), .Y(
        top_core_EC_mc_n318) );
  XOR2X1 U7724 ( .A(top_core_EC_mc_n312), .B(top_core_EC_mc_n313), .Y(
        top_core_EC_mc_n310) );
  XOR2X1 U7725 ( .A(top_core_EC_mc_n102), .B(top_core_EC_mc_n103), .Y(
        top_core_EC_mc_n99) );
  XOR2X1 U7726 ( .A(top_core_EC_mc_n9), .B(top_core_EC_mc_n10), .Y(
        top_core_EC_mc_n6) );
  XOR2X1 U7727 ( .A(top_core_EC_mc_n615), .B(top_core_EC_mc_n587), .Y(
        top_core_EC_mc_n613) );
  XOR2X1 U7728 ( .A(top_core_EC_mc_n608), .B(top_core_EC_mc_n500), .Y(
        top_core_EC_mc_n606) );
  XOR2X1 U7729 ( .A(top_core_EC_mc_n377), .B(top_core_EC_mc_n378), .Y(
        top_core_EC_mc_n375) );
  XOR2X1 U7730 ( .A(top_core_EC_mc_n361), .B(top_core_EC_mc_n362), .Y(
        top_core_EC_mc_n359) );
  XOR2X1 U7731 ( .A(top_core_EC_mc_n353), .B(top_core_EC_mc_n354), .Y(
        top_core_EC_mc_n351) );
  XOR2X1 U7732 ( .A(top_core_EC_mc_n328), .B(top_core_EC_mc_n329), .Y(
        top_core_EC_mc_n326) );
  XOR2X1 U7733 ( .A(top_core_EC_mc_mix_in_8[2]), .B(
        top_core_EC_mc_mix_in_8[18]), .Y(top_core_EC_mc_n657) );
  XOR2X1 U7734 ( .A(top_core_EC_mc_mix_in_8[5]), .B(
        top_core_EC_mc_mix_in_8[21]), .Y(top_core_EC_mc_n432) );
  NAND2X1 U7735 ( .A(n17057), .B(n2852), .Y(n17230) );
  NAND2X1 U7736 ( .A(n13907), .B(n3453), .Y(n14080) );
  NAND2X1 U7737 ( .A(n15167), .B(n3212), .Y(n15340) );
  NAND2X1 U7738 ( .A(n18317), .B(n2610), .Y(n18490) );
  NAND2X1 U7739 ( .A(n15482), .B(n3151), .Y(n15655) );
  NAND2X1 U7740 ( .A(n16742), .B(n2913), .Y(n16915) );
  NAND2X1 U7741 ( .A(n18632), .B(n2549), .Y(n18805) );
  NAND2X1 U7742 ( .A(n14852), .B(n3273), .Y(n15025) );
  NAND2X1 U7743 ( .A(n16427), .B(n2974), .Y(n16600) );
  NAND2X1 U7744 ( .A(n18002), .B(n2671), .Y(n18175) );
  NAND2X1 U7745 ( .A(n14537), .B(n3334), .Y(n14710) );
  NAND2X1 U7746 ( .A(n16112), .B(n3032), .Y(n16285) );
  NAND2X1 U7747 ( .A(n17687), .B(n2731), .Y(n17860) );
  NAND2X1 U7748 ( .A(n14222), .B(n3392), .Y(n14395) );
  NAND2X1 U7749 ( .A(n15797), .B(n3093), .Y(n15970) );
  NAND2X1 U7750 ( .A(n17372), .B(n2792), .Y(n17545) );
  NAND2X1 U7751 ( .A(n17195), .B(n2881), .Y(n17231) );
  NAND2X1 U7752 ( .A(n14045), .B(n3482), .Y(n14081) );
  NAND2X1 U7753 ( .A(n15305), .B(n3241), .Y(n15341) );
  NAND2X1 U7754 ( .A(n18455), .B(n2639), .Y(n18491) );
  NAND2X1 U7755 ( .A(n15620), .B(n3180), .Y(n15656) );
  NAND2X1 U7756 ( .A(n16880), .B(n2942), .Y(n16916) );
  NAND2X1 U7757 ( .A(n18770), .B(n2578), .Y(n18806) );
  NAND2X1 U7758 ( .A(n14990), .B(n3302), .Y(n15026) );
  NAND2X1 U7759 ( .A(n16565), .B(n3003), .Y(n16601) );
  NAND2X1 U7760 ( .A(n18140), .B(n2700), .Y(n18176) );
  NAND2X1 U7761 ( .A(n14675), .B(n3363), .Y(n14711) );
  NAND2X1 U7762 ( .A(n16250), .B(n3061), .Y(n16286) );
  NAND2X1 U7763 ( .A(n17825), .B(n2760), .Y(n17861) );
  NAND2X1 U7764 ( .A(n14360), .B(n3421), .Y(n14396) );
  NAND2X1 U7765 ( .A(n15935), .B(n3122), .Y(n15971) );
  NAND2X1 U7766 ( .A(n17510), .B(n2821), .Y(n17546) );
  INVX1 U7767 ( .A(n13455), .Y(n6558) );
  INVX1 U7768 ( .A(n12825), .Y(n6853) );
  INVX1 U7769 ( .A(n13140), .Y(n6899) );
  NAND2X1 U7770 ( .A(n6825), .B(n605), .Y(n11685) );
  NAND2X1 U7771 ( .A(n6803), .B(n606), .Y(top_core_KE_sb1_n110) );
  NAND2X1 U7772 ( .A(n6529), .B(n601), .Y(n12316) );
  NAND2X1 U7773 ( .A(n6471), .B(n1174), .Y(n13262) );
  NAND2X1 U7774 ( .A(n6506), .B(n608), .Y(n12001) );
  NAND2X1 U7775 ( .A(n6814), .B(n1220), .Y(n12947) );
  NAND2X1 U7776 ( .A(n6518), .B(n1179), .Y(n13577) );
  NAND2X1 U7777 ( .A(n6774), .B(n1214), .Y(n12632) );
  NAND2X1 U7778 ( .A(n3452), .B(n3450), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n171) );
  NAND2X1 U7779 ( .A(n2851), .B(n2848), .Y(n9985) );
  NAND2X1 U7780 ( .A(n2609), .B(n2606), .Y(n11153) );
  NAND2X1 U7781 ( .A(n3211), .B(n3208), .Y(n8233) );
  NAND2X1 U7782 ( .A(n2670), .B(n2667), .Y(n10861) );
  NAND2X1 U7783 ( .A(n3031), .B(n3028), .Y(n9109) );
  NAND2X1 U7784 ( .A(n3391), .B(n3388), .Y(n7357) );
  NAND2X1 U7785 ( .A(n2791), .B(n2788), .Y(n10277) );
  NAND2X1 U7786 ( .A(n2973), .B(n2970), .Y(n9401) );
  NAND2X1 U7787 ( .A(n3150), .B(n3147), .Y(n8525) );
  NAND2X1 U7788 ( .A(n3333), .B(n3330), .Y(n7649) );
  NAND2X1 U7789 ( .A(n2548), .B(n2545), .Y(n11445) );
  NAND2X1 U7790 ( .A(n2730), .B(n2727), .Y(n10569) );
  NAND2X1 U7791 ( .A(n2912), .B(n2909), .Y(n9693) );
  NAND2X1 U7792 ( .A(n3092), .B(n3089), .Y(n8817) );
  NAND2X1 U7793 ( .A(n3272), .B(n3269), .Y(n7941) );
  XNOR2X1 U7794 ( .A(top_core_EC_mc_mix_in_4_26_), .B(top_core_EC_mc_n8), .Y(
        top_core_EC_mc_n618) );
  XNOR2X1 U7795 ( .A(top_core_EC_mc_mix_in_8[30]), .B(top_core_EC_mc_n433), 
        .Y(top_core_EC_mc_n597) );
  XNOR2X1 U7796 ( .A(top_core_EC_mc_mix_in_2_27_), .B(top_core_EC_mc_n498), 
        .Y(top_core_EC_mc_n604) );
  NAND2XL U7797 ( .A(n30), .B(n17162), .Y(n16998) );
  NAND2XL U7798 ( .A(n31), .B(n14012), .Y(n13848) );
  NAND2XL U7799 ( .A(n32), .B(n18422), .Y(n18258) );
  NAND2XL U7800 ( .A(n33), .B(n15272), .Y(n15108) );
  NAND2XL U7801 ( .A(n34), .B(n15587), .Y(n15423) );
  NAND2XL U7802 ( .A(n36), .B(n16847), .Y(n16683) );
  NAND2XL U7803 ( .A(n35), .B(n18737), .Y(n18573) );
  NAND2XL U7804 ( .A(n37), .B(n14957), .Y(n14793) );
  NAND2XL U7805 ( .A(n38), .B(n16532), .Y(n16368) );
  NAND2XL U7806 ( .A(n39), .B(n18107), .Y(n17943) );
  NAND2XL U7807 ( .A(n40), .B(n14642), .Y(n14478) );
  NAND2XL U7808 ( .A(n41), .B(n16217), .Y(n16053) );
  NAND2XL U7809 ( .A(n42), .B(n17792), .Y(n17628) );
  NAND2XL U7810 ( .A(n43), .B(n14327), .Y(n14163) );
  NAND2XL U7811 ( .A(n44), .B(n15902), .Y(n15738) );
  NAND2XL U7812 ( .A(n45), .B(n17477), .Y(n17313) );
  AOI21X1 U7813 ( .A0(n17029), .A1(n17130), .B0(n17030), .Y(n17137) );
  AOI21X1 U7814 ( .A0(n13879), .A1(n13980), .B0(n13880), .Y(n13987) );
  AOI21X1 U7815 ( .A0(n18289), .A1(n18390), .B0(n18290), .Y(n18397) );
  AOI21X1 U7816 ( .A0(n15139), .A1(n15240), .B0(n15140), .Y(n15247) );
  AOI21X1 U7817 ( .A0(n15454), .A1(n15555), .B0(n15455), .Y(n15562) );
  AOI21X1 U7818 ( .A0(n18604), .A1(n18705), .B0(n18605), .Y(n18712) );
  AOI21X1 U7819 ( .A0(n16714), .A1(n16815), .B0(n16715), .Y(n16822) );
  AOI21X1 U7820 ( .A0(n14824), .A1(n14925), .B0(n14825), .Y(n14932) );
  AOI21X1 U7821 ( .A0(n16399), .A1(n16500), .B0(n16400), .Y(n16507) );
  AOI21X1 U7822 ( .A0(n17974), .A1(n18075), .B0(n17975), .Y(n18082) );
  AOI21X1 U7823 ( .A0(n14509), .A1(n14610), .B0(n14510), .Y(n14617) );
  AOI21X1 U7824 ( .A0(n16084), .A1(n16185), .B0(n16085), .Y(n16192) );
  AOI21X1 U7825 ( .A0(n17659), .A1(n17760), .B0(n17660), .Y(n17767) );
  AOI21X1 U7826 ( .A0(n14194), .A1(n14295), .B0(n14195), .Y(n14302) );
  AOI21X1 U7827 ( .A0(n15769), .A1(n15870), .B0(n15770), .Y(n15877) );
  AOI21X1 U7828 ( .A0(n17344), .A1(n17445), .B0(n17345), .Y(n17452) );
  XNOR2X1 U7829 ( .A(n4058), .B(n2395), .Y(top_core_EC_n1021) );
  OAI21XL U7830 ( .A0(n2880), .A1(n30), .B0(n17025), .Y(n17100) );
  OAI21XL U7831 ( .A0(n3481), .A1(n31), .B0(n13875), .Y(n13950) );
  OAI21XL U7832 ( .A0(n2638), .A1(n32), .B0(n18285), .Y(n18360) );
  OAI21XL U7833 ( .A0(n3240), .A1(n33), .B0(n15135), .Y(n15210) );
  OAI21XL U7834 ( .A0(n3179), .A1(n34), .B0(n15450), .Y(n15525) );
  OAI21XL U7835 ( .A0(n2577), .A1(n35), .B0(n18600), .Y(n18675) );
  OAI21XL U7836 ( .A0(n2941), .A1(n36), .B0(n16710), .Y(n16785) );
  OAI21XL U7837 ( .A0(n3301), .A1(n37), .B0(n14820), .Y(n14895) );
  OAI21XL U7838 ( .A0(n3002), .A1(n38), .B0(n16395), .Y(n16470) );
  OAI21XL U7839 ( .A0(n2699), .A1(n39), .B0(n17970), .Y(n18045) );
  OAI21XL U7840 ( .A0(n3362), .A1(n40), .B0(n14505), .Y(n14580) );
  OAI21XL U7841 ( .A0(n3060), .A1(n41), .B0(n16080), .Y(n16155) );
  OAI21XL U7842 ( .A0(n2759), .A1(n42), .B0(n17655), .Y(n17730) );
  OAI21XL U7843 ( .A0(n3420), .A1(n43), .B0(n14190), .Y(n14265) );
  OAI21XL U7844 ( .A0(n3121), .A1(n44), .B0(n15765), .Y(n15840) );
  OAI21XL U7845 ( .A0(n2820), .A1(n45), .B0(n17340), .Y(n17415) );
  AOI21X1 U7846 ( .A0(n6920), .A1(n689), .B0(n6913), .Y(n11923) );
  AOI21X1 U7847 ( .A0(n6874), .A1(n690), .B0(n6867), .Y(top_core_KE_sb1_n352)
         );
  AOI21X1 U7848 ( .A0(n6556), .A1(n692), .B0(n6548), .Y(n13499) );
  AOI21X1 U7849 ( .A0(n6580), .A1(n693), .B0(n6573), .Y(n12239) );
  AOI21X1 U7850 ( .A0(n6851), .A1(n694), .B0(n6843), .Y(n12869) );
  AOI21X1 U7851 ( .A0(n6604), .A1(n695), .B0(n6596), .Y(n13814) );
  AOI21X1 U7852 ( .A0(n6897), .A1(n696), .B0(n6889), .Y(n13184) );
  AOI21X1 U7853 ( .A0(n17073), .A1(n17062), .B0(n337), .Y(n17188) );
  AOI21X1 U7854 ( .A0(n13923), .A1(n13912), .B0(n338), .Y(n14038) );
  AOI21X1 U7855 ( .A0(n18333), .A1(n18322), .B0(n339), .Y(n18448) );
  AOI21X1 U7856 ( .A0(n15183), .A1(n15172), .B0(n340), .Y(n15298) );
  AOI21X1 U7857 ( .A0(n15498), .A1(n15487), .B0(n341), .Y(n15613) );
  AOI21X1 U7858 ( .A0(n16758), .A1(n16747), .B0(n342), .Y(n16873) );
  AOI21X1 U7859 ( .A0(n18648), .A1(n18637), .B0(n343), .Y(n18763) );
  AOI21X1 U7860 ( .A0(n14868), .A1(n14857), .B0(n344), .Y(n14983) );
  AOI21X1 U7861 ( .A0(n16443), .A1(n16432), .B0(n345), .Y(n16558) );
  AOI21X1 U7862 ( .A0(n18018), .A1(n18007), .B0(n346), .Y(n18133) );
  AOI21X1 U7863 ( .A0(n14553), .A1(n14542), .B0(n347), .Y(n14668) );
  AOI21X1 U7864 ( .A0(n16128), .A1(n16117), .B0(n348), .Y(n16243) );
  AOI21X1 U7865 ( .A0(n17703), .A1(n17692), .B0(n349), .Y(n17818) );
  AOI21X1 U7866 ( .A0(n14238), .A1(n14227), .B0(n350), .Y(n14353) );
  AOI21X1 U7867 ( .A0(n15813), .A1(n15802), .B0(n351), .Y(n15928) );
  AOI21X1 U7868 ( .A0(n17388), .A1(n17377), .B0(n352), .Y(n17503) );
  CLKINVX3 U7869 ( .A(n4022), .Y(n3990) );
  CLKINVX3 U7870 ( .A(n4025), .Y(n4009) );
  CLKINVX3 U7871 ( .A(n4023), .Y(n4001) );
  CLKINVX3 U7872 ( .A(n4024), .Y(n4008) );
  CLKINVX3 U7873 ( .A(n4022), .Y(n3991) );
  CLKINVX3 U7874 ( .A(n4027), .Y(n3999) );
  CLKINVX3 U7875 ( .A(n4023), .Y(n3998) );
  CLKINVX3 U7876 ( .A(n4027), .Y(n4003) );
  CLKINVX3 U7877 ( .A(n4024), .Y(n3994) );
  CLKINVX3 U7878 ( .A(n4023), .Y(n4000) );
  CLKINVX3 U7879 ( .A(n4026), .Y(n4011) );
  CLKINVX3 U7880 ( .A(n4028), .Y(n4006) );
  CLKINVX3 U7881 ( .A(n4024), .Y(n3996) );
  CLKINVX3 U7882 ( .A(n4022), .Y(n3995) );
  CLKINVX3 U7883 ( .A(n4023), .Y(n3997) );
  CLKINVX3 U7884 ( .A(n4026), .Y(n4002) );
  CLKINVX3 U7885 ( .A(n4024), .Y(n4007) );
  CLKINVX3 U7886 ( .A(n4025), .Y(n3993) );
  CLKINVX3 U7887 ( .A(n4021), .Y(n3992) );
  CLKINVX3 U7888 ( .A(n4025), .Y(n4010) );
  CLKINVX3 U7889 ( .A(n4021), .Y(n4005) );
  CLKINVX3 U7890 ( .A(n4022), .Y(n4004) );
  INVX1 U7891 ( .A(n11677), .Y(n6824) );
  INVX1 U7892 ( .A(top_core_KE_sb1_n102), .Y(n6802) );
  INVX1 U7893 ( .A(n12308), .Y(n6528) );
  INVX1 U7894 ( .A(n13254), .Y(n6470) );
  INVX1 U7895 ( .A(n11993), .Y(n6505) );
  INVX1 U7896 ( .A(n12624), .Y(n6773) );
  INVX1 U7897 ( .A(n13569), .Y(n6517) );
  INVX1 U7898 ( .A(n12939), .Y(n6813) );
  CLKINVX3 U7899 ( .A(n4026), .Y(n4012) );
  CLKINVX3 U7900 ( .A(n2395), .Y(n2367) );
  CLKINVX3 U7901 ( .A(n4025), .Y(n4016) );
  CLKINVX3 U7902 ( .A(n4027), .Y(n4015) );
  CLKINVX3 U7903 ( .A(n4023), .Y(n4014) );
  CLKINVX3 U7904 ( .A(n4026), .Y(n4017) );
  CLKINVX3 U7905 ( .A(n4027), .Y(n4013) );
  CLKINVX3 U7906 ( .A(n4027), .Y(n4019) );
  NAND4XL U7907 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n135), .B(n14), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n315), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n316), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n314) );
  NAND4XL U7908 ( .A(n9950), .B(n15), .C(n10129), .D(n10130), .Y(n10128) );
  NAND4XL U7909 ( .A(n11118), .B(n16), .C(n11297), .D(n11298), .Y(n11296) );
  NAND4XL U7910 ( .A(n8198), .B(n17), .C(n8377), .D(n8378), .Y(n8376) );
  NAND4XL U7911 ( .A(n10826), .B(n18), .C(n11005), .D(n11006), .Y(n11004) );
  NAND4XL U7912 ( .A(n9074), .B(n19), .C(n9253), .D(n9254), .Y(n9252) );
  NAND4XL U7913 ( .A(n7322), .B(n20), .C(n7501), .D(n7502), .Y(n7500) );
  NAND4XL U7914 ( .A(n10242), .B(n21), .C(n10421), .D(n10422), .Y(n10420) );
  NAND4XL U7915 ( .A(n9366), .B(n22), .C(n9545), .D(n9546), .Y(n9544) );
  NAND4XL U7916 ( .A(n8490), .B(n23), .C(n8669), .D(n8670), .Y(n8668) );
  NAND4XL U7917 ( .A(n7614), .B(n24), .C(n7793), .D(n7794), .Y(n7792) );
  NAND4XL U7918 ( .A(n11410), .B(n25), .C(n11589), .D(n11590), .Y(n11588) );
  NAND4XL U7919 ( .A(n10534), .B(n26), .C(n10713), .D(n10714), .Y(n10712) );
  NAND4XL U7920 ( .A(n9658), .B(n27), .C(n9837), .D(n9838), .Y(n9836) );
  NAND4XL U7921 ( .A(n8782), .B(n28), .C(n8961), .D(n8962), .Y(n8960) );
  NAND4XL U7922 ( .A(n7906), .B(n29), .C(n8085), .D(n8086), .Y(n8084) );
  CLKINVX3 U7923 ( .A(n4091), .Y(n4035) );
  CLKINVX3 U7924 ( .A(n4021), .Y(n3989) );
  CLKINVX3 U7925 ( .A(n4075), .Y(n4036) );
  CLKINVX3 U7926 ( .A(n4077), .Y(n4038) );
  CLKINVX3 U7927 ( .A(n4034), .Y(n4044) );
  CLKINVX3 U7928 ( .A(n4081), .Y(n4040) );
  CLKINVX3 U7929 ( .A(n4086), .Y(n4042) );
  CLKINVX3 U7930 ( .A(n4084), .Y(n4037) );
  CLKINVX3 U7931 ( .A(n4089), .Y(n4047) );
  CLKINVX3 U7932 ( .A(n4073), .Y(n4046) );
  CLKINVX3 U7933 ( .A(n4080), .Y(n4041) );
  CLKINVX3 U7934 ( .A(n4085), .Y(n4049) );
  CLKINVX3 U7935 ( .A(n4094), .Y(n4048) );
  CLKINVX3 U7936 ( .A(n4076), .Y(n4043) );
  CLKINVX3 U7937 ( .A(n4111), .Y(n4045) );
  CLKINVX3 U7938 ( .A(n4076), .Y(n4039) );
  AOI21X1 U7939 ( .A0(n2854), .A1(n10005), .B0(n10006), .Y(n9978) );
  NAND4BXL U7940 ( .AN(n10004), .B(n10013), .C(n10014), .D(n10015), .Y(n10005)
         );
  AOI31X1 U7941 ( .A0(n10007), .A1(n10008), .A2(n10009), .B0(n2862), .Y(n10006) );
  AOI21X1 U7942 ( .A0(n3455), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n191), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n192), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n164) );
  NAND4BXL U7943 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n190), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n199), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n200), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n201), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n191) );
  AOI31X1 U7944 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n193), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n194), .A2(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n195), .B0(n3462), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n192) );
  AOI21X1 U7945 ( .A0(n2612), .A1(n11173), .B0(n11174), .Y(n11146) );
  NAND4BXL U7946 ( .AN(n11172), .B(n11181), .C(n11182), .D(n11183), .Y(n11173)
         );
  AOI31X1 U7947 ( .A0(n11175), .A1(n11176), .A2(n11177), .B0(n2619), .Y(n11174) );
  AOI21X1 U7948 ( .A0(n3214), .A1(n8253), .B0(n8254), .Y(n8226) );
  NAND4BXL U7949 ( .AN(n8252), .B(n8261), .C(n8262), .D(n8263), .Y(n8253) );
  AOI31X1 U7950 ( .A0(n8255), .A1(n8256), .A2(n8257), .B0(n3222), .Y(n8254) );
  AOI21X1 U7951 ( .A0(n2673), .A1(n10881), .B0(n10882), .Y(n10854) );
  NAND4BXL U7952 ( .AN(n10880), .B(n10889), .C(n10890), .D(n10891), .Y(n10881)
         );
  AOI31X1 U7953 ( .A0(n10883), .A1(n10884), .A2(n10885), .B0(n2681), .Y(n10882) );
  AOI21X1 U7954 ( .A0(n3034), .A1(n9129), .B0(n9130), .Y(n9102) );
  NAND4BXL U7955 ( .AN(n9128), .B(n9137), .C(n9138), .D(n9139), .Y(n9129) );
  AOI31X1 U7956 ( .A0(n9131), .A1(n9132), .A2(n9133), .B0(n3041), .Y(n9130) );
  AOI21X1 U7957 ( .A0(n3394), .A1(n7377), .B0(n7378), .Y(n7350) );
  NAND4BXL U7958 ( .AN(n7376), .B(n7385), .C(n7386), .D(n7387), .Y(n7377) );
  AOI31X1 U7959 ( .A0(n7379), .A1(n7380), .A2(n7381), .B0(n3401), .Y(n7378) );
  AOI21X1 U7960 ( .A0(n2794), .A1(n10297), .B0(n10298), .Y(n10270) );
  NAND4BXL U7961 ( .AN(n10296), .B(n10305), .C(n10306), .D(n10307), .Y(n10297)
         );
  AOI31X1 U7962 ( .A0(n10299), .A1(n10300), .A2(n10301), .B0(n2801), .Y(n10298) );
  AOI21X1 U7963 ( .A0(n2976), .A1(n9421), .B0(n9422), .Y(n9394) );
  NAND4BXL U7964 ( .AN(n9420), .B(n9429), .C(n9430), .D(n9431), .Y(n9421) );
  AOI31X1 U7965 ( .A0(n9423), .A1(n9424), .A2(n9425), .B0(n2983), .Y(n9422) );
  AOI21X1 U7966 ( .A0(n3153), .A1(n8545), .B0(n8546), .Y(n8518) );
  NAND4BXL U7967 ( .AN(n8544), .B(n8553), .C(n8554), .D(n8555), .Y(n8545) );
  AOI31X1 U7968 ( .A0(n8547), .A1(n8548), .A2(n8549), .B0(n3160), .Y(n8546) );
  AOI21X1 U7969 ( .A0(n3336), .A1(n7669), .B0(n7670), .Y(n7642) );
  NAND4BXL U7970 ( .AN(n7668), .B(n7677), .C(n7678), .D(n7679), .Y(n7669) );
  AOI31X1 U7971 ( .A0(n7671), .A1(n7672), .A2(n7673), .B0(n3343), .Y(n7670) );
  AOI21X1 U7972 ( .A0(n2551), .A1(n11465), .B0(n11466), .Y(n11438) );
  NAND4BXL U7973 ( .AN(n11464), .B(n11473), .C(n11474), .D(n11475), .Y(n11465)
         );
  AOI31X1 U7974 ( .A0(n11467), .A1(n11468), .A2(n11469), .B0(n2555), .Y(n11466) );
  AOI21X1 U7975 ( .A0(n2733), .A1(n10589), .B0(n10590), .Y(n10562) );
  NAND4BXL U7976 ( .AN(n10588), .B(n10597), .C(n10598), .D(n10599), .Y(n10589)
         );
  AOI31X1 U7977 ( .A0(n10591), .A1(n10592), .A2(n10593), .B0(n2741), .Y(n10590) );
  AOI21X1 U7978 ( .A0(n2915), .A1(n9713), .B0(n9714), .Y(n9686) );
  NAND4BXL U7979 ( .AN(n9712), .B(n9721), .C(n9722), .D(n9723), .Y(n9713) );
  AOI31X1 U7980 ( .A0(n9715), .A1(n9716), .A2(n9717), .B0(n2922), .Y(n9714) );
  AOI21X1 U7981 ( .A0(n3095), .A1(n8837), .B0(n8838), .Y(n8810) );
  NAND4BXL U7982 ( .AN(n8836), .B(n8845), .C(n8846), .D(n8847), .Y(n8837) );
  AOI31X1 U7983 ( .A0(n8839), .A1(n8840), .A2(n8841), .B0(n3103), .Y(n8838) );
  AOI21X1 U7984 ( .A0(n3275), .A1(n7961), .B0(n7962), .Y(n7934) );
  NAND4BXL U7985 ( .AN(n7960), .B(n7969), .C(n7970), .D(n7971), .Y(n7961) );
  AOI31X1 U7986 ( .A0(n7963), .A1(n7964), .A2(n7965), .B0(n3282), .Y(n7962) );
  NAND4X1 U7987 ( .A(n17240), .B(n17164), .C(n17279), .D(n17280), .Y(n17278)
         );
  AOI21X1 U7988 ( .A0(n5380), .A1(n498), .B0(n5361), .Y(n17279) );
  NAND4X1 U7989 ( .A(n14090), .B(n14014), .C(n14129), .D(n14130), .Y(n14128)
         );
  AOI21X1 U7990 ( .A0(n6151), .A1(n497), .B0(n6129), .Y(n14129) );
  NAND4X1 U7991 ( .A(n15350), .B(n15274), .C(n15389), .D(n15390), .Y(n15388)
         );
  AOI21X1 U7992 ( .A0(n5852), .A1(n500), .B0(n5833), .Y(n15389) );
  NAND4X1 U7993 ( .A(n18500), .B(n18424), .C(n18539), .D(n18540), .Y(n18538)
         );
  AOI21X1 U7994 ( .A0(n5026), .A1(n501), .B0(n5007), .Y(n18539) );
  NAND4X1 U7995 ( .A(n15665), .B(n15589), .C(n15704), .D(n15705), .Y(n15703)
         );
  AOI21X1 U7996 ( .A0(n5768), .A1(n499), .B0(n5749), .Y(n15704) );
  NAND4X1 U7997 ( .A(n16925), .B(n16849), .C(n16964), .D(n16965), .Y(n16963)
         );
  AOI21X1 U7998 ( .A0(n5464), .A1(n503), .B0(n5445), .Y(n16964) );
  NAND4X1 U7999 ( .A(n18815), .B(n18739), .C(n18854), .D(n18855), .Y(n18853)
         );
  AOI21X1 U8000 ( .A0(n4910), .A1(n502), .B0(n4891), .Y(n18854) );
  NAND4X1 U8001 ( .A(n15035), .B(n14959), .C(n15074), .D(n15075), .Y(n15073)
         );
  AOI21X1 U8002 ( .A0(n5928), .A1(n504), .B0(n5909), .Y(n15074) );
  NAND4X1 U8003 ( .A(n16610), .B(n16534), .C(n16649), .D(n16650), .Y(n16648)
         );
  AOI21X1 U8004 ( .A0(n5540), .A1(n505), .B0(n5521), .Y(n16649) );
  NAND4X1 U8005 ( .A(n18185), .B(n18109), .C(n18224), .D(n18225), .Y(n18223)
         );
  AOI21X1 U8006 ( .A0(n5110), .A1(n506), .B0(n5091), .Y(n18224) );
  NAND4X1 U8007 ( .A(n14720), .B(n14644), .C(n14759), .D(n14760), .Y(n14758)
         );
  AOI21X1 U8008 ( .A0(n6004), .A1(n507), .B0(n5985), .Y(n14759) );
  NAND4X1 U8009 ( .A(n16295), .B(n16219), .C(n16334), .D(n16335), .Y(n16333)
         );
  AOI21X1 U8010 ( .A0(n5616), .A1(n508), .B0(n5597), .Y(n16334) );
  NAND4X1 U8011 ( .A(n17870), .B(n17794), .C(n17909), .D(n17910), .Y(n17908)
         );
  AOI21X1 U8012 ( .A0(n5218), .A1(n509), .B0(n5199), .Y(n17909) );
  NAND4X1 U8013 ( .A(n14405), .B(n14329), .C(n14444), .D(n14445), .Y(n14443)
         );
  AOI21X1 U8014 ( .A0(n6080), .A1(n510), .B0(n6061), .Y(n14444) );
  NAND4X1 U8015 ( .A(n15980), .B(n15904), .C(n16019), .D(n16020), .Y(n16018)
         );
  AOI21X1 U8016 ( .A0(n5692), .A1(n511), .B0(n5673), .Y(n16019) );
  NAND4X1 U8017 ( .A(n17555), .B(n17479), .C(n17594), .D(n17595), .Y(n17593)
         );
  AOI21X1 U8018 ( .A0(n5296), .A1(n512), .B0(n5277), .Y(n17594) );
  NAND4BXL U8019 ( .AN(n17218), .B(n17219), .C(n17164), .D(n17143), .Y(n17217)
         );
  NAND4BXL U8020 ( .AN(n14068), .B(n14069), .C(n14014), .D(n13993), .Y(n14067)
         );
  NAND4BXL U8021 ( .AN(n15328), .B(n15329), .C(n15274), .D(n15253), .Y(n15327)
         );
  NAND4BXL U8022 ( .AN(n18478), .B(n18479), .C(n18424), .D(n18403), .Y(n18477)
         );
  NAND4BXL U8023 ( .AN(n15643), .B(n15644), .C(n15589), .D(n15568), .Y(n15642)
         );
  NAND4BXL U8024 ( .AN(n16903), .B(n16904), .C(n16849), .D(n16828), .Y(n16902)
         );
  NAND4BXL U8025 ( .AN(n18793), .B(n18794), .C(n18739), .D(n18718), .Y(n18792)
         );
  NAND4BXL U8026 ( .AN(n15013), .B(n15014), .C(n14959), .D(n14938), .Y(n15012)
         );
  NAND4BXL U8027 ( .AN(n16588), .B(n16589), .C(n16534), .D(n16513), .Y(n16587)
         );
  NAND4BXL U8028 ( .AN(n18163), .B(n18164), .C(n18109), .D(n18088), .Y(n18162)
         );
  NAND4BXL U8029 ( .AN(n14698), .B(n14699), .C(n14644), .D(n14623), .Y(n14697)
         );
  NAND4BXL U8030 ( .AN(n16273), .B(n16274), .C(n16219), .D(n16198), .Y(n16272)
         );
  NAND4BXL U8031 ( .AN(n17848), .B(n17849), .C(n17794), .D(n17773), .Y(n17847)
         );
  NAND4BXL U8032 ( .AN(n14383), .B(n14384), .C(n14329), .D(n14308), .Y(n14382)
         );
  NAND4BXL U8033 ( .AN(n15958), .B(n15959), .C(n15904), .D(n15883), .Y(n15957)
         );
  NAND4BXL U8034 ( .AN(n17533), .B(n17534), .C(n17479), .D(n17458), .Y(n17532)
         );
  CLKINVX3 U8035 ( .A(n1876), .Y(n1860) );
  CLKINVX3 U8036 ( .A(n1876), .Y(n1857) );
  CLKINVX3 U8037 ( .A(n1873), .Y(n1858) );
  CLKINVX3 U8038 ( .A(n1876), .Y(n1859) );
  CLKINVX3 U8039 ( .A(n1873), .Y(n1861) );
  CLKINVX3 U8040 ( .A(n1875), .Y(n1865) );
  CLKINVX3 U8041 ( .A(n1875), .Y(n1864) );
  CLKINVX3 U8042 ( .A(n1876), .Y(n1863) );
  CLKINVX3 U8043 ( .A(n1875), .Y(n1862) );
  CLKINVX3 U8044 ( .A(n1854), .Y(n1845) );
  CLKINVX3 U8045 ( .A(n2869), .Y(n2866) );
  CLKINVX3 U8046 ( .A(n2627), .Y(n2624) );
  CLKINVX3 U8047 ( .A(n3229), .Y(n3226) );
  CLKINVX3 U8048 ( .A(n3168), .Y(n3165) );
  CLKINVX3 U8049 ( .A(n3469), .Y(n3467) );
  CLKINVX3 U8050 ( .A(n2566), .Y(n2563) );
  CLKINVX3 U8051 ( .A(n2930), .Y(n2927) );
  CLKINVX3 U8052 ( .A(n3290), .Y(n3287) );
  CLKINVX3 U8053 ( .A(n2991), .Y(n2988) );
  CLKINVX3 U8054 ( .A(n2688), .Y(n2685) );
  CLKINVX3 U8055 ( .A(n3351), .Y(n3348) );
  CLKINVX3 U8056 ( .A(n3049), .Y(n3046) );
  CLKINVX3 U8057 ( .A(n2749), .Y(n2745) );
  CLKINVX3 U8058 ( .A(n3409), .Y(n3406) );
  CLKINVX3 U8059 ( .A(n3110), .Y(n3107) );
  CLKINVX3 U8060 ( .A(n2809), .Y(n2806) );
  CLKINVX3 U8061 ( .A(n1875), .Y(n1866) );
  CLKINVX3 U8062 ( .A(n1914), .Y(n1908) );
  CLKINVX3 U8063 ( .A(n1954), .Y(n1948) );
  CLKINVX3 U8064 ( .A(n1994), .Y(n1988) );
  CLKINVX3 U8065 ( .A(n2074), .Y(n2068) );
  CLKINVX3 U8066 ( .A(n2114), .Y(n2108) );
  CLKINVX3 U8067 ( .A(n1915), .Y(n1905) );
  CLKINVX3 U8068 ( .A(n1955), .Y(n1945) );
  CLKINVX3 U8069 ( .A(n1995), .Y(n1985) );
  CLKINVX3 U8070 ( .A(n2075), .Y(n2065) );
  CLKINVX3 U8071 ( .A(n2115), .Y(n2105) );
  CLKINVX3 U8072 ( .A(n1914), .Y(n1906) );
  CLKINVX3 U8073 ( .A(n1954), .Y(n1946) );
  CLKINVX3 U8074 ( .A(n1994), .Y(n1986) );
  CLKINVX3 U8075 ( .A(n2074), .Y(n2066) );
  CLKINVX3 U8076 ( .A(n2114), .Y(n2106) );
  CLKINVX3 U8077 ( .A(n1914), .Y(n1909) );
  CLKINVX3 U8078 ( .A(n1954), .Y(n1949) );
  CLKINVX3 U8079 ( .A(n1994), .Y(n1989) );
  CLKINVX3 U8080 ( .A(n2074), .Y(n2069) );
  CLKINVX3 U8081 ( .A(n2114), .Y(n2109) );
  CLKINVX3 U8082 ( .A(n1913), .Y(n1910) );
  CLKINVX3 U8083 ( .A(n1953), .Y(n1950) );
  CLKINVX3 U8084 ( .A(n1993), .Y(n1990) );
  CLKINVX3 U8085 ( .A(n2073), .Y(n2070) );
  CLKINVX3 U8086 ( .A(n2113), .Y(n2110) );
  CLKINVX3 U8087 ( .A(n1854), .Y(n1852) );
  CLKINVX3 U8088 ( .A(n1875), .Y(n1872) );
  CLKINVX3 U8089 ( .A(n1853), .Y(n1851) );
  CLKINVX3 U8090 ( .A(n1874), .Y(n1871) );
  CLKINVX3 U8091 ( .A(n1913), .Y(n1911) );
  CLKINVX3 U8092 ( .A(n1953), .Y(n1951) );
  CLKINVX3 U8093 ( .A(n1993), .Y(n1991) );
  CLKINVX3 U8094 ( .A(n2073), .Y(n2071) );
  CLKINVX3 U8095 ( .A(n2113), .Y(n2111) );
  CLKINVX3 U8096 ( .A(n1856), .Y(n1850) );
  CLKINVX3 U8097 ( .A(n1874), .Y(n1870) );
  CLKINVX3 U8098 ( .A(n1853), .Y(n1846) );
  CLKINVX3 U8099 ( .A(n1874), .Y(n1868) );
  CLKINVX3 U8100 ( .A(n1874), .Y(n1869) );
  CLKINVX3 U8101 ( .A(n1856), .Y(n1847) );
  CLKINVX3 U8102 ( .A(n1914), .Y(n1912) );
  CLKINVX3 U8103 ( .A(n1954), .Y(n1952) );
  CLKINVX3 U8104 ( .A(n1994), .Y(n1992) );
  CLKINVX3 U8105 ( .A(n2074), .Y(n2072) );
  CLKINVX3 U8106 ( .A(n2114), .Y(n2112) );
  CLKINVX3 U8107 ( .A(n1855), .Y(n1848) );
  CLKINVX3 U8108 ( .A(n1876), .Y(n1867) );
  CLKINVX3 U8109 ( .A(n1855), .Y(n1849) );
  CLKINVX3 U8110 ( .A(n1914), .Y(n1907) );
  CLKINVX3 U8111 ( .A(n1954), .Y(n1947) );
  CLKINVX3 U8112 ( .A(n1994), .Y(n1987) );
  CLKINVX3 U8113 ( .A(n2074), .Y(n2067) );
  CLKINVX3 U8114 ( .A(n2114), .Y(n2107) );
  CLKINVX3 U8115 ( .A(n2035), .Y(n2025) );
  CLKINVX3 U8116 ( .A(n2034), .Y(n2026) );
  CLKINVX3 U8117 ( .A(n2034), .Y(n2028) );
  CLKINVX3 U8118 ( .A(n2034), .Y(n2029) );
  CLKINVX3 U8119 ( .A(n2033), .Y(n2030) );
  CLKINVX3 U8120 ( .A(n2033), .Y(n2031) );
  CLKINVX3 U8121 ( .A(n2034), .Y(n2032) );
  CLKINVX3 U8122 ( .A(n2034), .Y(n2027) );
  CLKINVX3 U8123 ( .A(n2326), .Y(n2321) );
  CLKINVX3 U8124 ( .A(n2326), .Y(n2324) );
  CLKINVX3 U8125 ( .A(n2325), .Y(n2323) );
  CLKINVX3 U8126 ( .A(n2325), .Y(n2322) );
  CLKINVX3 U8127 ( .A(n738), .Y(n2137) );
  CLKINVX3 U8128 ( .A(n738), .Y(n2138) );
  CLKINVX3 U8129 ( .A(n738), .Y(n2139) );
  CLKINVX3 U8130 ( .A(n738), .Y(n2140) );
  CLKINVX3 U8131 ( .A(n738), .Y(n2141) );
  CLKINVX3 U8132 ( .A(n738), .Y(n2142) );
  CLKINVX3 U8133 ( .A(n738), .Y(n2143) );
  CLKINVX3 U8134 ( .A(n738), .Y(n2144) );
  CLKINVX3 U8135 ( .A(n1913), .Y(n1904) );
  CLKINVX3 U8136 ( .A(n1953), .Y(n1944) );
  CLKINVX3 U8137 ( .A(n1993), .Y(n1984) );
  CLKINVX3 U8138 ( .A(n2073), .Y(n2064) );
  CLKINVX3 U8139 ( .A(n2113), .Y(n2104) );
  CLKINVX3 U8140 ( .A(n2033), .Y(n2024) );
  CLKINVX3 U8141 ( .A(n1854), .Y(n1840) );
  CLKINVX3 U8142 ( .A(n1856), .Y(n1837) );
  CLKINVX3 U8143 ( .A(n1855), .Y(n1838) );
  CLKINVX3 U8144 ( .A(n1855), .Y(n1839) );
  CLKINVX3 U8145 ( .A(n1854), .Y(n1841) );
  CLKINVX3 U8146 ( .A(n1853), .Y(n1842) );
  CLKINVX3 U8147 ( .A(n1854), .Y(n1844) );
  CLKINVX3 U8148 ( .A(n1853), .Y(n1843) );
  CLKINVX3 U8149 ( .A(n9944), .Y(n5366) );
  CLKINVX3 U8150 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n129), .Y(n6156) );
  CLKINVX3 U8151 ( .A(n11112), .Y(n5012) );
  CLKINVX3 U8152 ( .A(n8192), .Y(n5838) );
  CLKINVX3 U8153 ( .A(n10820), .Y(n5096) );
  CLKINVX3 U8154 ( .A(n9068), .Y(n5602) );
  CLKINVX3 U8155 ( .A(n7316), .Y(n6066) );
  CLKINVX3 U8156 ( .A(n10236), .Y(n5282) );
  CLKINVX3 U8157 ( .A(n9360), .Y(n5526) );
  CLKINVX3 U8158 ( .A(n8484), .Y(n5754) );
  CLKINVX3 U8159 ( .A(n7608), .Y(n5990) );
  CLKINVX3 U8160 ( .A(n11404), .Y(n4896) );
  CLKINVX3 U8161 ( .A(n10528), .Y(n5204) );
  CLKINVX3 U8162 ( .A(n9652), .Y(n5450) );
  CLKINVX3 U8163 ( .A(n8776), .Y(n5678) );
  CLKINVX3 U8164 ( .A(n7900), .Y(n5914) );
  CLKINVX3 U8165 ( .A(n14058), .Y(n6121) );
  CLKINVX3 U8166 ( .A(n17208), .Y(n5353) );
  CLKINVX3 U8167 ( .A(n18468), .Y(n4999) );
  CLKINVX3 U8168 ( .A(n15318), .Y(n5825) );
  CLKINVX3 U8169 ( .A(n15633), .Y(n5741) );
  CLKINVX3 U8170 ( .A(n16893), .Y(n5437) );
  CLKINVX3 U8171 ( .A(n18783), .Y(n4883) );
  CLKINVX3 U8172 ( .A(n15003), .Y(n5901) );
  CLKINVX3 U8173 ( .A(n16578), .Y(n5513) );
  CLKINVX3 U8174 ( .A(n18153), .Y(n5083) );
  CLKINVX3 U8175 ( .A(n14688), .Y(n5977) );
  CLKINVX3 U8176 ( .A(n16263), .Y(n5589) );
  CLKINVX3 U8177 ( .A(n17838), .Y(n5191) );
  CLKINVX3 U8178 ( .A(n14373), .Y(n6053) );
  CLKINVX3 U8179 ( .A(n15948), .Y(n5665) );
  CLKINVX3 U8180 ( .A(n17523), .Y(n5269) );
  CLKINVX3 U8181 ( .A(n3675), .Y(n3645) );
  CLKINVX3 U8182 ( .A(n3675), .Y(n3646) );
  CLKINVX3 U8183 ( .A(n3676), .Y(n3647) );
  CLKINVX3 U8184 ( .A(n3676), .Y(n3648) );
  CLKINVX3 U8185 ( .A(n3677), .Y(n3649) );
  CLKINVX3 U8186 ( .A(n3678), .Y(n3650) );
  CLKINVX3 U8187 ( .A(n1916), .Y(n1898) );
  CLKINVX3 U8188 ( .A(n1996), .Y(n1977) );
  CLKINVX3 U8189 ( .A(n2076), .Y(n2057) );
  CLKINVX3 U8190 ( .A(n2116), .Y(n2097) );
  CLKINVX3 U8191 ( .A(n1916), .Y(n1897) );
  CLKINVX3 U8192 ( .A(n1956), .Y(n1937) );
  CLKINVX3 U8193 ( .A(n1956), .Y(n1938) );
  CLKINVX3 U8194 ( .A(n1996), .Y(n1978) );
  CLKINVX3 U8195 ( .A(n2076), .Y(n2058) );
  CLKINVX3 U8196 ( .A(n2116), .Y(n2098) );
  CLKINVX3 U8197 ( .A(n1916), .Y(n1899) );
  CLKINVX3 U8198 ( .A(n1956), .Y(n1939) );
  CLKINVX3 U8199 ( .A(n1996), .Y(n1979) );
  CLKINVX3 U8200 ( .A(n2076), .Y(n2059) );
  CLKINVX3 U8201 ( .A(n2116), .Y(n2099) );
  CLKINVX3 U8202 ( .A(n1916), .Y(n1900) );
  CLKINVX3 U8203 ( .A(n1956), .Y(n1940) );
  CLKINVX3 U8204 ( .A(n1996), .Y(n1980) );
  CLKINVX3 U8205 ( .A(n2076), .Y(n2060) );
  CLKINVX3 U8206 ( .A(n2116), .Y(n2100) );
  CLKINVX3 U8207 ( .A(n1915), .Y(n1901) );
  CLKINVX3 U8208 ( .A(n1955), .Y(n1941) );
  CLKINVX3 U8209 ( .A(n1995), .Y(n1981) );
  CLKINVX3 U8210 ( .A(n2075), .Y(n2061) );
  CLKINVX3 U8211 ( .A(n2115), .Y(n2101) );
  CLKINVX3 U8212 ( .A(n1915), .Y(n1902) );
  CLKINVX3 U8213 ( .A(n1955), .Y(n1942) );
  CLKINVX3 U8214 ( .A(n1995), .Y(n1982) );
  CLKINVX3 U8215 ( .A(n2075), .Y(n2062) );
  CLKINVX3 U8216 ( .A(n2115), .Y(n2102) );
  CLKINVX3 U8217 ( .A(n1915), .Y(n1903) );
  CLKINVX3 U8218 ( .A(n1955), .Y(n1943) );
  CLKINVX3 U8219 ( .A(n1995), .Y(n1983) );
  CLKINVX3 U8220 ( .A(n2075), .Y(n2063) );
  CLKINVX3 U8221 ( .A(n2115), .Y(n2103) );
  CLKINVX3 U8222 ( .A(n2036), .Y(n2017) );
  CLKINVX3 U8223 ( .A(n2036), .Y(n2018) );
  CLKINVX3 U8224 ( .A(n2036), .Y(n2019) );
  CLKINVX3 U8225 ( .A(n2036), .Y(n2020) );
  CLKINVX3 U8226 ( .A(n2035), .Y(n2021) );
  CLKINVX3 U8227 ( .A(n2035), .Y(n2022) );
  CLKINVX3 U8228 ( .A(n2035), .Y(n2023) );
  CLKINVX3 U8229 ( .A(n2316), .Y(n2314) );
  CLKINVX3 U8230 ( .A(n741), .Y(n2315) );
  AND2X2 U8231 ( .A(n6144), .B(n3473), .Y(n545) );
  AND2X2 U8232 ( .A(n5348), .B(n2872), .Y(n546) );
  AND2X2 U8233 ( .A(n4994), .B(n2630), .Y(n547) );
  AND2X2 U8234 ( .A(n5820), .B(n3232), .Y(n548) );
  AND2X2 U8235 ( .A(n5078), .B(n2691), .Y(n549) );
  AND2X2 U8236 ( .A(n5584), .B(n3052), .Y(n550) );
  AND2X2 U8237 ( .A(n6048), .B(n3412), .Y(n551) );
  AND2X2 U8238 ( .A(n5264), .B(n2812), .Y(n552) );
  AND2X2 U8239 ( .A(n5508), .B(n2994), .Y(n553) );
  AND2X2 U8240 ( .A(n5736), .B(n3171), .Y(n554) );
  AND2X2 U8241 ( .A(n5972), .B(n3354), .Y(n555) );
  AND2X2 U8242 ( .A(n4878), .B(n2569), .Y(n556) );
  AND2X2 U8243 ( .A(n5186), .B(n2751), .Y(n557) );
  AND2X2 U8244 ( .A(n5432), .B(n2933), .Y(n558) );
  AND2X2 U8245 ( .A(n5660), .B(n3113), .Y(n559) );
  AND2X2 U8246 ( .A(n5896), .B(n3293), .Y(n560) );
  CLKINVX3 U8247 ( .A(n742), .Y(n3563) );
  CLKINVX3 U8248 ( .A(n742), .Y(n3562) );
  CLKINVX3 U8249 ( .A(n742), .Y(n3561) );
  CLKINVX3 U8250 ( .A(n3543), .Y(n3540) );
  CLKINVX3 U8251 ( .A(n3542), .Y(n3539) );
  CLKINVX3 U8252 ( .A(n3542), .Y(n3538) );
  CLKINVX3 U8253 ( .A(n3542), .Y(n3537) );
  CLKINVX3 U8254 ( .A(n3543), .Y(n3536) );
  CLKINVX3 U8255 ( .A(n3543), .Y(n3535) );
  CLKINVX3 U8256 ( .A(n2326), .Y(n2320) );
  CLKINVX3 U8257 ( .A(n2325), .Y(n2319) );
  CLKINVX3 U8258 ( .A(n2326), .Y(n2318) );
  INVX1 U8259 ( .A(n14089), .Y(n6117) );
  INVX1 U8260 ( .A(n17239), .Y(n5334) );
  INVX1 U8261 ( .A(n18499), .Y(n4980) );
  INVX1 U8262 ( .A(n15349), .Y(n5806) );
  INVX1 U8263 ( .A(n15664), .Y(n5722) );
  INVX1 U8264 ( .A(n18814), .Y(n4864) );
  INVX1 U8265 ( .A(n16924), .Y(n5418) );
  INVX1 U8266 ( .A(n15034), .Y(n5882) );
  INVX1 U8267 ( .A(n16609), .Y(n5494) );
  INVX1 U8268 ( .A(n18184), .Y(n5064) );
  INVX1 U8269 ( .A(n14719), .Y(n5958) );
  INVX1 U8270 ( .A(n16294), .Y(n5570) );
  INVX1 U8271 ( .A(n17869), .Y(n5172) );
  INVX1 U8272 ( .A(n14404), .Y(n6034) );
  INVX1 U8273 ( .A(n15979), .Y(n5646) );
  INVX1 U8274 ( .A(n17554), .Y(n5250) );
  NAND3X1 U8275 ( .A(n1144), .B(n3476), .C(n649), .Y(n13845) );
  NAND3X1 U8276 ( .A(n1005), .B(n2878), .C(n650), .Y(n16995) );
  NAND3X1 U8277 ( .A(n949), .B(n2636), .C(n651), .Y(n18255) );
  NAND3X1 U8278 ( .A(n1089), .B(n3236), .C(n652), .Y(n15105) );
  NAND3X1 U8279 ( .A(n1075), .B(n3175), .C(n653), .Y(n15420) );
  NAND3X1 U8280 ( .A(n935), .B(n2575), .C(n654), .Y(n18570) );
  NAND3X1 U8281 ( .A(n1019), .B(n2939), .C(n655), .Y(n16680) );
  NAND3X1 U8282 ( .A(n1103), .B(n3299), .C(n656), .Y(n14790) );
  NAND3X1 U8283 ( .A(n1033), .B(n3000), .C(n657), .Y(n16365) );
  NAND3X1 U8284 ( .A(n963), .B(n2697), .C(n658), .Y(n17940) );
  NAND3X1 U8285 ( .A(n1117), .B(n3358), .C(n659), .Y(n14475) );
  NAND3X1 U8286 ( .A(n1047), .B(n3058), .C(n660), .Y(n16050) );
  NAND3X1 U8287 ( .A(n977), .B(n2755), .C(n661), .Y(n17625) );
  NAND3X1 U8288 ( .A(n1131), .B(n3418), .C(n662), .Y(n14160) );
  NAND3X1 U8289 ( .A(n1061), .B(n3119), .C(n663), .Y(n15735) );
  NAND3X1 U8290 ( .A(n991), .B(n2818), .C(n664), .Y(n17310) );
  BUFX3 U8291 ( .A(n6123), .Y(n1133) );
  INVXL U8292 ( .A(n31), .Y(n6123) );
  BUFX3 U8293 ( .A(n5355), .Y(n994) );
  INVXL U8294 ( .A(n30), .Y(n5355) );
  BUFX3 U8295 ( .A(n5001), .Y(n938) );
  INVXL U8296 ( .A(n32), .Y(n5001) );
  BUFX3 U8297 ( .A(n5827), .Y(n1078) );
  INVXL U8298 ( .A(n33), .Y(n5827) );
  BUFX3 U8299 ( .A(n5743), .Y(n1064) );
  INVXL U8300 ( .A(n34), .Y(n5743) );
  BUFX3 U8301 ( .A(n5439), .Y(n1008) );
  INVXL U8302 ( .A(n36), .Y(n5439) );
  BUFX3 U8303 ( .A(n4885), .Y(n924) );
  INVXL U8304 ( .A(n35), .Y(n4885) );
  BUFX3 U8305 ( .A(n5903), .Y(n1092) );
  INVXL U8306 ( .A(n37), .Y(n5903) );
  BUFX3 U8307 ( .A(n5515), .Y(n1022) );
  INVXL U8308 ( .A(n38), .Y(n5515) );
  BUFX3 U8309 ( .A(n5085), .Y(n952) );
  INVXL U8310 ( .A(n39), .Y(n5085) );
  BUFX3 U8311 ( .A(n5979), .Y(n1106) );
  INVXL U8312 ( .A(n40), .Y(n5979) );
  BUFX3 U8313 ( .A(n5591), .Y(n1036) );
  INVXL U8314 ( .A(n41), .Y(n5591) );
  BUFX3 U8315 ( .A(n5193), .Y(n966) );
  INVXL U8316 ( .A(n42), .Y(n5193) );
  BUFX3 U8317 ( .A(n6055), .Y(n1120) );
  INVXL U8318 ( .A(n43), .Y(n6055) );
  BUFX3 U8319 ( .A(n5667), .Y(n1050) );
  INVXL U8320 ( .A(n44), .Y(n5667) );
  BUFX3 U8321 ( .A(n5271), .Y(n980) );
  INVXL U8322 ( .A(n45), .Y(n5271) );
  CLKINVX3 U8323 ( .A(n2200), .Y(n2191) );
  CLKINVX3 U8324 ( .A(n2196), .Y(n2192) );
  CLKINVX3 U8325 ( .A(n2203), .Y(n2193) );
  CLKINVX3 U8326 ( .A(n2197), .Y(n2194) );
  CLKINVX3 U8327 ( .A(n2199), .Y(n2195) );
  CLKINVX3 U8328 ( .A(n2202), .Y(n2190) );
  CLKINVX3 U8329 ( .A(n740), .Y(n2154) );
  CLKINVX3 U8330 ( .A(n2211), .Y(n2210) );
  CLKINVX3 U8331 ( .A(n740), .Y(n2155) );
  CLKINVX3 U8332 ( .A(n740), .Y(n2156) );
  CLKINVX3 U8333 ( .A(n2211), .Y(n2209) );
  CLKINVX3 U8334 ( .A(n740), .Y(n2157) );
  CLKINVX3 U8335 ( .A(n2215), .Y(n2208) );
  CLKINVX3 U8336 ( .A(n740), .Y(n2158) );
  CLKINVX3 U8337 ( .A(n2211), .Y(n2207) );
  CLKINVX3 U8338 ( .A(n740), .Y(n2159) );
  CLKINVX3 U8339 ( .A(n2219), .Y(n2206) );
  CLKINVX3 U8340 ( .A(n740), .Y(n2160) );
  CLKINVX3 U8341 ( .A(n2218), .Y(n2205) );
  CLKINVX3 U8342 ( .A(n2284), .Y(n2290) );
  CLKINVX3 U8343 ( .A(n2284), .Y(n2288) );
  CLKINVX3 U8344 ( .A(n2292), .Y(n2287) );
  BUFX3 U8345 ( .A(n6152), .Y(n1137) );
  INVXL U8346 ( .A(n165), .Y(n6152) );
  BUFX3 U8347 ( .A(n5381), .Y(n998) );
  INVXL U8348 ( .A(n164), .Y(n5381) );
  BUFX3 U8349 ( .A(n5027), .Y(n942) );
  INVXL U8350 ( .A(n166), .Y(n5027) );
  BUFX3 U8351 ( .A(n5853), .Y(n1082) );
  INVXL U8352 ( .A(n167), .Y(n5853) );
  BUFX3 U8353 ( .A(n5769), .Y(n1068) );
  INVXL U8354 ( .A(n168), .Y(n5769) );
  BUFX3 U8355 ( .A(n5465), .Y(n1012) );
  INVXL U8356 ( .A(n170), .Y(n5465) );
  BUFX3 U8357 ( .A(n4911), .Y(n928) );
  INVXL U8358 ( .A(n169), .Y(n4911) );
  BUFX3 U8359 ( .A(n5929), .Y(n1096) );
  INVXL U8360 ( .A(n171), .Y(n5929) );
  BUFX3 U8361 ( .A(n5541), .Y(n1026) );
  INVXL U8362 ( .A(n172), .Y(n5541) );
  BUFX3 U8363 ( .A(n5111), .Y(n956) );
  INVXL U8364 ( .A(n173), .Y(n5111) );
  BUFX3 U8365 ( .A(n6005), .Y(n1110) );
  INVXL U8366 ( .A(n174), .Y(n6005) );
  BUFX3 U8367 ( .A(n5617), .Y(n1040) );
  INVXL U8368 ( .A(n175), .Y(n5617) );
  BUFX3 U8369 ( .A(n5219), .Y(n970) );
  INVXL U8370 ( .A(n176), .Y(n5219) );
  BUFX3 U8371 ( .A(n6081), .Y(n1124) );
  INVXL U8372 ( .A(n177), .Y(n6081) );
  BUFX3 U8373 ( .A(n5693), .Y(n1054) );
  INVXL U8374 ( .A(n178), .Y(n5693) );
  BUFX3 U8375 ( .A(n5297), .Y(n984) );
  INVXL U8376 ( .A(n179), .Y(n5297) );
  CLKINVX3 U8377 ( .A(n739), .Y(n2179) );
  CLKINVX3 U8378 ( .A(n739), .Y(n2178) );
  CLKINVX3 U8379 ( .A(n739), .Y(n2177) );
  CLKINVX3 U8380 ( .A(n739), .Y(n2176) );
  CLKINVX3 U8381 ( .A(n739), .Y(n2175) );
  CLKINVX3 U8382 ( .A(n739), .Y(n2174) );
  CLKINVX3 U8383 ( .A(n739), .Y(n2173) );
  CLKINVX3 U8384 ( .A(n3543), .Y(n3541) );
  CLKINVX3 U8385 ( .A(n2869), .Y(n2867) );
  CLKINVX3 U8386 ( .A(n3469), .Y(n3468) );
  CLKINVX3 U8387 ( .A(n2627), .Y(n2625) );
  CLKINVX3 U8388 ( .A(n3229), .Y(n3227) );
  CLKINVX3 U8389 ( .A(n3168), .Y(n3166) );
  CLKINVX3 U8390 ( .A(n2566), .Y(n2564) );
  CLKINVX3 U8391 ( .A(n2930), .Y(n2928) );
  CLKINVX3 U8392 ( .A(n3290), .Y(n3288) );
  CLKINVX3 U8393 ( .A(n2991), .Y(n2989) );
  CLKINVX3 U8394 ( .A(n2688), .Y(n2686) );
  CLKINVX3 U8395 ( .A(n3351), .Y(n3349) );
  CLKINVX3 U8396 ( .A(n3049), .Y(n3047) );
  CLKINVX3 U8397 ( .A(n2749), .Y(n2746) );
  CLKINVX3 U8398 ( .A(n3409), .Y(n3407) );
  CLKINVX3 U8399 ( .A(n3110), .Y(n3108) );
  CLKINVX3 U8400 ( .A(n2809), .Y(n2807) );
  BUFX3 U8401 ( .A(n625), .Y(n1221) );
  BUFX3 U8402 ( .A(n626), .Y(n1215) );
  BUFX3 U8403 ( .A(n627), .Y(n1183) );
  BUFX3 U8404 ( .A(n629), .Y(n1172) );
  BUFX3 U8405 ( .A(n628), .Y(n1175) );
  BUFX3 U8406 ( .A(n630), .Y(n1212) );
  BUFX3 U8407 ( .A(n631), .Y(n1180) );
  BUFX3 U8408 ( .A(n632), .Y(n1218) );
  CLKINVX3 U8409 ( .A(n4021), .Y(n4020) );
  XOR2X1 U8410 ( .A(top_core_EC_mc_n682), .B(top_core_EC_mc_n926), .Y(
        top_core_EC_mc_n925) );
  XOR2X1 U8411 ( .A(top_core_EC_mc_n448), .B(top_core_EC_mc_n561), .Y(
        top_core_EC_mc_n560) );
  XOR2X1 U8412 ( .A(top_core_EC_mc_n383), .B(top_core_EC_mc_n505), .Y(
        top_core_EC_mc_n504) );
  XOR2X1 U8413 ( .A(top_core_EC_mc_n577), .B(top_core_EC_mc_n695), .Y(
        top_core_EC_mc_n694) );
  XOR2X1 U8414 ( .A(top_core_EC_mc_n391), .B(top_core_EC_mc_n513), .Y(
        top_core_EC_mc_n512) );
  XOR2X1 U8415 ( .A(top_core_EC_mc_n360), .B(top_core_EC_mc_n481), .Y(
        top_core_EC_mc_n480) );
  XOR2X1 U8416 ( .A(top_core_EC_mc_n327), .B(top_core_EC_mc_n466), .Y(
        top_core_EC_mc_n465) );
  XOR2X1 U8417 ( .A(top_core_EC_mc_n92), .B(top_core_EC_mc_n222), .Y(
        top_core_EC_mc_n221) );
  XOR2X1 U8418 ( .A(top_core_EC_mc_n68), .B(top_core_EC_mc_n207), .Y(
        top_core_EC_mc_n206) );
  XOR2X1 U8419 ( .A(top_core_EC_mc_n756), .B(top_core_EC_mc_n873), .Y(
        top_core_EC_mc_n872) );
  XOR2X1 U8420 ( .A(top_core_EC_mc_n733), .B(top_core_EC_mc_n856), .Y(
        top_core_EC_mc_n855) );
  XOR2X1 U8421 ( .A(top_core_EC_mc_n423), .B(top_core_EC_mc_n545), .Y(
        top_core_EC_mc_n544) );
  XOR2X1 U8422 ( .A(top_core_EC_mc_n399), .B(top_core_EC_mc_n521), .Y(
        top_core_EC_mc_n520) );
  XOR2X1 U8423 ( .A(top_core_EC_mc_n440), .B(top_core_EC_mc_n553), .Y(
        top_core_EC_mc_n552) );
  XOR2X1 U8424 ( .A(top_core_EC_mc_n415), .B(top_core_EC_mc_n537), .Y(
        top_core_EC_mc_n536) );
  XOR2X1 U8425 ( .A(top_core_EC_mc_n407), .B(top_core_EC_mc_n529), .Y(
        top_core_EC_mc_n528) );
  XOR2X1 U8426 ( .A(top_core_EC_mc_n352), .B(top_core_EC_mc_n476), .Y(
        top_core_EC_mc_n475) );
  XOR2X1 U8427 ( .A(top_core_EC_mc_n351), .B(top_core_EC_mc_n352), .Y(
        top_core_EC_mc_n350) );
  XOR2X1 U8428 ( .A(top_core_EC_mc_n326), .B(top_core_EC_mc_n327), .Y(
        top_core_EC_mc_n325) );
  XOR2X1 U8429 ( .A(top_core_EC_mc_n84), .B(top_core_EC_mc_n217), .Y(
        top_core_EC_mc_n216) );
  XOR2X1 U8430 ( .A(top_core_EC_mc_n763), .B(top_core_EC_mc_n880), .Y(
        top_core_EC_mc_n879) );
  XOR2X1 U8431 ( .A(top_core_EC_mc_n656), .B(top_core_EC_mc_n657), .Y(
        top_core_EC_mc_n655) );
  XOR2X1 U8432 ( .A(top_core_EC_mc_n583), .B(top_core_EC_mc_n584), .Y(
        top_core_EC_mc_n582) );
  XOR2X1 U8433 ( .A(top_core_EC_mc_n496), .B(top_core_EC_mc_n497), .Y(
        top_core_EC_mc_n495) );
  XOR2X1 U8434 ( .A(top_core_EC_mc_n431), .B(top_core_EC_mc_n432), .Y(
        top_core_EC_mc_n430) );
  XOR2X1 U8435 ( .A(top_core_EC_mc_n342), .B(top_core_EC_mc_n343), .Y(
        top_core_EC_mc_n341) );
  XOR2X1 U8436 ( .A(top_core_EC_mc_n253), .B(top_core_EC_mc_n254), .Y(
        top_core_EC_mc_n252) );
  XOR2X1 U8437 ( .A(top_core_EC_mc_n188), .B(top_core_EC_mc_n189), .Y(
        top_core_EC_mc_n187) );
  XOR2X1 U8438 ( .A(top_core_EC_mc_n99), .B(top_core_EC_mc_n100), .Y(
        top_core_EC_mc_n98) );
  XOR2X1 U8439 ( .A(top_core_EC_mc_n368), .B(top_core_EC_mc_n486), .Y(
        top_core_EC_mc_n485) );
  XOR2X1 U8440 ( .A(top_core_EC_mc_n335), .B(top_core_EC_mc_n471), .Y(
        top_core_EC_mc_n470) );
  XOR2X1 U8441 ( .A(top_core_EC_mc_n359), .B(top_core_EC_mc_n360), .Y(
        top_core_EC_mc_n358) );
  XOR2X1 U8442 ( .A(top_core_EC_mc_n334), .B(top_core_EC_mc_n335), .Y(
        top_core_EC_mc_n333) );
  XOR2X1 U8443 ( .A(top_core_EC_mc_n109), .B(top_core_EC_mc_n227), .Y(
        top_core_EC_mc_n226) );
  XOR2X1 U8444 ( .A(top_core_EC_mc_n76), .B(top_core_EC_mc_n212), .Y(
        top_core_EC_mc_n211) );
  XOR2X1 U8445 ( .A(top_core_EC_mc_n570), .B(top_core_EC_mc_n688), .Y(
        top_core_EC_mc_n687) );
  XOR2X1 U8446 ( .A(top_core_EC_mc_n108), .B(top_core_EC_mc_n109), .Y(
        top_core_EC_mc_n107) );
  XOR2X1 U8447 ( .A(top_core_EC_mc_n91), .B(top_core_EC_mc_n92), .Y(
        top_core_EC_mc_n90) );
  XOR2X1 U8448 ( .A(top_core_EC_mc_n83), .B(top_core_EC_mc_n84), .Y(
        top_core_EC_mc_n82) );
  XOR2X1 U8449 ( .A(top_core_EC_mc_n75), .B(top_core_EC_mc_n76), .Y(
        top_core_EC_mc_n74) );
  XOR2X1 U8450 ( .A(top_core_EC_mc_n67), .B(top_core_EC_mc_n68), .Y(
        top_core_EC_mc_n66) );
  XOR2X1 U8451 ( .A(top_core_EC_mc_n749), .B(top_core_EC_mc_n866), .Y(
        top_core_EC_mc_n865) );
  XOR2X1 U8452 ( .A(top_core_EC_mc_n741), .B(top_core_EC_mc_n861), .Y(
        top_core_EC_mc_n860) );
  XOR2X1 U8453 ( .A(top_core_EC_mc_n762), .B(top_core_EC_mc_n763), .Y(
        top_core_EC_mc_n761) );
  XOR2X1 U8454 ( .A(top_core_EC_mc_n755), .B(top_core_EC_mc_n756), .Y(
        top_core_EC_mc_n754) );
  XOR2X1 U8455 ( .A(top_core_EC_mc_n748), .B(top_core_EC_mc_n749), .Y(
        top_core_EC_mc_n747) );
  XOR2X1 U8456 ( .A(top_core_EC_mc_n740), .B(top_core_EC_mc_n741), .Y(
        top_core_EC_mc_n739) );
  XOR2X1 U8457 ( .A(top_core_EC_mc_n732), .B(top_core_EC_mc_n733), .Y(
        top_core_EC_mc_n731) );
  INVX1 U8458 ( .A(n17275), .Y(n5329) );
  INVX1 U8459 ( .A(n14125), .Y(n6113) );
  INVX1 U8460 ( .A(n18535), .Y(n4975) );
  INVX1 U8461 ( .A(n15385), .Y(n5801) );
  INVX1 U8462 ( .A(n15700), .Y(n5717) );
  INVX1 U8463 ( .A(n16960), .Y(n5413) );
  INVX1 U8464 ( .A(n18850), .Y(n4859) );
  INVX1 U8465 ( .A(n15070), .Y(n5877) );
  INVX1 U8466 ( .A(n16645), .Y(n5489) );
  INVX1 U8467 ( .A(n18220), .Y(n5059) );
  INVX1 U8468 ( .A(n14755), .Y(n5953) );
  INVX1 U8469 ( .A(n16330), .Y(n5565) );
  INVX1 U8470 ( .A(n17905), .Y(n5167) );
  INVX1 U8471 ( .A(n14440), .Y(n6029) );
  INVX1 U8472 ( .A(n16015), .Y(n5641) );
  INVX1 U8473 ( .A(n17590), .Y(n5245) );
  INVX1 U8474 ( .A(n13617), .Y(n6596) );
  CLKINVX3 U8475 ( .A(n3451), .Y(n3448) );
  CLKINVX3 U8476 ( .A(n2850), .Y(n2847) );
  CLKINVX3 U8477 ( .A(n2608), .Y(n2605) );
  CLKINVX3 U8478 ( .A(n3210), .Y(n3207) );
  CLKINVX3 U8479 ( .A(n2972), .Y(n2969) );
  CLKINVX3 U8480 ( .A(n2669), .Y(n2666) );
  CLKINVX3 U8481 ( .A(n3149), .Y(n3146) );
  CLKINVX3 U8482 ( .A(n3332), .Y(n3329) );
  CLKINVX3 U8483 ( .A(n3030), .Y(n3027) );
  CLKINVX3 U8484 ( .A(n2547), .Y(n2544) );
  CLKINVX3 U8485 ( .A(n2729), .Y(n2726) );
  CLKINVX3 U8486 ( .A(n3390), .Y(n3387) );
  CLKINVX3 U8487 ( .A(n2911), .Y(n2908) );
  CLKINVX3 U8488 ( .A(n3091), .Y(n3088) );
  CLKINVX3 U8489 ( .A(n2790), .Y(n2787) );
  CLKINVX3 U8490 ( .A(n3271), .Y(n3268) );
  AOI221X1 U8491 ( .A0(n1615), .A1(n562), .B0(n1004), .B1(n5348), .C0(n9964), 
        .Y(n9963) );
  AOI221X1 U8492 ( .A0(n1625), .A1(n561), .B0(n1145), .B1(n6144), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n149), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n148) );
  AOI221X1 U8493 ( .A0(n1611), .A1(n563), .B0(n948), .B1(n4994), .C0(n11132), 
        .Y(n11131) );
  AOI221X1 U8494 ( .A0(n1621), .A1(n564), .B0(n1088), .B1(n5820), .C0(n8212), 
        .Y(n8211) );
  AOI221X1 U8495 ( .A0(n1612), .A1(n565), .B0(n962), .B1(n5078), .C0(n10840), 
        .Y(n10839) );
  AOI221X1 U8496 ( .A0(n1618), .A1(n566), .B0(n1046), .B1(n5584), .C0(n9088), 
        .Y(n9087) );
  AOI221X1 U8497 ( .A0(n1624), .A1(n567), .B0(n1130), .B1(n6048), .C0(n7336), 
        .Y(n7335) );
  AOI221X1 U8498 ( .A0(n1614), .A1(n568), .B0(n990), .B1(n5264), .C0(n10256), 
        .Y(n10255) );
  AOI221X1 U8499 ( .A0(n1617), .A1(n569), .B0(n1032), .B1(n5508), .C0(n9380), 
        .Y(n9379) );
  AOI221X1 U8500 ( .A0(n1620), .A1(n570), .B0(n1074), .B1(n5736), .C0(n8504), 
        .Y(n8503) );
  AOI221X1 U8501 ( .A0(n1623), .A1(n571), .B0(n1116), .B1(n5972), .C0(n7628), 
        .Y(n7627) );
  AOI221X1 U8502 ( .A0(n1610), .A1(n572), .B0(n934), .B1(n4878), .C0(n11424), 
        .Y(n11423) );
  AOI221X1 U8503 ( .A0(n1619), .A1(n575), .B0(n1060), .B1(n5660), .C0(n8796), 
        .Y(n8795) );
  AOI221X1 U8504 ( .A0(n1622), .A1(n576), .B0(n1102), .B1(n5896), .C0(n7920), 
        .Y(n7919) );
  AOI221X1 U8505 ( .A0(n1613), .A1(n573), .B0(n976), .B1(n5186), .C0(n10548), 
        .Y(n10547) );
  AOI221X1 U8506 ( .A0(n1616), .A1(n574), .B0(n1018), .B1(n5432), .C0(n9672), 
        .Y(n9671) );
  AND2X2 U8507 ( .A(n6165), .B(n3473), .Y(n561) );
  AND2X2 U8508 ( .A(n5375), .B(n2872), .Y(n562) );
  AND2X2 U8509 ( .A(n5021), .B(n2630), .Y(n563) );
  AND2X2 U8510 ( .A(n5847), .B(n3232), .Y(n564) );
  AND2X2 U8511 ( .A(n5105), .B(n2691), .Y(n565) );
  AND2X2 U8512 ( .A(n5611), .B(n3052), .Y(n566) );
  AND2X2 U8513 ( .A(n6075), .B(n3412), .Y(n567) );
  AND2X2 U8514 ( .A(n5291), .B(n2812), .Y(n568) );
  AND2X2 U8515 ( .A(n5535), .B(n2994), .Y(n569) );
  AND2X2 U8516 ( .A(n5763), .B(n3171), .Y(n570) );
  AND2X2 U8517 ( .A(n5999), .B(n3354), .Y(n571) );
  AND2X2 U8518 ( .A(n4905), .B(n2569), .Y(n572) );
  AND2X2 U8519 ( .A(n5213), .B(n2751), .Y(n573) );
  AND2X2 U8520 ( .A(n5459), .B(n2933), .Y(n574) );
  AND2X2 U8521 ( .A(n5687), .B(n3113), .Y(n575) );
  AND2X2 U8522 ( .A(n5923), .B(n3293), .Y(n576) );
  CLKINVX3 U8523 ( .A(n3678), .Y(n3651) );
  OAI21XL U8524 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .B0(n14), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n328) );
  OAI21XL U8525 ( .A0(n9896), .A1(n9913), .B0(n15), .Y(n10142) );
  OAI21XL U8526 ( .A0(n11064), .A1(n11081), .B0(n16), .Y(n11310) );
  OAI21XL U8527 ( .A0(n8144), .A1(n8161), .B0(n17), .Y(n8390) );
  OAI21XL U8528 ( .A0(n10772), .A1(n10789), .B0(n18), .Y(n11018) );
  OAI21XL U8529 ( .A0(n9020), .A1(n9037), .B0(n19), .Y(n9266) );
  OAI21XL U8530 ( .A0(n7268), .A1(n7285), .B0(n20), .Y(n7514) );
  OAI21XL U8531 ( .A0(n10188), .A1(n10205), .B0(n21), .Y(n10434) );
  OAI21XL U8532 ( .A0(n9312), .A1(n9329), .B0(n22), .Y(n9558) );
  OAI21XL U8533 ( .A0(n8436), .A1(n8453), .B0(n23), .Y(n8682) );
  OAI21XL U8534 ( .A0(n7560), .A1(n7577), .B0(n24), .Y(n7806) );
  OAI21XL U8535 ( .A0(n11356), .A1(n11373), .B0(n25), .Y(n11602) );
  OAI21XL U8536 ( .A0(n10480), .A1(n10497), .B0(n26), .Y(n10726) );
  OAI21XL U8537 ( .A0(n9604), .A1(n9621), .B0(n27), .Y(n9850) );
  OAI21XL U8538 ( .A0(n8728), .A1(n8745), .B0(n28), .Y(n8974) );
  OAI21XL U8539 ( .A0(n7852), .A1(n7869), .B0(n29), .Y(n8098) );
  OAI2BB1XL U8540 ( .A0N(n2902), .A1N(n17175), .B0(n164), .Y(n17174) );
  OAI2BB1XL U8541 ( .A0N(n3494), .A1N(n14025), .B0(n165), .Y(n14024) );
  OAI2BB1XL U8542 ( .A0N(n2651), .A1N(n18435), .B0(n166), .Y(n18434) );
  OAI2BB1XL U8543 ( .A0N(n3262), .A1N(n15285), .B0(n167), .Y(n15284) );
  OAI2BB1XL U8544 ( .A0N(n3201), .A1N(n15600), .B0(n168), .Y(n15599) );
  OAI2BB1XL U8545 ( .A0N(n2590), .A1N(n18750), .B0(n169), .Y(n18749) );
  OAI2BB1XL U8546 ( .A0N(n2963), .A1N(n16860), .B0(n170), .Y(n16859) );
  OAI2BB1XL U8547 ( .A0N(top_core_EC_ss_in[24]), .A1N(n14970), .B0(n171), .Y(
        n14969) );
  OAI2BB1XL U8548 ( .A0N(n3016), .A1N(n16545), .B0(n172), .Y(n16544) );
  OAI2BB1XL U8549 ( .A0N(n2711), .A1N(n18120), .B0(n173), .Y(n18119) );
  OAI2BB1XL U8550 ( .A0N(n3376), .A1N(n14655), .B0(n174), .Y(n14654) );
  OAI2BB1XL U8551 ( .A0N(n3073), .A1N(n16230), .B0(n175), .Y(n16229) );
  OAI2BB1XL U8552 ( .A0N(n2773), .A1N(n17805), .B0(n176), .Y(n17804) );
  OAI2BB1XL U8553 ( .A0N(n3433), .A1N(n14340), .B0(n177), .Y(n14339) );
  OAI2BB1XL U8554 ( .A0N(n3135), .A1N(n15915), .B0(n178), .Y(n15914) );
  OAI2BB1XL U8555 ( .A0N(n2834), .A1N(n17490), .B0(n179), .Y(n17489) );
  AOI211X1 U8556 ( .A0(n3483), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n298), 
        .B0(n1139), .C0(top_core_EC_ss_gen_tbox_0__sboxs_r_n86), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n312) );
  AOI211X1 U8557 ( .A0(n2882), .A1(n10112), .B0(n996), .C0(n9903), .Y(n10126)
         );
  AOI211X1 U8558 ( .A0(n2640), .A1(n11280), .B0(n940), .C0(n11071), .Y(n11294)
         );
  AOI211X1 U8559 ( .A0(n3242), .A1(n8360), .B0(n1080), .C0(n8151), .Y(n8374)
         );
  AOI211X1 U8560 ( .A0(n2701), .A1(n10988), .B0(n954), .C0(n10779), .Y(n11002)
         );
  AOI211X1 U8561 ( .A0(n3062), .A1(n9236), .B0(n1038), .C0(n9027), .Y(n9250)
         );
  AOI211X1 U8562 ( .A0(n3422), .A1(n7484), .B0(n1122), .C0(n7275), .Y(n7498)
         );
  AOI211X1 U8563 ( .A0(n2822), .A1(n10404), .B0(n982), .C0(n10195), .Y(n10418)
         );
  AOI211X1 U8564 ( .A0(n3004), .A1(n9528), .B0(n1024), .C0(n9319), .Y(n9542)
         );
  AOI211X1 U8565 ( .A0(n3181), .A1(n8652), .B0(n1066), .C0(n8443), .Y(n8666)
         );
  AOI211X1 U8566 ( .A0(n3364), .A1(n7776), .B0(n1108), .C0(n7567), .Y(n7790)
         );
  AOI211X1 U8567 ( .A0(n2579), .A1(n11572), .B0(n926), .C0(n11363), .Y(n11586)
         );
  AOI211X1 U8568 ( .A0(n2761), .A1(n10696), .B0(n968), .C0(n10487), .Y(n10710)
         );
  AOI211X1 U8569 ( .A0(n2943), .A1(n9820), .B0(n1010), .C0(n9611), .Y(n9834)
         );
  AOI211X1 U8570 ( .A0(n3123), .A1(n8944), .B0(n1052), .C0(n8735), .Y(n8958)
         );
  AOI211X1 U8571 ( .A0(n3303), .A1(n8068), .B0(n1094), .C0(n7859), .Y(n8082)
         );
  AOI211X1 U8572 ( .A0(n17057), .A1(n2904), .B0(n17058), .C0(n17059), .Y(
        n17055) );
  AOI211X1 U8573 ( .A0(n13907), .A1(n3507), .B0(n13908), .C0(n13909), .Y(
        n13905) );
  AOI211X1 U8574 ( .A0(n18317), .A1(n2662), .B0(n18318), .C0(n18319), .Y(
        n18315) );
  AOI211X1 U8575 ( .A0(n15167), .A1(n3264), .B0(n15168), .C0(n15169), .Y(
        n15165) );
  AOI211X1 U8576 ( .A0(n15482), .A1(n3203), .B0(n15483), .C0(n15484), .Y(
        n15480) );
  AOI211X1 U8577 ( .A0(n18632), .A1(n2601), .B0(n18633), .C0(n18634), .Y(
        n18630) );
  AOI211X1 U8578 ( .A0(n16742), .A1(n2965), .B0(n16743), .C0(n16744), .Y(
        n16740) );
  AOI211X1 U8579 ( .A0(n14852), .A1(n3327), .B0(n14853), .C0(n14854), .Y(
        n14850) );
  AOI211X1 U8580 ( .A0(n16427), .A1(n3024), .B0(n16428), .C0(n16429), .Y(
        n16425) );
  AOI211X1 U8581 ( .A0(n18002), .A1(n2722), .B0(n18003), .C0(n18004), .Y(
        n18000) );
  AOI211X1 U8582 ( .A0(n14537), .A1(n3384), .B0(n14538), .C0(n14539), .Y(
        n14535) );
  AOI211X1 U8583 ( .A0(n16112), .A1(n3084), .B0(n16113), .C0(n16114), .Y(
        n16110) );
  AOI211X1 U8584 ( .A0(n17687), .A1(n2785), .B0(n17688), .C0(n17689), .Y(
        n17685) );
  AOI211X1 U8585 ( .A0(n14222), .A1(n3444), .B0(n14223), .C0(n14224), .Y(
        n14220) );
  AOI211X1 U8586 ( .A0(n15797), .A1(n3143), .B0(n15798), .C0(n15799), .Y(
        n15795) );
  AOI211X1 U8587 ( .A0(n17372), .A1(n2845), .B0(n17373), .C0(n17374), .Y(
        n17370) );
  AOI221X1 U8588 ( .A0(n2859), .A1(n17236), .B0(n17237), .B1(n2852), .C0(
        n17238), .Y(n17210) );
  NAND4X1 U8589 ( .A(n5382), .B(n17073), .C(n17240), .D(n17241), .Y(n17237) );
  OAI221XL U8590 ( .A0(n1003), .A1(n17031), .B0(n17007), .B1(n17239), .C0(
        n17032), .Y(n17238) );
  AOI221X1 U8591 ( .A0(n3455), .A1(n14086), .B0(n14087), .B1(n3453), .C0(
        n14088), .Y(n14060) );
  NAND4X1 U8592 ( .A(n6153), .B(n13923), .C(n14090), .D(n14091), .Y(n14087) );
  OAI221XL U8593 ( .A0(n1142), .A1(n13881), .B0(n13857), .B1(n14089), .C0(
        n13882), .Y(n14088) );
  AOI221X1 U8594 ( .A0(n3219), .A1(n15346), .B0(n15347), .B1(n3212), .C0(
        n15348), .Y(n15320) );
  NAND4X1 U8595 ( .A(n5854), .B(n15183), .C(n15350), .D(n15351), .Y(n15347) );
  OAI221XL U8596 ( .A0(n1087), .A1(n15141), .B0(n15117), .B1(n15349), .C0(
        n15142), .Y(n15348) );
  AOI221X1 U8597 ( .A0(n2618), .A1(n18496), .B0(n18497), .B1(n2622), .C0(
        n18498), .Y(n18470) );
  NAND4X1 U8598 ( .A(n5028), .B(n18333), .C(n18500), .D(n18501), .Y(n18497) );
  OAI221XL U8599 ( .A0(n947), .A1(n18291), .B0(n18267), .B1(n18499), .C0(
        n18292), .Y(n18498) );
  AOI221X1 U8600 ( .A0(n3159), .A1(n15661), .B0(n15662), .B1(n3151), .C0(
        n15663), .Y(n15635) );
  NAND4X1 U8601 ( .A(n5770), .B(n15498), .C(n15665), .D(n15666), .Y(n15662) );
  OAI221XL U8602 ( .A0(n1073), .A1(n15456), .B0(n15432), .B1(n15664), .C0(
        n15457), .Y(n15663) );
  AOI221X1 U8603 ( .A0(n2921), .A1(n16921), .B0(n16922), .B1(n2913), .C0(
        n16923), .Y(n16895) );
  NAND4X1 U8604 ( .A(n5466), .B(n16758), .C(n16925), .D(n16926), .Y(n16922) );
  OAI221XL U8605 ( .A0(n1017), .A1(n16716), .B0(n16692), .B1(n16924), .C0(
        n16717), .Y(n16923) );
  AOI221X1 U8606 ( .A0(n2559), .A1(n18811), .B0(n18812), .B1(n2548), .C0(
        n18813), .Y(n18785) );
  NAND4X1 U8607 ( .A(n4912), .B(n18648), .C(n18815), .D(n18816), .Y(n18812) );
  OAI221XL U8608 ( .A0(n933), .A1(n18606), .B0(n18582), .B1(n18814), .C0(
        n18607), .Y(n18813) );
  AOI221X1 U8609 ( .A0(n3281), .A1(n15031), .B0(n15032), .B1(n3273), .C0(
        n15033), .Y(n15005) );
  NAND4X1 U8610 ( .A(n5930), .B(n14868), .C(n15035), .D(n15036), .Y(n15032) );
  OAI221XL U8611 ( .A0(n1101), .A1(n14826), .B0(n14802), .B1(n15034), .C0(
        n14827), .Y(n15033) );
  AOI221X1 U8612 ( .A0(n2982), .A1(n16606), .B0(n16607), .B1(n2974), .C0(
        n16608), .Y(n16580) );
  NAND4X1 U8613 ( .A(n5542), .B(n16443), .C(n16610), .D(n16611), .Y(n16607) );
  OAI221XL U8614 ( .A0(n1031), .A1(n16401), .B0(n16377), .B1(n16609), .C0(
        n16402), .Y(n16608) );
  AOI221X1 U8615 ( .A0(n2678), .A1(n18181), .B0(n18182), .B1(n2671), .C0(
        n18183), .Y(n18155) );
  NAND4X1 U8616 ( .A(n5112), .B(n18018), .C(n18185), .D(n18186), .Y(n18182) );
  OAI221XL U8617 ( .A0(n961), .A1(n17976), .B0(n17952), .B1(n18184), .C0(
        n17977), .Y(n18183) );
  AOI221X1 U8618 ( .A0(n3342), .A1(n14716), .B0(n14717), .B1(n3346), .C0(
        n14718), .Y(n14690) );
  NAND4X1 U8619 ( .A(n6006), .B(n14553), .C(n14720), .D(n14721), .Y(n14717) );
  OAI221XL U8620 ( .A0(n1115), .A1(n14511), .B0(n14487), .B1(n14719), .C0(
        n14512), .Y(n14718) );
  AOI221X1 U8621 ( .A0(n3040), .A1(n16291), .B0(n16292), .B1(n3044), .C0(
        n16293), .Y(n16265) );
  NAND4X1 U8622 ( .A(n5618), .B(n16128), .C(n16295), .D(n16296), .Y(n16292) );
  OAI221XL U8623 ( .A0(n1045), .A1(n16086), .B0(n16062), .B1(n16294), .C0(
        n16087), .Y(n16293) );
  AOI221X1 U8624 ( .A0(n2738), .A1(n17866), .B0(n17867), .B1(n2731), .C0(
        n17868), .Y(n17840) );
  NAND4X1 U8625 ( .A(n5220), .B(n17703), .C(n17870), .D(n17871), .Y(n17867) );
  OAI221XL U8626 ( .A0(n975), .A1(n17661), .B0(n17637), .B1(n17869), .C0(
        n17662), .Y(n17868) );
  AOI221X1 U8627 ( .A0(n3400), .A1(n14401), .B0(n14402), .B1(n3404), .C0(
        n14403), .Y(n14375) );
  NAND4X1 U8628 ( .A(n6082), .B(n14238), .C(n14405), .D(n14406), .Y(n14402) );
  OAI221XL U8629 ( .A0(n1129), .A1(n14196), .B0(n14172), .B1(n14404), .C0(
        n14197), .Y(n14403) );
  AOI221X1 U8630 ( .A0(n3100), .A1(n15976), .B0(n15977), .B1(n3093), .C0(
        n15978), .Y(n15950) );
  NAND4X1 U8631 ( .A(n5694), .B(n15813), .C(n15980), .D(n15981), .Y(n15977) );
  OAI221XL U8632 ( .A0(n1059), .A1(n15771), .B0(n15747), .B1(n15979), .C0(
        n15772), .Y(n15978) );
  AOI221X1 U8633 ( .A0(n2800), .A1(n17551), .B0(n17552), .B1(n2792), .C0(
        n17553), .Y(n17525) );
  NAND4X1 U8634 ( .A(n5298), .B(n17388), .C(n17555), .D(n17556), .Y(n17552) );
  OAI221XL U8635 ( .A0(n989), .A1(n17346), .B0(n17322), .B1(n17554), .C0(
        n17347), .Y(n17553) );
  AOI222X1 U8636 ( .A0(n5333), .A1(n586), .B0(n2857), .B1(n10042), .C0(n10043), 
        .C1(n2853), .Y(n10023) );
  NAND4BXL U8637 ( .AN(n10044), .B(n10045), .C(n10046), .D(n10047), .Y(n10043)
         );
  AOI222X1 U8638 ( .A0(n5375), .A1(n2901), .B0(n5366), .B1(n433), .C0(n1001), 
        .C1(n5347), .Y(n10047) );
  AOI222X1 U8639 ( .A0(n6119), .A1(n585), .B0(n3462), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n228), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n229), .C1(n3454), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n209) );
  NAND4BXL U8640 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n230), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n231), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n232), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n233), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n229) );
  AOI222X1 U8641 ( .A0(n6165), .A1(n3500), .B0(n6156), .B1(n434), .C0(n1143), 
        .C1(n6143), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n233) );
  AOI222X1 U8642 ( .A0(n4979), .A1(n587), .B0(n2612), .B1(n11210), .C0(n11211), 
        .C1(n2611), .Y(n11191) );
  NAND4BXL U8643 ( .AN(n11212), .B(n11213), .C(n11214), .D(n11215), .Y(n11211)
         );
  AOI222X1 U8644 ( .A0(n5021), .A1(n2656), .B0(n5012), .B1(n435), .C0(n945), 
        .C1(n4993), .Y(n11215) );
  AOI222X1 U8645 ( .A0(n5805), .A1(n588), .B0(n3217), .B1(n8290), .C0(n8291), 
        .C1(n3213), .Y(n8271) );
  NAND4BXL U8646 ( .AN(n8292), .B(n8293), .C(n8294), .D(n8295), .Y(n8291) );
  AOI222X1 U8647 ( .A0(n5847), .A1(n3261), .B0(n5838), .B1(n436), .C0(n1085), 
        .C1(n5819), .Y(n8295) );
  AOI222X1 U8648 ( .A0(n5063), .A1(n589), .B0(n2676), .B1(n10918), .C0(n10919), 
        .C1(n2672), .Y(n10899) );
  NAND4BXL U8649 ( .AN(n10920), .B(n10921), .C(n10922), .D(n10923), .Y(n10919)
         );
  AOI222X1 U8650 ( .A0(n5105), .A1(n2719), .B0(n5096), .B1(n442), .C0(n959), 
        .C1(n5077), .Y(n10923) );
  AOI222X1 U8651 ( .A0(n5569), .A1(n590), .B0(n3034), .B1(n9166), .C0(n9167), 
        .C1(n3033), .Y(n9147) );
  NAND4BXL U8652 ( .AN(n9168), .B(n9169), .C(n9170), .D(n9171), .Y(n9167) );
  AOI222X1 U8653 ( .A0(n5611), .A1(n3078), .B0(n5602), .B1(n444), .C0(n1043), 
        .C1(n5583), .Y(n9171) );
  AOI222X1 U8654 ( .A0(n6033), .A1(n591), .B0(n3394), .B1(n7414), .C0(n7415), 
        .C1(n3393), .Y(n7395) );
  NAND4BXL U8655 ( .AN(n7416), .B(n7417), .C(n7418), .D(n7419), .Y(n7415) );
  AOI222X1 U8656 ( .A0(n6075), .A1(n3441), .B0(n6066), .B1(n446), .C0(n1127), 
        .C1(n6047), .Y(n7419) );
  AOI222X1 U8657 ( .A0(n5249), .A1(n592), .B0(n2794), .B1(n10334), .C0(n10335), 
        .C1(n2793), .Y(n10315) );
  NAND4BXL U8658 ( .AN(n10336), .B(n10337), .C(n10338), .D(n10339), .Y(n10335)
         );
  AOI222X1 U8659 ( .A0(n5291), .A1(n2839), .B0(n5282), .B1(n448), .C0(n987), 
        .C1(n5263), .Y(n10339) );
  AOI222X1 U8660 ( .A0(n5493), .A1(n593), .B0(n2976), .B1(n9458), .C0(n9459), 
        .C1(n2975), .Y(n9439) );
  NAND4BXL U8661 ( .AN(n9460), .B(n9461), .C(n9462), .D(n9463), .Y(n9459) );
  AOI222X1 U8662 ( .A0(n5535), .A1(n3017), .B0(n5526), .B1(n441), .C0(n1029), 
        .C1(n5507), .Y(n9463) );
  AOI222X1 U8663 ( .A0(n5721), .A1(n594), .B0(n3153), .B1(n8582), .C0(n8583), 
        .C1(n3152), .Y(n8563) );
  NAND4BXL U8664 ( .AN(n8584), .B(n8585), .C(n8586), .D(n8587), .Y(n8583) );
  AOI222X1 U8665 ( .A0(n5763), .A1(n3200), .B0(n5754), .B1(n437), .C0(n1071), 
        .C1(n5735), .Y(n8587) );
  AOI222X1 U8666 ( .A0(n5957), .A1(n595), .B0(n3336), .B1(n7706), .C0(n7707), 
        .C1(n3335), .Y(n7687) );
  NAND4BXL U8667 ( .AN(n7708), .B(n7709), .C(n7710), .D(n7711), .Y(n7707) );
  AOI222X1 U8668 ( .A0(n5999), .A1(n3377), .B0(n5990), .B1(n443), .C0(n1113), 
        .C1(n5971), .Y(n7711) );
  AOI222X1 U8669 ( .A0(n4863), .A1(n596), .B0(n2553), .B1(n11502), .C0(n11503), 
        .C1(n2550), .Y(n11483) );
  NAND4BXL U8670 ( .AN(n11504), .B(n11505), .C(n11506), .D(n11507), .Y(n11503)
         );
  AOI222X1 U8671 ( .A0(n4905), .A1(n2595), .B0(n4896), .B1(n439), .C0(n931), 
        .C1(n4877), .Y(n11507) );
  AOI222X1 U8672 ( .A0(n5171), .A1(n597), .B0(n2736), .B1(n10626), .C0(n10627), 
        .C1(n2732), .Y(n10607) );
  NAND4BXL U8673 ( .AN(n10628), .B(n10629), .C(n10630), .D(n10631), .Y(n10627)
         );
  AOI222X1 U8674 ( .A0(n5213), .A1(n2785), .B0(n5204), .B1(n445), .C0(n973), 
        .C1(n5185), .Y(n10631) );
  AOI222X1 U8675 ( .A0(n5417), .A1(n598), .B0(n2915), .B1(n9750), .C0(n9751), 
        .C1(n2914), .Y(n9731) );
  NAND4BXL U8676 ( .AN(n9752), .B(n9753), .C(n9754), .D(n9755), .Y(n9751) );
  AOI222X1 U8677 ( .A0(n5459), .A1(n2962), .B0(n5450), .B1(n438), .C0(n1015), 
        .C1(n5431), .Y(n9755) );
  AOI222X1 U8678 ( .A0(n5645), .A1(n599), .B0(n3098), .B1(n8874), .C0(n8875), 
        .C1(n3094), .Y(n8855) );
  NAND4BXL U8679 ( .AN(n8876), .B(n8877), .C(n8878), .D(n8879), .Y(n8875) );
  AOI222X1 U8680 ( .A0(n5687), .A1(n3136), .B0(n5678), .B1(n447), .C0(n1057), 
        .C1(n5659), .Y(n8879) );
  AOI222X1 U8681 ( .A0(n5881), .A1(n600), .B0(n3275), .B1(n7998), .C0(n7999), 
        .C1(n3274), .Y(n7979) );
  NAND4BXL U8682 ( .AN(n8000), .B(n8001), .C(n8002), .D(n8003), .Y(n7999) );
  AOI222X1 U8683 ( .A0(n5923), .A1(n3321), .B0(n5914), .B1(n440), .C0(n1099), 
        .C1(n5895), .Y(n8003) );
  AOI211X1 U8684 ( .A0(n5336), .A1(n1615), .B0(n5350), .C0(n10019), .Y(n10151)
         );
  AOI211X1 U8685 ( .A0(n6132), .A1(n1625), .B0(n6146), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n205), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n337) );
  AOI211X1 U8686 ( .A0(n5808), .A1(n1621), .B0(n5822), .C0(n8267), .Y(n8399)
         );
  AOI211X1 U8687 ( .A0(n4982), .A1(n1611), .B0(n4996), .C0(n11187), .Y(n11319)
         );
  AOI211X1 U8688 ( .A0(n2863), .A1(n10104), .B0(n5369), .C0(n9926), .Y(n10103)
         );
  AOI211X1 U8689 ( .A0(n3464), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n290), 
        .B0(n6159), .C0(top_core_EC_ss_gen_tbox_0__sboxs_r_n111), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n289) );
  AOI211X1 U8690 ( .A0(n3223), .A1(n8352), .B0(n5841), .C0(n8174), .Y(n8351)
         );
  AOI211X1 U8691 ( .A0(n2621), .A1(n11272), .B0(n5015), .C0(n11094), .Y(n11271) );
  AOI211X1 U8692 ( .A0(n5066), .A1(n1612), .B0(n5080), .C0(n10895), .Y(n11027)
         );
  AOI211X1 U8693 ( .A0(n6036), .A1(n1624), .B0(n6050), .C0(n7391), .Y(n7523)
         );
  AOI211X1 U8694 ( .A0(n5572), .A1(n1618), .B0(n5586), .C0(n9143), .Y(n9275)
         );
  AOI211X1 U8695 ( .A0(n2682), .A1(n10980), .B0(n5099), .C0(n10802), .Y(n10979) );
  AOI211X1 U8696 ( .A0(n5252), .A1(n1614), .B0(n5266), .C0(n10311), .Y(n10443)
         );
  AOI211X1 U8697 ( .A0(n5496), .A1(n1617), .B0(n5510), .C0(n9435), .Y(n9567)
         );
  AOI211X1 U8698 ( .A0(n5724), .A1(n1620), .B0(n5738), .C0(n8559), .Y(n8691)
         );
  AOI211X1 U8699 ( .A0(n5960), .A1(n1623), .B0(n5974), .C0(n7683), .Y(n7815)
         );
  AOI211X1 U8700 ( .A0(n4866), .A1(n1610), .B0(n4880), .C0(n11479), .Y(n11611)
         );
  AOI211X1 U8701 ( .A0(n5174), .A1(n1613), .B0(n5188), .C0(n10603), .Y(n10735)
         );
  AOI211X1 U8702 ( .A0(n5420), .A1(n1616), .B0(n5434), .C0(n9727), .Y(n9859)
         );
  AOI211X1 U8703 ( .A0(n5648), .A1(n1619), .B0(n5662), .C0(n8851), .Y(n8983)
         );
  AOI211X1 U8704 ( .A0(n5884), .A1(n1622), .B0(n5898), .C0(n7975), .Y(n8107)
         );
  AOI211X1 U8705 ( .A0(n3403), .A1(n7476), .B0(n6069), .C0(n7298), .Y(n7475)
         );
  AOI211X1 U8706 ( .A0(n3043), .A1(n9228), .B0(n5605), .C0(n9050), .Y(n9227)
         );
  AOI211X1 U8707 ( .A0(n2803), .A1(n10396), .B0(n5285), .C0(n10218), .Y(n10395) );
  AOI211X1 U8708 ( .A0(n2985), .A1(n9520), .B0(n5529), .C0(n9342), .Y(n9519)
         );
  AOI211X1 U8709 ( .A0(n3162), .A1(n8644), .B0(n5757), .C0(n8466), .Y(n8643)
         );
  AOI211X1 U8710 ( .A0(n3345), .A1(n7768), .B0(n5993), .C0(n7590), .Y(n7767)
         );
  AOI211X1 U8711 ( .A0(n2560), .A1(n11564), .B0(n4899), .C0(n11386), .Y(n11563) );
  AOI211X1 U8712 ( .A0(n2742), .A1(n10688), .B0(n5207), .C0(n10510), .Y(n10687) );
  AOI211X1 U8713 ( .A0(n2924), .A1(n9812), .B0(n5453), .C0(n9634), .Y(n9811)
         );
  AOI211X1 U8714 ( .A0(n3104), .A1(n8936), .B0(n5681), .C0(n8758), .Y(n8935)
         );
  AOI211X1 U8715 ( .A0(n3284), .A1(n8060), .B0(n5917), .C0(n7882), .Y(n8059)
         );
  INVX1 U8716 ( .A(n9949), .Y(n5342) );
  INVX1 U8717 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n134), .Y(n6138) );
  INVX1 U8718 ( .A(n11117), .Y(n4988) );
  INVX1 U8719 ( .A(n8197), .Y(n5814) );
  INVX1 U8720 ( .A(n10825), .Y(n5072) );
  INVX1 U8721 ( .A(n9073), .Y(n5578) );
  INVX1 U8722 ( .A(n7321), .Y(n6042) );
  INVX1 U8723 ( .A(n10241), .Y(n5258) );
  INVX1 U8724 ( .A(n9365), .Y(n5502) );
  INVX1 U8725 ( .A(n8489), .Y(n5730) );
  INVX1 U8726 ( .A(n7613), .Y(n5966) );
  INVX1 U8727 ( .A(n11409), .Y(n4872) );
  INVX1 U8728 ( .A(n10533), .Y(n5180) );
  INVX1 U8729 ( .A(n9657), .Y(n5426) );
  INVX1 U8730 ( .A(n8781), .Y(n5654) );
  INVX1 U8731 ( .A(n7905), .Y(n5890) );
  INVX1 U8732 ( .A(n17028), .Y(n5352) );
  INVX1 U8733 ( .A(n13878), .Y(n6120) );
  INVX1 U8734 ( .A(n18288), .Y(n4998) );
  INVX1 U8735 ( .A(n15138), .Y(n5824) );
  INVX1 U8736 ( .A(n15453), .Y(n5740) );
  INVX1 U8737 ( .A(n18603), .Y(n4882) );
  INVX1 U8738 ( .A(n16713), .Y(n5436) );
  INVX1 U8739 ( .A(n14823), .Y(n5900) );
  INVX1 U8740 ( .A(n16398), .Y(n5512) );
  INVX1 U8741 ( .A(n17973), .Y(n5082) );
  INVX1 U8742 ( .A(n14508), .Y(n5976) );
  INVX1 U8743 ( .A(n16083), .Y(n5588) );
  INVX1 U8744 ( .A(n17658), .Y(n5190) );
  INVX1 U8745 ( .A(n14193), .Y(n6052) );
  INVX1 U8746 ( .A(n15768), .Y(n5664) );
  INVX1 U8747 ( .A(n17343), .Y(n5268) );
  INVX1 U8748 ( .A(n2889), .Y(n2885) );
  INVX1 U8749 ( .A(n3505), .Y(n3496) );
  INVX1 U8750 ( .A(n3490), .Y(n3486) );
  INVX1 U8751 ( .A(n3505), .Y(n3497) );
  INVX1 U8752 ( .A(n2906), .Y(n2894) );
  INVX1 U8753 ( .A(n3266), .Y(n3254) );
  INVX1 U8754 ( .A(n3205), .Y(n3193) );
  INVX1 U8755 ( .A(n2967), .Y(n2955) );
  INVX1 U8756 ( .A(top_core_EC_ss_in[96]), .Y(n2777) );
  INVX1 U8757 ( .A(n3325), .Y(n3318) );
  INVX1 U8758 ( .A(n2516), .Y(n2421) );
  INVX1 U8759 ( .A(n2520), .Y(n2403) );
  INVX1 U8760 ( .A(n2516), .Y(n2422) );
  INVX1 U8761 ( .A(n2382), .Y(n2412) );
  INVX1 U8762 ( .A(n2519), .Y(n2407) );
  INVX1 U8763 ( .A(n2380), .Y(n2413) );
  INVX1 U8764 ( .A(n2386), .Y(n2410) );
  INVX1 U8765 ( .A(n2517), .Y(n2418) );
  INVX1 U8766 ( .A(n2520), .Y(n2404) );
  INVX1 U8767 ( .A(top_core_EC_operation), .Y(n2400) );
  INVX1 U8768 ( .A(n2518), .Y(n2415) );
  INVX1 U8769 ( .A(n2388), .Y(n2409) );
  INVX1 U8770 ( .A(n2515), .Y(n2424) );
  INVX1 U8771 ( .A(n2387), .Y(n2408) );
  INVX1 U8772 ( .A(n2517), .Y(n2419) );
  INVX1 U8773 ( .A(n2515), .Y(n2423) );
  INVX1 U8774 ( .A(n2519), .Y(n2405) );
  INVX1 U8775 ( .A(n2518), .Y(n2416) );
  INVX1 U8776 ( .A(n2517), .Y(n2417) );
  INVX1 U8777 ( .A(n2378), .Y(n2411) );
  INVX1 U8778 ( .A(n2515), .Y(n2425) );
  INVX1 U8779 ( .A(n2518), .Y(n2414) );
  INVX1 U8780 ( .A(n2520), .Y(n2402) );
  INVX1 U8781 ( .A(n2383), .Y(n2401) );
  INVX1 U8782 ( .A(n2516), .Y(n2420) );
  INVX1 U8783 ( .A(n2519), .Y(n2406) );
  INVX1 U8784 ( .A(n2514), .Y(n2427) );
  INVX1 U8785 ( .A(n2514), .Y(n2428) );
  INVX1 U8786 ( .A(n2514), .Y(n2426) );
  INVX1 U8787 ( .A(n2865), .Y(n2855) );
  INVX1 U8788 ( .A(n3225), .Y(n3215) );
  INVX1 U8789 ( .A(n2610), .Y(n2613) );
  INVX1 U8790 ( .A(n3466), .Y(n3456) );
  INVX1 U8791 ( .A(n2684), .Y(n2674) );
  INVX1 U8792 ( .A(n3392), .Y(n3395) );
  INVX1 U8793 ( .A(n3032), .Y(n3035) );
  INVX1 U8794 ( .A(n2805), .Y(n2795) );
  INVX1 U8795 ( .A(n2987), .Y(n2977) );
  INVX1 U8796 ( .A(n3164), .Y(n3154) );
  INVX1 U8797 ( .A(n3334), .Y(n3337) );
  INVX1 U8798 ( .A(n2562), .Y(n2552) );
  INVX1 U8799 ( .A(n2744), .Y(n2734) );
  INVX1 U8800 ( .A(n2926), .Y(n2916) );
  INVX1 U8801 ( .A(n3106), .Y(n3096) );
  INVX1 U8802 ( .A(n3286), .Y(n3276) );
  INVX1 U8803 ( .A(n2864), .Y(n2856) );
  INVX1 U8804 ( .A(n3224), .Y(n3216) );
  INVX1 U8805 ( .A(n2683), .Y(n2675) );
  INVX1 U8806 ( .A(n2743), .Y(n2735) );
  INVX1 U8807 ( .A(n3105), .Y(n3097) );
  INVX1 U8808 ( .A(n3505), .Y(n3495) );
  INVX1 U8809 ( .A(n2844), .Y(n2835) );
  INVX1 U8810 ( .A(n2720), .Y(n2712) );
  INVX1 U8811 ( .A(n3442), .Y(n3434) );
  INVX1 U8812 ( .A(n3326), .Y(n3315) );
  INVX1 U8813 ( .A(n2784), .Y(n2774) );
  INVX1 U8814 ( .A(n2844), .Y(n2836) );
  INVX1 U8815 ( .A(n3016), .Y(n3017) );
  INVX1 U8816 ( .A(n3376), .Y(n3377) );
  INVX1 U8817 ( .A(n2784), .Y(n2775) );
  INVX1 U8818 ( .A(n3135), .Y(n3136) );
  INVX1 U8819 ( .A(n3326), .Y(n3316) );
  INVX1 U8820 ( .A(n3465), .Y(n3457) );
  INVX1 U8821 ( .A(n2623), .Y(n2614) );
  INVX1 U8822 ( .A(n3163), .Y(n3155) );
  INVX1 U8823 ( .A(n2925), .Y(n2917) );
  INVX1 U8824 ( .A(n2561), .Y(n2553) );
  INVX1 U8825 ( .A(n3285), .Y(n3277) );
  INVX1 U8826 ( .A(n2986), .Y(n2978) );
  INVX1 U8827 ( .A(n3347), .Y(n3338) );
  INVX1 U8828 ( .A(n3045), .Y(n3036) );
  INVX1 U8829 ( .A(n3405), .Y(n3396) );
  INVX1 U8830 ( .A(n2804), .Y(n2796) );
  INVX1 U8831 ( .A(n2852), .Y(n2857) );
  INVX1 U8832 ( .A(n3453), .Y(n3458) );
  INVX1 U8833 ( .A(n2610), .Y(n2615) );
  INVX1 U8834 ( .A(n3212), .Y(n3217) );
  INVX1 U8835 ( .A(n3151), .Y(n3156) );
  INVX1 U8836 ( .A(n2913), .Y(n2918) );
  INVX1 U8837 ( .A(n2549), .Y(n2554) );
  INVX1 U8838 ( .A(n3273), .Y(n3278) );
  INVX1 U8839 ( .A(n2974), .Y(n2979) );
  INVX1 U8840 ( .A(n3334), .Y(n3339) );
  INVX1 U8841 ( .A(n2731), .Y(n2736) );
  INVX1 U8842 ( .A(n3093), .Y(n3098) );
  INVX1 U8843 ( .A(n2671), .Y(n2676) );
  INVX1 U8844 ( .A(n3032), .Y(n3037) );
  INVX1 U8845 ( .A(n3392), .Y(n3397) );
  INVX1 U8846 ( .A(n2792), .Y(n2797) );
  INVX1 U8847 ( .A(top_core_EC_ss_in[81]), .Y(n2883) );
  INVX1 U8848 ( .A(n2647), .Y(n2641) );
  INVX1 U8849 ( .A(n2724), .Y(n2713) );
  INVX1 U8850 ( .A(n3446), .Y(n3435) );
  INVX1 U8851 ( .A(n3429), .Y(n3423) );
  INVX1 U8852 ( .A(n3069), .Y(n3063) );
  INVX1 U8853 ( .A(n2844), .Y(n2837) );
  INVX1 U8854 ( .A(n2829), .Y(n2823) );
  INVX1 U8855 ( .A(n3016), .Y(n3018) );
  INVX1 U8856 ( .A(n3376), .Y(n3378) );
  INVX1 U8857 ( .A(n2784), .Y(n2776) );
  INVX1 U8858 ( .A(n2950), .Y(n2944) );
  INVX1 U8859 ( .A(n3135), .Y(n3137) );
  INVX1 U8860 ( .A(n3326), .Y(n3317) );
  INVX1 U8861 ( .A(n3481), .Y(n3484) );
  INVX1 U8862 ( .A(n2880), .Y(n2884) );
  INVX1 U8863 ( .A(n3240), .Y(n3243) );
  INVX1 U8864 ( .A(n3301), .Y(n3304) );
  INVX1 U8865 ( .A(n3002), .Y(n3005) );
  INVX1 U8866 ( .A(n3480), .Y(n3477) );
  INVX1 U8867 ( .A(n3473), .Y(n3478) );
  INVX1 U8868 ( .A(n2872), .Y(n2875) );
  INVX1 U8869 ( .A(n2630), .Y(n2633) );
  INVX1 U8870 ( .A(n3232), .Y(n3236) );
  INVX1 U8871 ( .A(n2932), .Y(n2936) );
  INVX1 U8872 ( .A(n3171), .Y(n3175) );
  INVX1 U8873 ( .A(n2569), .Y(n2572) );
  INVX1 U8874 ( .A(n2993), .Y(n2997) );
  INVX1 U8875 ( .A(n3113), .Y(n3116) );
  INVX1 U8876 ( .A(n2690), .Y(n2694) );
  INVX1 U8877 ( .A(n3052), .Y(n3055) );
  INVX1 U8878 ( .A(n3411), .Y(n3415) );
  INVX1 U8879 ( .A(n3354), .Y(n3358) );
  INVX1 U8880 ( .A(n2751), .Y(n2755) );
  INVX1 U8881 ( .A(n3490), .Y(n3485) );
  INVX1 U8882 ( .A(n2882), .Y(n2886) );
  INVX1 U8883 ( .A(n3249), .Y(n3244) );
  INVX1 U8884 ( .A(n3189), .Y(n3182) );
  INVX1 U8885 ( .A(n2950), .Y(n2945) );
  INVX1 U8886 ( .A(n2587), .Y(n2580) );
  INVX1 U8887 ( .A(n3310), .Y(n3305) );
  INVX1 U8888 ( .A(n3011), .Y(n3006) );
  INVX1 U8889 ( .A(n2701), .Y(n2702) );
  INVX1 U8890 ( .A(n3372), .Y(n3365) );
  INVX1 U8891 ( .A(n3069), .Y(n3064) );
  INVX1 U8892 ( .A(n2769), .Y(n2762) );
  INVX1 U8893 ( .A(n3131), .Y(n3124) );
  INVX1 U8894 ( .A(n2829), .Y(n2824) );
  INVX1 U8895 ( .A(n2871), .Y(n2876) );
  INVX1 U8896 ( .A(n2629), .Y(n2634) );
  INVX1 U8897 ( .A(n2690), .Y(n2695) );
  INVX1 U8898 ( .A(n3411), .Y(n3416) );
  INVX1 U8899 ( .A(n3051), .Y(n3056) );
  INVX1 U8900 ( .A(n2932), .Y(n2937) );
  INVX1 U8901 ( .A(n2819), .Y(n2815) );
  INVX1 U8902 ( .A(n2568), .Y(n2573) );
  INVX1 U8903 ( .A(n3300), .Y(n3296) );
  INVX1 U8904 ( .A(n2993), .Y(n2998) );
  INVX1 U8905 ( .A(n3112), .Y(n3117) );
  INVX1 U8906 ( .A(n3480), .Y(n3479) );
  INVX1 U8907 ( .A(n2879), .Y(n2877) );
  INVX1 U8908 ( .A(n2637), .Y(n2635) );
  INVX1 U8909 ( .A(n3239), .Y(n3237) );
  INVX1 U8910 ( .A(n3178), .Y(n3176) );
  INVX1 U8911 ( .A(n3059), .Y(n3057) );
  INVX1 U8912 ( .A(n2819), .Y(n2816) );
  INVX1 U8913 ( .A(n2576), .Y(n2574) );
  INVX1 U8914 ( .A(n3300), .Y(n3297) );
  INVX1 U8915 ( .A(n3361), .Y(n3359) );
  INVX1 U8916 ( .A(n2758), .Y(n2756) );
  INVX1 U8917 ( .A(n3120), .Y(n3118) );
  INVX1 U8918 ( .A(n2494), .Y(n2492) );
  INVX1 U8919 ( .A(n2494), .Y(n2491) );
  INVX1 U8920 ( .A(n2495), .Y(n2490) );
  INVX1 U8921 ( .A(n2541), .Y(n2509) );
  INVX1 U8922 ( .A(n2541), .Y(n2510) );
  INVX1 U8923 ( .A(n2530), .Y(n2503) );
  INVX1 U8924 ( .A(n2530), .Y(n2504) );
  INVX1 U8925 ( .A(n2526), .Y(n2511) );
  INVX1 U8926 ( .A(n2366), .Y(n2513) );
  INVX1 U8927 ( .A(n2496), .Y(n2486) );
  INVX1 U8928 ( .A(n2496), .Y(n2485) );
  INVX1 U8929 ( .A(n2526), .Y(n2512) );
  INVX1 U8930 ( .A(n2528), .Y(n2508) );
  INVX1 U8931 ( .A(n2528), .Y(n2507) );
  INVX1 U8932 ( .A(n2529), .Y(n2506) );
  INVX1 U8933 ( .A(n2494), .Y(n2493) );
  INVX1 U8934 ( .A(n2529), .Y(n2505) );
  INVX1 U8935 ( .A(n2532), .Y(n2500) );
  INVX1 U8936 ( .A(n2531), .Y(n2501) );
  INVX1 U8937 ( .A(n2531), .Y(n2502) );
  INVX1 U8938 ( .A(n2533), .Y(n2498) );
  INVX1 U8939 ( .A(n2533), .Y(n2497) );
  INVX1 U8940 ( .A(n2495), .Y(n2489) );
  INVX1 U8941 ( .A(n2532), .Y(n2499) );
  INVX1 U8942 ( .A(n2496), .Y(n2487) );
  INVX1 U8943 ( .A(n2495), .Y(n2488) );
  INVX1 U8944 ( .A(top_core_EC_ss_in[41]), .Y(n3183) );
  INVX1 U8945 ( .A(top_core_EC_ss_in[121]), .Y(n2581) );
  INVX1 U8946 ( .A(top_core_EC_ss_in[105]), .Y(n2703) );
  INVX1 U8947 ( .A(top_core_EC_ss_in[17]), .Y(n3366) );
  INVX1 U8948 ( .A(top_core_EC_ss_in[97]), .Y(n2763) );
  INVX1 U8949 ( .A(top_core_EC_ss_in[49]), .Y(n3125) );
  INVX1 U8950 ( .A(n3465), .Y(n3459) );
  INVX1 U8951 ( .A(n2864), .Y(n2858) );
  INVX1 U8952 ( .A(n2623), .Y(n2616) );
  INVX1 U8953 ( .A(n3224), .Y(n3218) );
  INVX1 U8954 ( .A(n2683), .Y(n2677) );
  INVX1 U8955 ( .A(n3045), .Y(n3038) );
  INVX1 U8956 ( .A(n3405), .Y(n3398) );
  INVX1 U8957 ( .A(n2804), .Y(n2798) );
  INVX1 U8958 ( .A(n2986), .Y(n2980) );
  INVX1 U8959 ( .A(n3163), .Y(n3157) );
  INVX1 U8960 ( .A(n3347), .Y(n3340) );
  INVX1 U8961 ( .A(n2561), .Y(n2555) );
  INVX1 U8962 ( .A(n2743), .Y(n2737) );
  INVX1 U8963 ( .A(n2925), .Y(n2919) );
  INVX1 U8964 ( .A(n3105), .Y(n3099) );
  INVX1 U8965 ( .A(n3285), .Y(n3279) );
  INVX1 U8966 ( .A(n2851), .Y(n2859) );
  INVX1 U8967 ( .A(n3452), .Y(n3460) );
  INVX1 U8968 ( .A(n2623), .Y(n2617) );
  INVX1 U8969 ( .A(n3211), .Y(n3219) );
  INVX1 U8970 ( .A(n2670), .Y(n2678) );
  INVX1 U8971 ( .A(n3405), .Y(n3399) );
  INVX1 U8972 ( .A(n3045), .Y(n3039) );
  INVX1 U8973 ( .A(n3150), .Y(n3158) );
  INVX1 U8974 ( .A(n2561), .Y(n2556) );
  INVX1 U8975 ( .A(n2912), .Y(n2920) );
  INVX1 U8976 ( .A(n2973), .Y(n2981) );
  INVX1 U8977 ( .A(n3347), .Y(n3341) );
  INVX1 U8978 ( .A(n2730), .Y(n2738) );
  INVX1 U8979 ( .A(n3092), .Y(n3100) );
  INVX1 U8980 ( .A(n3272), .Y(n3280) );
  INVX1 U8981 ( .A(n2791), .Y(n2799) );
  INVX1 U8982 ( .A(n3466), .Y(n3461) );
  INVX1 U8983 ( .A(n2865), .Y(n2860) );
  INVX1 U8984 ( .A(n2611), .Y(n2618) );
  INVX1 U8985 ( .A(n3225), .Y(n3220) );
  INVX1 U8986 ( .A(n2684), .Y(n2679) );
  INVX1 U8987 ( .A(n3393), .Y(n3400) );
  INVX1 U8988 ( .A(n3033), .Y(n3040) );
  INVX1 U8989 ( .A(n2805), .Y(n2800) );
  INVX1 U8990 ( .A(n2987), .Y(n2982) );
  INVX1 U8991 ( .A(n3164), .Y(n3159) );
  INVX1 U8992 ( .A(n3335), .Y(n3342) );
  INVX1 U8993 ( .A(n2562), .Y(n2557) );
  INVX1 U8994 ( .A(n2744), .Y(n2739) );
  INVX1 U8995 ( .A(n2926), .Y(n2921) );
  INVX1 U8996 ( .A(n3106), .Y(n3101) );
  INVX1 U8997 ( .A(n3286), .Y(n3281) );
  INVX1 U8998 ( .A(n3465), .Y(n3462) );
  INVX1 U8999 ( .A(n2864), .Y(n2861) );
  INVX1 U9000 ( .A(n3224), .Y(n3221) );
  INVX1 U9001 ( .A(n2683), .Y(n2680) );
  INVX1 U9002 ( .A(n2743), .Y(n2740) );
  INVX1 U9003 ( .A(n3105), .Y(n3102) );
  INVX1 U9004 ( .A(n2903), .Y(n2895) );
  INVX1 U9005 ( .A(n2660), .Y(n2652) );
  INVX1 U9006 ( .A(n3263), .Y(n3255) );
  INVX1 U9007 ( .A(n3082), .Y(n3074) );
  INVX1 U9008 ( .A(top_core_EC_ss_in[64]), .Y(n3019) );
  INVX1 U9009 ( .A(top_core_EC_ss_in[16]), .Y(n3379) );
  INVX1 U9010 ( .A(n2783), .Y(n2778) );
  INVX1 U9011 ( .A(top_core_EC_ss_in[48]), .Y(n3138) );
  INVX1 U9012 ( .A(n2844), .Y(n2838) );
  INVX1 U9013 ( .A(n3202), .Y(n3194) );
  INVX1 U9014 ( .A(n2599), .Y(n2591) );
  INVX1 U9015 ( .A(n2964), .Y(n2956) );
  INVX1 U9016 ( .A(n2903), .Y(n2896) );
  INVX1 U9017 ( .A(n2660), .Y(n2653) );
  INVX1 U9018 ( .A(n3263), .Y(n3256) );
  INVX1 U9019 ( .A(n3202), .Y(n3195) );
  INVX1 U9020 ( .A(n2964), .Y(n2957) );
  INVX1 U9021 ( .A(n2932), .Y(n2938) );
  INVX1 U9022 ( .A(n2690), .Y(n2696) );
  INVX1 U9023 ( .A(n3411), .Y(n3417) );
  INVX1 U9024 ( .A(n2599), .Y(n2592) );
  INVX1 U9025 ( .A(n3292), .Y(n3298) );
  INVX1 U9026 ( .A(top_core_EC_ss_in[64]), .Y(n3020) );
  INVX1 U9027 ( .A(n2993), .Y(n2999) );
  INVX1 U9028 ( .A(n2721), .Y(n2714) );
  INVX1 U9029 ( .A(top_core_EC_ss_in[16]), .Y(n3380) );
  INVX1 U9030 ( .A(n3082), .Y(n3075) );
  INVX1 U9031 ( .A(n2783), .Y(n2779) );
  INVX1 U9032 ( .A(n3443), .Y(n3436) );
  INVX1 U9033 ( .A(top_core_EC_ss_in[48]), .Y(n3139) );
  INVX1 U9034 ( .A(top_core_EC_ss_in[88]), .Y(n2839) );
  INVX1 U9035 ( .A(n3325), .Y(n3319) );
  INVX1 U9036 ( .A(n2811), .Y(n2817) );
  INVX1 U9037 ( .A(n2880), .Y(n2887) );
  INVX1 U9038 ( .A(n2647), .Y(n2642) );
  INVX1 U9039 ( .A(n2699), .Y(n2704) );
  INVX1 U9040 ( .A(n3060), .Y(n3065) );
  INVX1 U9041 ( .A(n3429), .Y(n3424) );
  INVX1 U9042 ( .A(n2820), .Y(n2825) );
  INVX1 U9043 ( .A(n3189), .Y(n3184) );
  INVX1 U9044 ( .A(n3372), .Y(n3367) );
  INVX1 U9045 ( .A(n2587), .Y(n2582) );
  INVX1 U9046 ( .A(n2769), .Y(n2764) );
  INVX1 U9047 ( .A(n2941), .Y(n2946) );
  INVX1 U9048 ( .A(n3131), .Y(n3126) );
  INVX1 U9049 ( .A(n2903), .Y(n2897) );
  INVX1 U9050 ( .A(n3504), .Y(n3498) );
  INVX1 U9051 ( .A(n2660), .Y(n2654) );
  INVX1 U9052 ( .A(n3263), .Y(n3257) );
  INVX1 U9053 ( .A(n3202), .Y(n3196) );
  INVX1 U9054 ( .A(n2964), .Y(n2958) );
  INVX1 U9055 ( .A(n2599), .Y(n2593) );
  INVX1 U9056 ( .A(n3325), .Y(n3320) );
  INVX1 U9057 ( .A(n3016), .Y(n3021) );
  INVX1 U9058 ( .A(n2721), .Y(n2715) );
  INVX1 U9059 ( .A(n3376), .Y(n3381) );
  INVX1 U9060 ( .A(n3082), .Y(n3076) );
  INVX1 U9061 ( .A(n2783), .Y(n2780) );
  INVX1 U9062 ( .A(n3443), .Y(n3437) );
  INVX1 U9063 ( .A(n3135), .Y(n3140) );
  INVX1 U9064 ( .A(n2834), .Y(n2840) );
  INVX1 U9065 ( .A(n3503), .Y(n3499) );
  INVX1 U9066 ( .A(n2902), .Y(n2898) );
  INVX1 U9067 ( .A(n2659), .Y(n2655) );
  INVX1 U9068 ( .A(n3262), .Y(n3258) );
  INVX1 U9069 ( .A(n2720), .Y(n2716) );
  INVX1 U9070 ( .A(n3081), .Y(n3077) );
  INVX1 U9071 ( .A(n3442), .Y(n3438) );
  INVX1 U9072 ( .A(top_core_EC_ss_in[88]), .Y(n2841) );
  INVX1 U9073 ( .A(n3016), .Y(n3022) );
  INVX1 U9074 ( .A(n3201), .Y(n3197) );
  INVX1 U9075 ( .A(n3376), .Y(n3382) );
  INVX1 U9076 ( .A(n2598), .Y(n2594) );
  INVX1 U9077 ( .A(n2963), .Y(n2959) );
  INVX1 U9078 ( .A(n3135), .Y(n3141) );
  INVX1 U9079 ( .A(n3324), .Y(n3321) );
  INVX1 U9080 ( .A(n2902), .Y(n2899) );
  INVX1 U9081 ( .A(n3503), .Y(n3500) );
  INVX1 U9082 ( .A(n3262), .Y(n3259) );
  INVX1 U9083 ( .A(n2659), .Y(n2656) );
  INVX1 U9084 ( .A(n3201), .Y(n3198) );
  INVX1 U9085 ( .A(n2720), .Y(n2717) );
  INVX1 U9086 ( .A(n3081), .Y(n3078) );
  INVX1 U9087 ( .A(n2963), .Y(n2960) );
  INVX1 U9088 ( .A(n3442), .Y(n3439) );
  INVX1 U9089 ( .A(n2598), .Y(n2595) );
  INVX1 U9090 ( .A(top_core_EC_ss_in[88]), .Y(n2842) );
  INVX1 U9091 ( .A(n3324), .Y(n3322) );
  INVX1 U9092 ( .A(n2902), .Y(n2900) );
  INVX1 U9093 ( .A(n3503), .Y(n3501) );
  INVX1 U9094 ( .A(n2659), .Y(n2657) );
  INVX1 U9095 ( .A(n3262), .Y(n3260) );
  INVX1 U9096 ( .A(n3201), .Y(n3199) );
  INVX1 U9097 ( .A(n2963), .Y(n2961) );
  INVX1 U9098 ( .A(n2598), .Y(n2596) );
  INVX1 U9099 ( .A(n3324), .Y(n3323) );
  INVX1 U9100 ( .A(n2720), .Y(n2718) );
  INVX1 U9101 ( .A(n3081), .Y(n3079) );
  INVX1 U9102 ( .A(top_core_EC_ss_in[96]), .Y(n2781) );
  INVX1 U9103 ( .A(n3442), .Y(n3440) );
  INVX1 U9104 ( .A(n2844), .Y(n2843) );
  INVX1 U9105 ( .A(n3466), .Y(n3463) );
  INVX1 U9106 ( .A(n2865), .Y(n2862) );
  INVX1 U9107 ( .A(n2623), .Y(n2619) );
  INVX1 U9108 ( .A(n3225), .Y(n3222) );
  INVX1 U9109 ( .A(n3164), .Y(n3160) );
  INVX1 U9110 ( .A(n2926), .Y(n2922) );
  INVX1 U9111 ( .A(n3286), .Y(n3282) );
  INVX1 U9112 ( .A(n2987), .Y(n2983) );
  INVX1 U9113 ( .A(n2684), .Y(n2681) );
  INVX1 U9114 ( .A(n3347), .Y(n3343) );
  INVX1 U9115 ( .A(n3045), .Y(n3041) );
  INVX1 U9116 ( .A(n2744), .Y(n2741) );
  INVX1 U9117 ( .A(n3405), .Y(n3401) );
  INVX1 U9118 ( .A(n3106), .Y(n3103) );
  INVX1 U9119 ( .A(n2805), .Y(n2801) );
  INVX1 U9120 ( .A(n2222), .Y(n2228) );
  INVX1 U9121 ( .A(n2226), .Y(n2229) );
  INVX1 U9122 ( .A(n2220), .Y(n2230) );
  INVX1 U9123 ( .A(n2220), .Y(n2231) );
  INVX1 U9124 ( .A(n2220), .Y(n2232) );
  INVX1 U9125 ( .A(n2622), .Y(n2620) );
  INVX1 U9126 ( .A(n3163), .Y(n3161) );
  INVX1 U9127 ( .A(n2925), .Y(n2923) );
  INVX1 U9128 ( .A(n2550), .Y(n2558) );
  INVX1 U9129 ( .A(n3285), .Y(n3283) );
  INVX1 U9130 ( .A(n2986), .Y(n2984) );
  INVX1 U9131 ( .A(n3346), .Y(n3344) );
  INVX1 U9132 ( .A(n3044), .Y(n3042) );
  INVX1 U9133 ( .A(n3404), .Y(n3402) );
  INVX1 U9134 ( .A(n2804), .Y(n2802) );
  INVX1 U9135 ( .A(n2561), .Y(n2559) );
  INVX1 U9136 ( .A(n2349), .Y(n2351) );
  INVX1 U9137 ( .A(n2348), .Y(n2352) );
  INVX1 U9138 ( .A(n2363), .Y(n2358) );
  INVX1 U9139 ( .A(n2364), .Y(n2359) );
  INVX1 U9140 ( .A(n2364), .Y(n2353) );
  INVX1 U9141 ( .A(n2364), .Y(n2354) );
  INVX1 U9142 ( .A(n2363), .Y(n2355) );
  INVX1 U9143 ( .A(n2363), .Y(n2356) );
  INVX1 U9144 ( .A(n2364), .Y(n2362) );
  INVX1 U9145 ( .A(n2364), .Y(n2357) );
  INVX1 U9146 ( .A(n2363), .Y(n2360) );
  INVX1 U9147 ( .A(n2363), .Y(n2361) );
  INVX1 U9148 ( .A(n2661), .Y(n2658) );
  INVX1 U9149 ( .A(n2600), .Y(n2597) );
  INVX1 U9150 ( .A(n2783), .Y(n2782) );
  INVX1 U9151 ( .A(n3083), .Y(n3080) );
  INVX1 U9152 ( .A(n3249), .Y(n3245) );
  INVX1 U9153 ( .A(top_core_EC_ss_in[113]), .Y(n2643) );
  INVX1 U9154 ( .A(n2700), .Y(n2705) );
  INVX1 U9155 ( .A(n3490), .Y(n3487) );
  INVX1 U9156 ( .A(n2647), .Y(n2644) );
  INVX1 U9157 ( .A(top_core_EC_ss_in[33]), .Y(n3246) );
  INVX1 U9158 ( .A(top_core_EC_ss_in[41]), .Y(n3186) );
  INVX1 U9159 ( .A(top_core_EC_ss_in[121]), .Y(n2584) );
  INVX1 U9160 ( .A(top_core_EC_ss_in[9]), .Y(n3425) );
  INVX1 U9161 ( .A(n2724), .Y(n2719) );
  INVX1 U9162 ( .A(n3446), .Y(n3441) );
  INVX1 U9163 ( .A(top_core_EC_ss_in[25]), .Y(n3307) );
  INVX1 U9164 ( .A(top_core_EC_ss_in[65]), .Y(n3007) );
  INVX1 U9165 ( .A(top_core_EC_ss_in[65]), .Y(n3008) );
  INVX1 U9166 ( .A(n3189), .Y(n3185) );
  INVX1 U9167 ( .A(n2699), .Y(n2706) );
  INVX1 U9168 ( .A(top_core_EC_ss_in[17]), .Y(n3368) );
  INVX1 U9169 ( .A(n3372), .Y(n3369) );
  INVX1 U9170 ( .A(n2587), .Y(n2583) );
  INVX1 U9171 ( .A(n3069), .Y(n3066) );
  INVX1 U9172 ( .A(top_core_EC_ss_in[97]), .Y(n2765) );
  INVX1 U9173 ( .A(n2769), .Y(n2766) );
  INVX1 U9174 ( .A(n2950), .Y(n2947) );
  INVX1 U9175 ( .A(n3429), .Y(n3426) );
  INVX1 U9176 ( .A(top_core_EC_ss_in[49]), .Y(n3127) );
  INVX1 U9177 ( .A(n3131), .Y(n3128) );
  INVX1 U9178 ( .A(top_core_EC_ss_in[25]), .Y(n3306) );
  INVX1 U9179 ( .A(n2829), .Y(n2826) );
  INVX1 U9180 ( .A(n2879), .Y(n2878) );
  INVX1 U9181 ( .A(n2637), .Y(n2636) );
  INVX1 U9182 ( .A(n3239), .Y(n3238) );
  INVX1 U9183 ( .A(n3178), .Y(n3177) );
  INVX1 U9184 ( .A(n2576), .Y(n2575) );
  INVX1 U9185 ( .A(n2940), .Y(n2939) );
  INVX1 U9186 ( .A(n3300), .Y(n3299) );
  INVX1 U9187 ( .A(n3001), .Y(n3000) );
  INVX1 U9188 ( .A(n2698), .Y(n2697) );
  INVX1 U9189 ( .A(n3361), .Y(n3360) );
  INVX1 U9190 ( .A(n3059), .Y(n3058) );
  INVX1 U9191 ( .A(n2758), .Y(n2757) );
  INVX1 U9192 ( .A(n3419), .Y(n3418) );
  INVX1 U9193 ( .A(n3120), .Y(n3119) );
  INVX1 U9194 ( .A(n2819), .Y(n2818) );
  INVX1 U9195 ( .A(n3482), .Y(n3488) );
  INVX1 U9196 ( .A(n2906), .Y(n2901) );
  INVX1 U9197 ( .A(n2640), .Y(n2645) );
  INVX1 U9198 ( .A(n3249), .Y(n3247) );
  INVX1 U9199 ( .A(n3266), .Y(n3261) );
  INVX1 U9200 ( .A(n3205), .Y(n3200) );
  INVX1 U9201 ( .A(n2967), .Y(n2962) );
  INVX1 U9202 ( .A(n3179), .Y(n3187) );
  INVX1 U9203 ( .A(n2577), .Y(n2585) );
  INVX1 U9204 ( .A(n2950), .Y(n2948) );
  INVX1 U9205 ( .A(n3310), .Y(n3308) );
  INVX1 U9206 ( .A(n3011), .Y(n3009) );
  INVX1 U9207 ( .A(n2701), .Y(n2707) );
  INVX1 U9208 ( .A(n3362), .Y(n3370) );
  INVX1 U9209 ( .A(n3069), .Y(n3067) );
  INVX1 U9210 ( .A(n2759), .Y(n2767) );
  INVX1 U9211 ( .A(n3422), .Y(n3427) );
  INVX1 U9212 ( .A(n3121), .Y(n3129) );
  INVX1 U9213 ( .A(n2829), .Y(n2827) );
  INVX1 U9214 ( .A(n3505), .Y(n3502) );
  INVX1 U9215 ( .A(n3016), .Y(n3023) );
  INVX1 U9216 ( .A(n3376), .Y(n3383) );
  INVX1 U9217 ( .A(n3135), .Y(n3142) );
  INVX1 U9218 ( .A(n3626), .Y(n3625) );
  INVX1 U9219 ( .A(n3626), .Y(n3624) );
  INVX1 U9220 ( .A(n2220), .Y(n2234) );
  INVX1 U9221 ( .A(n2227), .Y(n2233) );
  CLKINVX2 U9222 ( .A(n274), .Y(n4176) );
  CLKINVX2 U9223 ( .A(n275), .Y(n4180) );
  CLKINVX2 U9224 ( .A(n276), .Y(n4184) );
  CLKINVX2 U9225 ( .A(n277), .Y(n4188) );
  CLKINVX2 U9226 ( .A(n282), .Y(n4177) );
  CLKINVX2 U9227 ( .A(n283), .Y(n4181) );
  CLKINVX2 U9228 ( .A(n284), .Y(n4185) );
  CLKINVX2 U9229 ( .A(n285), .Y(n4189) );
  CLKINVX2 U9230 ( .A(n267), .Y(n4178) );
  CLKINVX2 U9231 ( .A(n268), .Y(n4182) );
  CLKINVX2 U9232 ( .A(n269), .Y(n4186) );
  CLKINVX2 U9233 ( .A(n270), .Y(n4190) );
  CLKINVX2 U9234 ( .A(n47), .Y(n4179) );
  CLKINVX2 U9235 ( .A(n48), .Y(n4183) );
  CLKINVX2 U9236 ( .A(n49), .Y(n4187) );
  CLKINVX2 U9237 ( .A(n87), .Y(n4191) );
  CLKINVX2 U9238 ( .A(n278), .Y(n4145) );
  CLKINVX2 U9239 ( .A(n279), .Y(n4149) );
  CLKINVX2 U9240 ( .A(n280), .Y(n4153) );
  CLKINVX2 U9241 ( .A(n281), .Y(n4157) );
  CLKINVX2 U9242 ( .A(n286), .Y(n4146) );
  CLKINVX2 U9243 ( .A(n287), .Y(n4150) );
  CLKINVX2 U9244 ( .A(n288), .Y(n4154) );
  CLKINVX2 U9245 ( .A(n289), .Y(n4158) );
  CLKINVX2 U9246 ( .A(n271), .Y(n4147) );
  CLKINVX2 U9247 ( .A(n84), .Y(n4151) );
  CLKINVX2 U9248 ( .A(n272), .Y(n4155) );
  CLKINVX2 U9249 ( .A(n273), .Y(n4159) );
  CLKINVX2 U9250 ( .A(n7), .Y(n4148) );
  CLKINVX2 U9251 ( .A(n9), .Y(n4152) );
  CLKINVX2 U9252 ( .A(n10), .Y(n4156) );
  CLKINVX2 U9253 ( .A(n11), .Y(n4160) );
  CLKINVX2 U9254 ( .A(n294), .Y(n4161) );
  CLKINVX2 U9255 ( .A(n295), .Y(n4165) );
  CLKINVX2 U9256 ( .A(n296), .Y(n4168) );
  CLKINVX2 U9257 ( .A(n297), .Y(n4172) );
  CLKINVX2 U9258 ( .A(n298), .Y(n4162) );
  CLKINVX2 U9259 ( .A(n299), .Y(n4166) );
  CLKINVX2 U9260 ( .A(n300), .Y(n4169) );
  CLKINVX2 U9261 ( .A(n301), .Y(n4173) );
  CLKINVX2 U9262 ( .A(n290), .Y(n4163) );
  CLKINVX2 U9263 ( .A(n291), .Y(n4167) );
  CLKINVX2 U9264 ( .A(n292), .Y(n4170) );
  CLKINVX2 U9265 ( .A(n293), .Y(n4174) );
  CLKINVX2 U9266 ( .A(n8), .Y(n4164) );
  CLKINVX2 U9267 ( .A(n12), .Y(n4171) );
  CLKINVX2 U9268 ( .A(n88), .Y(n4175) );
  NAND2X2 U9269 ( .A(n6550), .B(n1674), .Y(n13293) );
  NAND2X2 U9270 ( .A(n6845), .B(n1732), .Y(n12663) );
  NAND2X2 U9271 ( .A(n6891), .B(n1703), .Y(n12978) );
  NAND2X2 U9272 ( .A(n5388), .B(n2867), .Y(n9944) );
  NAND2X2 U9273 ( .A(n6175), .B(n3468), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n129) );
  NAND2X2 U9274 ( .A(n5034), .B(n2625), .Y(n11112) );
  NAND2X2 U9275 ( .A(n5860), .B(n3227), .Y(n8192) );
  NAND2X2 U9276 ( .A(n5118), .B(n2686), .Y(n10820) );
  NAND2X2 U9277 ( .A(n5624), .B(n3047), .Y(n9068) );
  NAND2X2 U9278 ( .A(n6088), .B(n3407), .Y(n7316) );
  NAND2X2 U9279 ( .A(n5304), .B(n2807), .Y(n10236) );
  NAND2X2 U9280 ( .A(n5548), .B(n2989), .Y(n9360) );
  NAND2X2 U9281 ( .A(n5776), .B(n3166), .Y(n8484) );
  NAND2X2 U9282 ( .A(n6012), .B(n3349), .Y(n7608) );
  NAND2X2 U9283 ( .A(n4918), .B(n2564), .Y(n11404) );
  NAND2X2 U9284 ( .A(n5226), .B(n2746), .Y(n10528) );
  NAND2X2 U9285 ( .A(n5472), .B(n2928), .Y(n9652) );
  NAND2X2 U9286 ( .A(n5700), .B(n3108), .Y(n8776) );
  NAND2X2 U9287 ( .A(n5936), .B(n3288), .Y(n7900) );
  NAND2X2 U9288 ( .A(n5388), .B(n2868), .Y(n9887) );
  NAND2X2 U9289 ( .A(n6175), .B(n3471), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n69) );
  NAND2X2 U9290 ( .A(n5034), .B(n2626), .Y(n11055) );
  NAND2X2 U9291 ( .A(n5860), .B(n3228), .Y(n8135) );
  NAND2X2 U9292 ( .A(n5118), .B(n2688), .Y(n10763) );
  NAND2X2 U9293 ( .A(n5624), .B(n3049), .Y(n9011) );
  NAND2X2 U9294 ( .A(n6088), .B(n3409), .Y(n7259) );
  NAND2X2 U9295 ( .A(n5304), .B(n2808), .Y(n10179) );
  NAND2X2 U9296 ( .A(n5548), .B(n2990), .Y(n9303) );
  NAND2X2 U9297 ( .A(n5776), .B(n3167), .Y(n8427) );
  NAND2X2 U9298 ( .A(n6012), .B(n3350), .Y(n7551) );
  NAND2X2 U9299 ( .A(n4918), .B(n2565), .Y(n11347) );
  NAND2X2 U9300 ( .A(n5226), .B(n2747), .Y(n10471) );
  NAND2X2 U9301 ( .A(n5472), .B(n2929), .Y(n9595) );
  NAND2X2 U9302 ( .A(n5700), .B(n3109), .Y(n8719) );
  NAND2X2 U9303 ( .A(n5936), .B(n3289), .Y(n7843) );
  NAND2X2 U9304 ( .A(n5387), .B(n2869), .Y(n9943) );
  NAND2X2 U9305 ( .A(n6174), .B(n3470), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n128) );
  NAND2X2 U9306 ( .A(n5033), .B(n2627), .Y(n11111) );
  NAND2X2 U9307 ( .A(n5859), .B(n3229), .Y(n8191) );
  NAND2X2 U9308 ( .A(n5117), .B(n2687), .Y(n10819) );
  NAND2X2 U9309 ( .A(n6087), .B(n3408), .Y(n7315) );
  NAND2X2 U9310 ( .A(n5623), .B(n3048), .Y(n9067) );
  NAND2X2 U9311 ( .A(n5303), .B(n2809), .Y(n10235) );
  NAND2X2 U9312 ( .A(n5547), .B(n2991), .Y(n9359) );
  NAND2X2 U9313 ( .A(n5775), .B(n3168), .Y(n8483) );
  NAND2X2 U9314 ( .A(n6011), .B(n3351), .Y(n7607) );
  NAND2X2 U9315 ( .A(n4917), .B(n2566), .Y(n11403) );
  NAND2X2 U9316 ( .A(n5225), .B(n2748), .Y(n10527) );
  NAND2X2 U9317 ( .A(n5471), .B(n2930), .Y(n9651) );
  NAND2X2 U9318 ( .A(n5699), .B(n3110), .Y(n8775) );
  NAND2X2 U9319 ( .A(n5935), .B(n3290), .Y(n7899) );
  NAND2X2 U9320 ( .A(n995), .B(n2872), .Y(n17208) );
  NAND2X2 U9321 ( .A(n1134), .B(n3473), .Y(n14058) );
  NAND2X2 U9322 ( .A(n1079), .B(n3232), .Y(n15318) );
  NAND2X2 U9323 ( .A(n939), .B(n2630), .Y(n18468) );
  NAND2X2 U9324 ( .A(n1065), .B(n3171), .Y(n15633) );
  NAND2X2 U9325 ( .A(n1009), .B(n2933), .Y(n16893) );
  NAND2X2 U9326 ( .A(n925), .B(n2569), .Y(n18783) );
  NAND2X2 U9327 ( .A(n1093), .B(n3293), .Y(n15003) );
  NAND2X2 U9328 ( .A(n1023), .B(n2994), .Y(n16578) );
  NAND2X2 U9329 ( .A(n953), .B(n2691), .Y(n18153) );
  NAND2X2 U9330 ( .A(n1107), .B(n3354), .Y(n14688) );
  NAND2X2 U9331 ( .A(n1037), .B(n3052), .Y(n16263) );
  NAND2X2 U9332 ( .A(n967), .B(n2751), .Y(n17838) );
  NAND2X2 U9333 ( .A(n1121), .B(n3412), .Y(n14373) );
  NAND2X2 U9334 ( .A(n1051), .B(n3113), .Y(n15948) );
  NAND2X2 U9335 ( .A(n981), .B(n2812), .Y(n17523) );
  XOR2X1 U9336 ( .A(n1542), .B(top_core_EC_mix_in[40]), .Y(
        top_core_EC_mc_mix_in_4_42_) );
  XOR2X1 U9337 ( .A(n1542), .B(top_core_EC_mix_in[43]), .Y(
        top_core_EC_mc_mix_in_8[46]) );
  NAND2X1 U9338 ( .A(n685), .B(n1160), .Y(n13699) );
  NOR2X1 U9339 ( .A(n11852), .B(n1259), .Y(n11741) );
  NOR2X1 U9340 ( .A(top_core_KE_sb1_n281), .B(n1331), .Y(top_core_KE_sb1_n168)
         );
  NOR2X1 U9341 ( .A(n13428), .B(n1275), .Y(n13318) );
  NOR2X1 U9342 ( .A(n12168), .B(n1262), .Y(n12057) );
  NOR2X1 U9343 ( .A(n12798), .B(n1269), .Y(n12688) );
  NOR2X1 U9344 ( .A(n13113), .B(n1272), .Y(n13003) );
  NOR2X1 U9345 ( .A(n13743), .B(n1278), .Y(n13633) );
  NOR2X1 U9346 ( .A(n13282), .B(n180), .Y(n13258) );
  NOR2X1 U9347 ( .A(n12967), .B(n182), .Y(n12943) );
  NOR2X1 U9348 ( .A(n12652), .B(n181), .Y(n12628) );
  NOR2X1 U9349 ( .A(n3), .B(n686), .Y(n13241) );
  NOR2X1 U9350 ( .A(n4), .B(n688), .Y(n12611) );
  NOR2X1 U9351 ( .A(n5), .B(n687), .Y(n12926) );
  NAND2X1 U9352 ( .A(n999), .B(n2872), .Y(n17062) );
  NAND2X1 U9353 ( .A(n1138), .B(n3473), .Y(n13912) );
  NAND2X1 U9354 ( .A(n943), .B(n2630), .Y(n18322) );
  NAND2X1 U9355 ( .A(n1083), .B(n3232), .Y(n15172) );
  NAND2X1 U9356 ( .A(n1069), .B(n3171), .Y(n15487) );
  NAND2X1 U9357 ( .A(n929), .B(n2569), .Y(n18637) );
  NAND2X1 U9358 ( .A(n1013), .B(n2933), .Y(n16747) );
  NAND2X1 U9359 ( .A(n1097), .B(n3293), .Y(n14857) );
  NAND2X1 U9360 ( .A(n1027), .B(n2994), .Y(n16432) );
  NAND2X1 U9361 ( .A(n957), .B(n2691), .Y(n18007) );
  NAND2X1 U9362 ( .A(n1111), .B(n3354), .Y(n14542) );
  NAND2X1 U9363 ( .A(n1041), .B(n3052), .Y(n16117) );
  NAND2X1 U9364 ( .A(n971), .B(n2751), .Y(n17692) );
  NAND2X1 U9365 ( .A(n1125), .B(n3412), .Y(n14227) );
  NAND2X1 U9366 ( .A(n1055), .B(n3113), .Y(n15802) );
  NAND2X1 U9367 ( .A(n985), .B(n2812), .Y(n17377) );
  NOR3XL U9368 ( .A(n13885), .B(n1144), .C(n107), .Y(n13859) );
  NOR3XL U9369 ( .A(n17035), .B(n1005), .C(n106), .Y(n17009) );
  NOR3XL U9370 ( .A(n18295), .B(n949), .C(n108), .Y(n18269) );
  NOR3XL U9371 ( .A(n15145), .B(n1089), .C(n109), .Y(n15119) );
  NOR3XL U9372 ( .A(n15460), .B(n1075), .C(n110), .Y(n15434) );
  NOR3XL U9373 ( .A(n18610), .B(n935), .C(n111), .Y(n18584) );
  NOR3XL U9374 ( .A(n16720), .B(n1019), .C(n112), .Y(n16694) );
  NOR3XL U9375 ( .A(n14830), .B(n1103), .C(n113), .Y(n14804) );
  NOR3XL U9376 ( .A(n16405), .B(n1033), .C(n114), .Y(n16379) );
  NOR3XL U9377 ( .A(n17980), .B(n963), .C(n115), .Y(n17954) );
  NOR3XL U9378 ( .A(n14515), .B(n1117), .C(n116), .Y(n14489) );
  NOR3XL U9379 ( .A(n16090), .B(n1047), .C(n117), .Y(n16064) );
  NOR3XL U9380 ( .A(n17665), .B(n977), .C(n118), .Y(n17639) );
  NOR3XL U9381 ( .A(n14200), .B(n1131), .C(n119), .Y(n14174) );
  NOR3XL U9382 ( .A(n15775), .B(n1061), .C(n120), .Y(n15749) );
  NOR3XL U9383 ( .A(n17350), .B(n991), .C(n121), .Y(n17324) );
  OAI222XL U9384 ( .A0(n2859), .A1(n17148), .B0(n17149), .B1(n17030), .C0(
        n17150), .C1(n2852), .Y(n17147) );
  AOI211X1 U9385 ( .A0(n370), .A1(n2870), .B0(n17154), .C0(n995), .Y(n17149)
         );
  NOR4BX1 U9386 ( .AN(n17151), .B(n17058), .C(n17152), .D(n5376), .Y(n17150)
         );
  OAI222XL U9387 ( .A0(n3460), .A1(n13998), .B0(n13999), .B1(n13880), .C0(
        n14000), .C1(n3453), .Y(n13997) );
  AOI211X1 U9388 ( .A0(n369), .A1(n3471), .B0(n14004), .C0(n1134), .Y(n13999)
         );
  NOR4BX1 U9389 ( .AN(n14001), .B(n13908), .C(n14002), .D(n6166), .Y(n14000)
         );
  OAI222XL U9390 ( .A0(n2617), .A1(n18408), .B0(n18409), .B1(n18290), .C0(
        n18410), .C1(n2610), .Y(n18407) );
  AOI211X1 U9391 ( .A0(n371), .A1(n2628), .B0(n18414), .C0(n939), .Y(n18409)
         );
  NOR4BX1 U9392 ( .AN(n18411), .B(n18318), .C(n18412), .D(n5022), .Y(n18410)
         );
  OAI222XL U9393 ( .A0(n3219), .A1(n15258), .B0(n15259), .B1(n15140), .C0(
        n15260), .C1(n3212), .Y(n15257) );
  AOI211X1 U9394 ( .A0(n372), .A1(n3230), .B0(n15264), .C0(n1079), .Y(n15259)
         );
  NOR4BX1 U9395 ( .AN(n15261), .B(n15168), .C(n15262), .D(n5848), .Y(n15260)
         );
  OAI222XL U9396 ( .A0(n3158), .A1(n15573), .B0(n15574), .B1(n15455), .C0(
        n15575), .C1(n3151), .Y(n15572) );
  AOI211X1 U9397 ( .A0(n373), .A1(n3169), .B0(n15579), .C0(n1065), .Y(n15574)
         );
  NOR4BX1 U9398 ( .AN(n15576), .B(n15483), .C(n15577), .D(n5764), .Y(n15575)
         );
  OAI222XL U9399 ( .A0(n2556), .A1(n18723), .B0(n18724), .B1(n18605), .C0(
        n18725), .C1(n2549), .Y(n18722) );
  AOI211X1 U9400 ( .A0(n374), .A1(n2567), .B0(n18729), .C0(n925), .Y(n18724)
         );
  NOR4BX1 U9401 ( .AN(n18726), .B(n18633), .C(n18727), .D(n4906), .Y(n18725)
         );
  OAI222XL U9402 ( .A0(n2920), .A1(n16833), .B0(n16834), .B1(n16715), .C0(
        n16835), .C1(n2913), .Y(n16832) );
  AOI211X1 U9403 ( .A0(n375), .A1(n2931), .B0(n16839), .C0(n1009), .Y(n16834)
         );
  NOR4BX1 U9404 ( .AN(n16836), .B(n16743), .C(n16837), .D(n5460), .Y(n16835)
         );
  OAI222XL U9405 ( .A0(n3280), .A1(n14943), .B0(n14944), .B1(n14825), .C0(
        n14945), .C1(n3273), .Y(n14942) );
  AOI211X1 U9406 ( .A0(n376), .A1(n3291), .B0(n14949), .C0(n1093), .Y(n14944)
         );
  NOR4BX1 U9407 ( .AN(n14946), .B(n14853), .C(n14947), .D(n5924), .Y(n14945)
         );
  OAI222XL U9408 ( .A0(n2981), .A1(n16518), .B0(n16519), .B1(n16400), .C0(
        n16520), .C1(n2974), .Y(n16517) );
  AOI211X1 U9409 ( .A0(n377), .A1(n2992), .B0(n16524), .C0(n1023), .Y(n16519)
         );
  NOR4BX1 U9410 ( .AN(n16521), .B(n16428), .C(n16522), .D(n5536), .Y(n16520)
         );
  OAI222XL U9411 ( .A0(n2678), .A1(n18093), .B0(n18094), .B1(n17975), .C0(
        n18095), .C1(n2671), .Y(n18092) );
  AOI211X1 U9412 ( .A0(n378), .A1(n2689), .B0(n18099), .C0(n953), .Y(n18094)
         );
  NOR4BX1 U9413 ( .AN(n18096), .B(n18003), .C(n18097), .D(n5106), .Y(n18095)
         );
  OAI222XL U9414 ( .A0(n3341), .A1(n14628), .B0(n14629), .B1(n14510), .C0(
        n14630), .C1(n3334), .Y(n14627) );
  AOI211X1 U9415 ( .A0(n379), .A1(n3352), .B0(n14634), .C0(n1107), .Y(n14629)
         );
  NOR4BX1 U9416 ( .AN(n14631), .B(n14538), .C(n14632), .D(n6000), .Y(n14630)
         );
  OAI222XL U9417 ( .A0(n3039), .A1(n16203), .B0(n16204), .B1(n16085), .C0(
        n16205), .C1(n3032), .Y(n16202) );
  AOI211X1 U9418 ( .A0(n380), .A1(n3050), .B0(n16209), .C0(n1037), .Y(n16204)
         );
  NOR4BX1 U9419 ( .AN(n16206), .B(n16113), .C(n16207), .D(n5612), .Y(n16205)
         );
  OAI222XL U9420 ( .A0(n2738), .A1(n17778), .B0(n17779), .B1(n17660), .C0(
        n17780), .C1(n2731), .Y(n17777) );
  AOI211X1 U9421 ( .A0(n381), .A1(n2747), .B0(n17784), .C0(n967), .Y(n17779)
         );
  NOR4BX1 U9422 ( .AN(n17781), .B(n17688), .C(n17782), .D(n5214), .Y(n17780)
         );
  OAI222XL U9423 ( .A0(n3399), .A1(n14313), .B0(n14314), .B1(n14195), .C0(
        n14315), .C1(n3392), .Y(n14312) );
  AOI211X1 U9424 ( .A0(n382), .A1(n3410), .B0(n14319), .C0(n1121), .Y(n14314)
         );
  NOR4BX1 U9425 ( .AN(n14316), .B(n14223), .C(n14317), .D(n6076), .Y(n14315)
         );
  OAI222XL U9426 ( .A0(n3100), .A1(n15888), .B0(n15889), .B1(n15770), .C0(
        n15890), .C1(n3093), .Y(n15887) );
  AOI211X1 U9427 ( .A0(n383), .A1(n3111), .B0(n15894), .C0(n1051), .Y(n15889)
         );
  NOR4BX1 U9428 ( .AN(n15891), .B(n15798), .C(n15892), .D(n5688), .Y(n15890)
         );
  OAI222XL U9429 ( .A0(n2799), .A1(n17463), .B0(n17464), .B1(n17345), .C0(
        n17465), .C1(n2792), .Y(n17462) );
  AOI211X1 U9430 ( .A0(n384), .A1(n2810), .B0(n17469), .C0(n981), .Y(n17464)
         );
  NOR4BX1 U9431 ( .AN(n17466), .B(n17373), .C(n17467), .D(n5292), .Y(n17465)
         );
  OAI222XL U9432 ( .A0(n1142), .A1(n13883), .B0(n13884), .B1(n3454), .C0(
        n13885), .C1(n13886), .Y(n13871) );
  OAI222XL U9433 ( .A0(n1003), .A1(n17033), .B0(n17034), .B1(n2853), .C0(
        n17035), .C1(n17036), .Y(n17021) );
  OAI222XL U9434 ( .A0(n947), .A1(n18293), .B0(n18294), .B1(n2611), .C0(n18295), .C1(n18296), .Y(n18281) );
  OAI222XL U9435 ( .A0(n1087), .A1(n15143), .B0(n15144), .B1(n3213), .C0(
        n15145), .C1(n15146), .Y(n15131) );
  OAI222XL U9436 ( .A0(n1073), .A1(n15458), .B0(n15459), .B1(n3152), .C0(
        n15460), .C1(n15461), .Y(n15446) );
  OAI222XL U9437 ( .A0(n933), .A1(n18608), .B0(n18609), .B1(n2550), .C0(n18610), .C1(n18611), .Y(n18596) );
  OAI222XL U9438 ( .A0(n1017), .A1(n16718), .B0(n16719), .B1(n2914), .C0(
        n16720), .C1(n16721), .Y(n16706) );
  OAI222XL U9439 ( .A0(n1101), .A1(n14828), .B0(n14829), .B1(n3274), .C0(
        n14830), .C1(n14831), .Y(n14816) );
  OAI222XL U9440 ( .A0(n1031), .A1(n16403), .B0(n16404), .B1(n2975), .C0(
        n16405), .C1(n16406), .Y(n16391) );
  OAI222XL U9441 ( .A0(n961), .A1(n17978), .B0(n17979), .B1(n2672), .C0(n17980), .C1(n17981), .Y(n17966) );
  OAI222XL U9442 ( .A0(n1115), .A1(n14513), .B0(n14514), .B1(n3335), .C0(
        n14515), .C1(n14516), .Y(n14501) );
  OAI222XL U9443 ( .A0(n1045), .A1(n16088), .B0(n16089), .B1(n3033), .C0(
        n16090), .C1(n16091), .Y(n16076) );
  OAI222XL U9444 ( .A0(n975), .A1(n17663), .B0(n17664), .B1(n2732), .C0(n17665), .C1(n17666), .Y(n17651) );
  OAI222XL U9445 ( .A0(n1129), .A1(n14198), .B0(n14199), .B1(n3393), .C0(
        n14200), .C1(n14201), .Y(n14186) );
  OAI222XL U9446 ( .A0(n1059), .A1(n15773), .B0(n15774), .B1(n3094), .C0(
        n15775), .C1(n15776), .Y(n15761) );
  OAI222XL U9447 ( .A0(n989), .A1(n17348), .B0(n17349), .B1(n2793), .C0(n17350), .C1(n17351), .Y(n17336) );
  NOR2X1 U9448 ( .A(n17030), .B(n17135), .Y(n17195) );
  NOR2X1 U9449 ( .A(n13880), .B(n13985), .Y(n14045) );
  NOR2X1 U9450 ( .A(n15140), .B(n15245), .Y(n15305) );
  NOR2X1 U9451 ( .A(n18290), .B(n18395), .Y(n18455) );
  NOR2X1 U9452 ( .A(n15455), .B(n15560), .Y(n15620) );
  NOR2X1 U9453 ( .A(n16715), .B(n16820), .Y(n16880) );
  NOR2X1 U9454 ( .A(n18605), .B(n18710), .Y(n18770) );
  NOR2X1 U9455 ( .A(n14825), .B(n14930), .Y(n14990) );
  NOR2X1 U9456 ( .A(n16400), .B(n16505), .Y(n16565) );
  NOR2X1 U9457 ( .A(n17975), .B(n18080), .Y(n18140) );
  NOR2X1 U9458 ( .A(n14510), .B(n14615), .Y(n14675) );
  NOR2X1 U9459 ( .A(n16085), .B(n16190), .Y(n16250) );
  NOR2X1 U9460 ( .A(n17660), .B(n17765), .Y(n17825) );
  NOR2X1 U9461 ( .A(n14195), .B(n14300), .Y(n14360) );
  NOR2X1 U9462 ( .A(n15770), .B(n15875), .Y(n15935) );
  NOR2X1 U9463 ( .A(n17345), .B(n17450), .Y(n17510) );
  NOR2X1 U9464 ( .A(n686), .B(n1673), .Y(n13286) );
  NOR2X1 U9465 ( .A(n688), .B(n1731), .Y(n12656) );
  NOR2X1 U9466 ( .A(n687), .B(n1702), .Y(n12971) );
  AOI22X1 U9467 ( .A0(n3481), .A1(n3477), .B0(n3472), .B1(n530), .Y(n13943) );
  XOR2X1 U9468 ( .A(n1542), .B(top_core_EC_mix_in[42]), .Y(
        top_core_EC_mc_mix_in_2_43_) );
  XOR2X1 U9469 ( .A(n1548), .B(top_core_EC_mix_in[10]), .Y(
        top_core_EC_mc_mix_in_2_11_) );
  NOR3XL U9470 ( .A(n17092), .B(n2855), .C(n106), .Y(n17189) );
  NOR3XL U9471 ( .A(n13942), .B(n3463), .C(n107), .Y(n14039) );
  NOR3XL U9472 ( .A(n18352), .B(n2613), .C(n108), .Y(n18449) );
  NOR3XL U9473 ( .A(n15202), .B(n3215), .C(n109), .Y(n15299) );
  NOR3XL U9474 ( .A(n15517), .B(n3154), .C(n110), .Y(n15614) );
  NOR3XL U9475 ( .A(n16777), .B(n2916), .C(n112), .Y(n16874) );
  NOR3XL U9476 ( .A(n18667), .B(n2552), .C(n111), .Y(n18764) );
  NOR3XL U9477 ( .A(n14887), .B(n3276), .C(n113), .Y(n14984) );
  NOR3XL U9478 ( .A(n16462), .B(n2977), .C(n114), .Y(n16559) );
  NOR3XL U9479 ( .A(n18037), .B(n2674), .C(n115), .Y(n18134) );
  NOR3XL U9480 ( .A(n14572), .B(n3337), .C(n116), .Y(n14669) );
  NOR3XL U9481 ( .A(n16147), .B(n3035), .C(n117), .Y(n16244) );
  NOR3XL U9482 ( .A(n17722), .B(n2734), .C(n118), .Y(n17819) );
  NOR3XL U9483 ( .A(n14257), .B(n3395), .C(n119), .Y(n14354) );
  NOR3XL U9484 ( .A(n15832), .B(n3096), .C(n120), .Y(n15929) );
  NOR3XL U9485 ( .A(n17407), .B(n2795), .C(n121), .Y(n17504) );
  NOR2X1 U9486 ( .A(n1161), .B(n6592), .Y(n13758) );
  NAND2X1 U9487 ( .A(n6626), .B(n607), .Y(n12418) );
  OAI222XL U9488 ( .A0(n17168), .A1(n2852), .B0(n17169), .B1(n17035), .C0(
        n2859), .C1(n17170), .Y(n17157) );
  AOI211X1 U9489 ( .A0(n5357), .A1(n2884), .B0(n17171), .C0(n17172), .Y(n17170) );
  AOI221X1 U9490 ( .A0(n5376), .A1(n498), .B0(n1002), .B1(n999), .C0(n17174), 
        .Y(n17168) );
  OAI222XL U9491 ( .A0(n14018), .A1(n3453), .B0(n14019), .B1(n13885), .C0(
        n3461), .C1(n14020), .Y(n14007) );
  AOI211X1 U9492 ( .A0(n6125), .A1(n3488), .B0(n14021), .C0(n14022), .Y(n14020) );
  AOI221X1 U9493 ( .A0(n6166), .A1(n497), .B0(n1141), .B1(n1138), .C0(n14024), 
        .Y(n14018) );
  OAI222XL U9494 ( .A0(n18428), .A1(n2610), .B0(n18429), .B1(n18295), .C0(
        n2617), .C1(n18430), .Y(n18417) );
  AOI211X1 U9495 ( .A0(n5003), .A1(n2645), .B0(n18431), .C0(n18432), .Y(n18430) );
  AOI221X1 U9496 ( .A0(n5022), .A1(n501), .B0(n946), .B1(n943), .C0(n18434), 
        .Y(n18428) );
  OAI222XL U9497 ( .A0(n15278), .A1(n3212), .B0(n15279), .B1(n15145), .C0(
        n3219), .C1(n15280), .Y(n15267) );
  AOI211X1 U9498 ( .A0(n5829), .A1(n3247), .B0(n15281), .C0(n15282), .Y(n15280) );
  AOI221X1 U9499 ( .A0(n5848), .A1(n500), .B0(n1086), .B1(n1083), .C0(n15284), 
        .Y(n15278) );
  OAI222XL U9500 ( .A0(n15593), .A1(n3151), .B0(n15594), .B1(n15460), .C0(
        n3158), .C1(n15595), .Y(n15582) );
  AOI211X1 U9501 ( .A0(n5745), .A1(n3187), .B0(n15596), .C0(n15597), .Y(n15595) );
  AOI221X1 U9502 ( .A0(n5764), .A1(n499), .B0(n1072), .B1(n1069), .C0(n15599), 
        .Y(n15593) );
  OAI222XL U9503 ( .A0(n18743), .A1(n2549), .B0(n18744), .B1(n18610), .C0(
        n2556), .C1(n18745), .Y(n18732) );
  AOI211X1 U9504 ( .A0(n4887), .A1(n2585), .B0(n18746), .C0(n18747), .Y(n18745) );
  AOI221X1 U9505 ( .A0(n4906), .A1(n502), .B0(n932), .B1(n929), .C0(n18749), 
        .Y(n18743) );
  OAI222XL U9506 ( .A0(n16853), .A1(n2913), .B0(n16854), .B1(n16720), .C0(
        n2920), .C1(n16855), .Y(n16842) );
  AOI211X1 U9507 ( .A0(n5441), .A1(n2948), .B0(n16856), .C0(n16857), .Y(n16855) );
  AOI221X1 U9508 ( .A0(n5460), .A1(n503), .B0(n1016), .B1(n1013), .C0(n16859), 
        .Y(n16853) );
  OAI222XL U9509 ( .A0(n14963), .A1(n3273), .B0(n14964), .B1(n14830), .C0(
        n3280), .C1(n14965), .Y(n14952) );
  AOI211X1 U9510 ( .A0(n5905), .A1(n3308), .B0(n14966), .C0(n14967), .Y(n14965) );
  AOI221X1 U9511 ( .A0(n5924), .A1(n504), .B0(n1100), .B1(n1097), .C0(n14969), 
        .Y(n14963) );
  OAI222XL U9512 ( .A0(n16538), .A1(n2974), .B0(n16539), .B1(n16405), .C0(
        n2981), .C1(n16540), .Y(n16527) );
  AOI211X1 U9513 ( .A0(n5517), .A1(n3009), .B0(n16541), .C0(n16542), .Y(n16540) );
  AOI221X1 U9514 ( .A0(n5536), .A1(n505), .B0(n1030), .B1(n1027), .C0(n16544), 
        .Y(n16538) );
  OAI222XL U9515 ( .A0(n18113), .A1(n2671), .B0(n18114), .B1(n17980), .C0(
        n2678), .C1(n18115), .Y(n18102) );
  AOI211X1 U9516 ( .A0(n5087), .A1(n2707), .B0(n18116), .C0(n18117), .Y(n18115) );
  AOI221X1 U9517 ( .A0(n5106), .A1(n506), .B0(n960), .B1(n957), .C0(n18119), 
        .Y(n18113) );
  OAI222XL U9518 ( .A0(n14648), .A1(n3334), .B0(n14649), .B1(n14515), .C0(
        n3341), .C1(n14650), .Y(n14637) );
  AOI211X1 U9519 ( .A0(n5981), .A1(n3370), .B0(n14651), .C0(n14652), .Y(n14650) );
  AOI221X1 U9520 ( .A0(n6000), .A1(n507), .B0(n1114), .B1(n1111), .C0(n14654), 
        .Y(n14648) );
  OAI222XL U9521 ( .A0(n16223), .A1(n3032), .B0(n16224), .B1(n16090), .C0(
        n3039), .C1(n16225), .Y(n16212) );
  AOI211X1 U9522 ( .A0(n5593), .A1(n3067), .B0(n16226), .C0(n16227), .Y(n16225) );
  AOI221X1 U9523 ( .A0(n5612), .A1(n508), .B0(n1044), .B1(n1041), .C0(n16229), 
        .Y(n16223) );
  OAI222XL U9524 ( .A0(n17798), .A1(n2731), .B0(n17799), .B1(n17665), .C0(
        n2738), .C1(n17800), .Y(n17787) );
  AOI211X1 U9525 ( .A0(n5195), .A1(n2767), .B0(n17801), .C0(n17802), .Y(n17800) );
  AOI221X1 U9526 ( .A0(n5214), .A1(n509), .B0(n974), .B1(n971), .C0(n17804), 
        .Y(n17798) );
  OAI222XL U9527 ( .A0(n14333), .A1(n3392), .B0(n14334), .B1(n14200), .C0(
        n3399), .C1(n14335), .Y(n14322) );
  AOI211X1 U9528 ( .A0(n6057), .A1(n3427), .B0(n14336), .C0(n14337), .Y(n14335) );
  AOI221X1 U9529 ( .A0(n6076), .A1(n510), .B0(n1128), .B1(n1125), .C0(n14339), 
        .Y(n14333) );
  OAI222XL U9530 ( .A0(n15908), .A1(n3093), .B0(n15909), .B1(n15775), .C0(
        n3100), .C1(n15910), .Y(n15897) );
  AOI211X1 U9531 ( .A0(n5669), .A1(n3129), .B0(n15911), .C0(n15912), .Y(n15910) );
  AOI221X1 U9532 ( .A0(n5688), .A1(n511), .B0(n1058), .B1(n1055), .C0(n15914), 
        .Y(n15908) );
  OAI222XL U9533 ( .A0(n17483), .A1(n2792), .B0(n17484), .B1(n17350), .C0(
        n2799), .C1(n17485), .Y(n17472) );
  AOI211X1 U9534 ( .A0(n5273), .A1(n2827), .B0(n17486), .C0(n17487), .Y(n17485) );
  AOI221X1 U9535 ( .A0(n5292), .A1(n512), .B0(n988), .B1(n985), .C0(n17489), 
        .Y(n17483) );
  XOR2X1 U9536 ( .A(n1545), .B(top_core_EC_mix_in[26]), .Y(
        top_core_EC_mc_mix_in_2_27_) );
  NOR2X1 U9537 ( .A(n11658), .B(n1222), .Y(n11702) );
  NOR2X1 U9538 ( .A(top_core_KE_sb1_n83), .B(n1216), .Y(top_core_KE_sb1_n127)
         );
  NOR2X1 U9539 ( .A(n13235), .B(n1173), .Y(n13279) );
  NOR2X1 U9540 ( .A(n11974), .B(n1176), .Y(n12018) );
  NOR2X1 U9541 ( .A(n12605), .B(n1213), .Y(n12649) );
  NOR2X1 U9542 ( .A(n13550), .B(n1178), .Y(n13594) );
  NOR2X1 U9543 ( .A(n12920), .B(n1219), .Y(n12964) );
  NOR2X1 U9544 ( .A(n670), .B(n1666), .Y(n13231) );
  NOR2X1 U9545 ( .A(n672), .B(n1695), .Y(n12916) );
  NOR2X1 U9546 ( .A(n671), .B(n1724), .Y(n12601) );
  NAND2X1 U9547 ( .A(n1161), .B(n1178), .Y(n13649) );
  NOR2X1 U9548 ( .A(n1246), .B(n9946), .Y(n10019) );
  NOR2X1 U9549 ( .A(n1328), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n131), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n205) );
  NOR2X1 U9550 ( .A(n1254), .B(n11114), .Y(n11187) );
  NOR2X1 U9551 ( .A(n1234), .B(n8194), .Y(n8267) );
  NOR2X1 U9552 ( .A(n1252), .B(n10822), .Y(n10895) );
  NOR2X1 U9553 ( .A(n1228), .B(n7318), .Y(n7391) );
  NOR2X1 U9554 ( .A(n1240), .B(n9070), .Y(n9143) );
  NOR2X1 U9555 ( .A(n1248), .B(n10238), .Y(n10311) );
  NOR2X1 U9556 ( .A(n1242), .B(n9362), .Y(n9435) );
  NOR2X1 U9557 ( .A(n1236), .B(n8486), .Y(n8559) );
  NOR2X1 U9558 ( .A(n1230), .B(n7610), .Y(n7683) );
  NOR2X1 U9559 ( .A(n1256), .B(n11406), .Y(n11479) );
  NOR2X1 U9560 ( .A(n1250), .B(n10530), .Y(n10603) );
  NOR2X1 U9561 ( .A(n1244), .B(n9654), .Y(n9727) );
  NOR2X1 U9562 ( .A(n1238), .B(n8778), .Y(n8851) );
  NOR2X1 U9563 ( .A(n1232), .B(n7902), .Y(n7975) );
  OAI222XL U9564 ( .A0(n10069), .A1(n9895), .B0(n10070), .B1(n2853), .C0(n2859), .C1(n10071), .Y(n10058) );
  AOI211X1 U9565 ( .A0(n433), .A1(n9899), .B0(n10073), .C0(n9926), .Y(n10070)
         );
  NAND2X1 U9566 ( .A(n10074), .B(n9999), .Y(n10073) );
  OAI222XL U9567 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n255), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n78), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n256), .B1(n3454), .C0(n3460), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n257), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n244) );
  AOI211X1 U9568 ( .A0(n434), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n82), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n259), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n111), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n256) );
  NAND2X1 U9569 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n260), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n185), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n259) );
  OAI222XL U9570 ( .A0(n11237), .A1(n11063), .B0(n11238), .B1(n2611), .C0(
        n2617), .C1(n11239), .Y(n11226) );
  AOI211X1 U9571 ( .A0(n435), .A1(n11067), .B0(n11241), .C0(n11094), .Y(n11238) );
  NAND2X1 U9572 ( .A(n11242), .B(n11167), .Y(n11241) );
  OAI222XL U9573 ( .A0(n8317), .A1(n8143), .B0(n8318), .B1(n3213), .C0(n3219), 
        .C1(n8319), .Y(n8306) );
  AOI211X1 U9574 ( .A0(n436), .A1(n8147), .B0(n8321), .C0(n8174), .Y(n8318) );
  NAND2X1 U9575 ( .A(n8322), .B(n8247), .Y(n8321) );
  OAI222XL U9576 ( .A0(n10945), .A1(n10771), .B0(n10946), .B1(n2672), .C0(
        n2678), .C1(n10947), .Y(n10934) );
  AOI211X1 U9577 ( .A0(n442), .A1(n10775), .B0(n10949), .C0(n10802), .Y(n10946) );
  NAND2X1 U9578 ( .A(n10950), .B(n10875), .Y(n10949) );
  OAI222XL U9579 ( .A0(n7441), .A1(n7267), .B0(n7442), .B1(n3393), .C0(n3399), 
        .C1(n7443), .Y(n7430) );
  AOI211X1 U9580 ( .A0(n446), .A1(n7271), .B0(n7445), .C0(n7298), .Y(n7442) );
  NAND2X1 U9581 ( .A(n7446), .B(n7371), .Y(n7445) );
  OAI222XL U9582 ( .A0(n9193), .A1(n9019), .B0(n9194), .B1(n3033), .C0(n3039), 
        .C1(n9195), .Y(n9182) );
  AOI211X1 U9583 ( .A0(n444), .A1(n9023), .B0(n9197), .C0(n9050), .Y(n9194) );
  NAND2X1 U9584 ( .A(n9198), .B(n9123), .Y(n9197) );
  OAI222XL U9585 ( .A0(n10361), .A1(n10187), .B0(n10362), .B1(n2793), .C0(
        n2799), .C1(n10363), .Y(n10350) );
  AOI211X1 U9586 ( .A0(n448), .A1(n10191), .B0(n10365), .C0(n10218), .Y(n10362) );
  NAND2X1 U9587 ( .A(n10366), .B(n10291), .Y(n10365) );
  OAI222XL U9588 ( .A0(n9485), .A1(n9311), .B0(n9486), .B1(n2975), .C0(n2981), 
        .C1(n9487), .Y(n9474) );
  AOI211X1 U9589 ( .A0(n441), .A1(n9315), .B0(n9489), .C0(n9342), .Y(n9486) );
  NAND2X1 U9590 ( .A(n9490), .B(n9415), .Y(n9489) );
  OAI222XL U9591 ( .A0(n8609), .A1(n8435), .B0(n8610), .B1(n3152), .C0(n3158), 
        .C1(n8611), .Y(n8598) );
  AOI211X1 U9592 ( .A0(n437), .A1(n8439), .B0(n8613), .C0(n8466), .Y(n8610) );
  NAND2X1 U9593 ( .A(n8614), .B(n8539), .Y(n8613) );
  OAI222XL U9594 ( .A0(n7733), .A1(n7559), .B0(n7734), .B1(n3335), .C0(n3341), 
        .C1(n7735), .Y(n7722) );
  AOI211X1 U9595 ( .A0(n443), .A1(n7563), .B0(n7737), .C0(n7590), .Y(n7734) );
  NAND2X1 U9596 ( .A(n7738), .B(n7663), .Y(n7737) );
  OAI222XL U9597 ( .A0(n11529), .A1(n11355), .B0(n11530), .B1(n2550), .C0(
        n2556), .C1(n11531), .Y(n11518) );
  AOI211X1 U9598 ( .A0(n439), .A1(n11359), .B0(n11533), .C0(n11386), .Y(n11530) );
  NAND2X1 U9599 ( .A(n11534), .B(n11459), .Y(n11533) );
  OAI222XL U9600 ( .A0(n10653), .A1(n10479), .B0(n10654), .B1(n2732), .C0(
        n2738), .C1(n10655), .Y(n10642) );
  AOI211X1 U9601 ( .A0(n445), .A1(n10483), .B0(n10657), .C0(n10510), .Y(n10654) );
  NAND2X1 U9602 ( .A(n10658), .B(n10583), .Y(n10657) );
  OAI222XL U9603 ( .A0(n9777), .A1(n9603), .B0(n9778), .B1(n2914), .C0(n2920), 
        .C1(n9779), .Y(n9766) );
  AOI211X1 U9604 ( .A0(n438), .A1(n9607), .B0(n9781), .C0(n9634), .Y(n9778) );
  NAND2X1 U9605 ( .A(n9782), .B(n9707), .Y(n9781) );
  OAI222XL U9606 ( .A0(n8901), .A1(n8727), .B0(n8902), .B1(n3094), .C0(n3100), 
        .C1(n8903), .Y(n8890) );
  AOI211X1 U9607 ( .A0(n447), .A1(n8731), .B0(n8905), .C0(n8758), .Y(n8902) );
  NAND2X1 U9608 ( .A(n8906), .B(n8831), .Y(n8905) );
  OAI222XL U9609 ( .A0(n8025), .A1(n7851), .B0(n8026), .B1(n3274), .C0(n3280), 
        .C1(n8027), .Y(n8014) );
  AOI211X1 U9610 ( .A0(n440), .A1(n7855), .B0(n8029), .C0(n7882), .Y(n8026) );
  NAND2X1 U9611 ( .A(n8030), .B(n7955), .Y(n8029) );
  NAND2X1 U9612 ( .A(n1152), .B(n1687), .Y(n13311) );
  NAND2X1 U9613 ( .A(n1192), .B(n1745), .Y(n12681) );
  NAND2X1 U9614 ( .A(n1201), .B(n1716), .Y(n12996) );
  NAND2X1 U9615 ( .A(n1161), .B(n1658), .Y(n13626) );
  NOR2XL U9616 ( .A(n3), .B(n580), .Y(n13341) );
  NOR2XL U9617 ( .A(n4), .B(n584), .Y(n12711) );
  NOR2XL U9618 ( .A(n5), .B(n582), .Y(n13026) );
  NOR2X1 U9619 ( .A(n17205), .B(n2866), .Y(n17057) );
  NOR2X1 U9620 ( .A(n14055), .B(n3467), .Y(n13907) );
  NOR2X1 U9621 ( .A(n15315), .B(n3226), .Y(n15167) );
  NOR2X1 U9622 ( .A(n18465), .B(n2624), .Y(n18317) );
  NOR2X1 U9623 ( .A(n15630), .B(n3165), .Y(n15482) );
  NOR2X1 U9624 ( .A(n16890), .B(n2927), .Y(n16742) );
  NOR2X1 U9625 ( .A(n18780), .B(n2563), .Y(n18632) );
  NOR2X1 U9626 ( .A(n15000), .B(n3287), .Y(n14852) );
  NOR2X1 U9627 ( .A(n16575), .B(n2988), .Y(n16427) );
  NOR2X1 U9628 ( .A(n18150), .B(n2685), .Y(n18002) );
  NOR2X1 U9629 ( .A(n14685), .B(n3348), .Y(n14537) );
  NOR2X1 U9630 ( .A(n16260), .B(n3046), .Y(n16112) );
  NOR2X1 U9631 ( .A(n17835), .B(n2745), .Y(n17687) );
  NOR2X1 U9632 ( .A(n14370), .B(n3406), .Y(n14222) );
  NOR2X1 U9633 ( .A(n15945), .B(n3107), .Y(n15797) );
  NOR2X1 U9634 ( .A(n17520), .B(n2806), .Y(n17372) );
  OAI22X1 U9635 ( .A0(top_core_EC_mc_n922), .A1(n2465), .B0(n2375), .B1(
        top_core_EC_mc_n923), .Y(top_core_EC_mix_out_0_) );
  XOR2X1 U9636 ( .A(top_core_EC_mc_n924), .B(top_core_EC_mc_n925), .Y(
        top_core_EC_mc_n923) );
  XNOR2X1 U9637 ( .A(top_core_EC_mix_in[24]), .B(top_core_EC_mc_n926), .Y(
        top_core_EC_mc_n922) );
  XNOR2X1 U9638 ( .A(top_core_EC_mix_in[24]), .B(top_core_EC_mc_n101), .Y(
        top_core_EC_mc_n924) );
  OAI22X1 U9639 ( .A0(top_core_EC_mc_n652), .A1(n2415), .B0(n2378), .B1(
        top_core_EC_mc_n653), .Y(top_core_EC_mix_out_1_) );
  XOR2X1 U9640 ( .A(top_core_EC_mc_n654), .B(top_core_EC_mc_n655), .Y(
        top_core_EC_mc_n653) );
  XNOR2X1 U9641 ( .A(top_core_EC_mc_mix_in_2_26_), .B(top_core_EC_mc_n656), 
        .Y(top_core_EC_mc_n652) );
  XNOR2X1 U9642 ( .A(top_core_EC_mc_mix_in_2_26_), .B(top_core_EC_mc_n8), .Y(
        top_core_EC_mc_n654) );
  OAI22X1 U9643 ( .A0(top_core_EC_mc_n579), .A1(n2479), .B0(n2379), .B1(
        top_core_EC_mc_n580), .Y(top_core_EC_mix_out_2_) );
  XOR2X1 U9644 ( .A(top_core_EC_mc_n581), .B(top_core_EC_mc_n582), .Y(
        top_core_EC_mc_n580) );
  XNOR2X1 U9645 ( .A(top_core_EC_mix_in[26]), .B(top_core_EC_mc_n583), .Y(
        top_core_EC_mc_n579) );
  XNOR2X1 U9646 ( .A(top_core_EC_mix_in[26]), .B(top_core_EC_mc_n585), .Y(
        top_core_EC_mc_n581) );
  OAI22X1 U9647 ( .A0(top_core_EC_mc_n492), .A1(n2482), .B0(n2380), .B1(
        top_core_EC_mc_n493), .Y(top_core_EC_mix_out_3_) );
  XOR2X1 U9648 ( .A(top_core_EC_mc_n494), .B(top_core_EC_mc_n495), .Y(
        top_core_EC_mc_n493) );
  XNOR2X1 U9649 ( .A(top_core_EC_mix_in[27]), .B(top_core_EC_mc_n496), .Y(
        top_core_EC_mc_n492) );
  XNOR2X1 U9650 ( .A(top_core_EC_mix_in[27]), .B(top_core_EC_mc_n498), .Y(
        top_core_EC_mc_n494) );
  OAI22X1 U9651 ( .A0(top_core_EC_mc_n427), .A1(n2466), .B0(n2381), .B1(
        top_core_EC_mc_n428), .Y(top_core_EC_mix_out_4_) );
  XOR2X1 U9652 ( .A(top_core_EC_mc_n429), .B(top_core_EC_mc_n430), .Y(
        top_core_EC_mc_n428) );
  XNOR2X1 U9653 ( .A(top_core_EC_mc_mix_in_8[31]), .B(top_core_EC_mc_n431), 
        .Y(top_core_EC_mc_n427) );
  XNOR2X1 U9654 ( .A(top_core_EC_mc_mix_in_8[31]), .B(top_core_EC_mc_n433), 
        .Y(top_core_EC_mc_n429) );
  OAI22X1 U9655 ( .A0(top_core_EC_mc_n338), .A1(n2432), .B0(n2381), .B1(
        top_core_EC_mc_n339), .Y(top_core_EC_mix_out_5_) );
  XOR2X1 U9656 ( .A(top_core_EC_mc_n340), .B(top_core_EC_mc_n341), .Y(
        top_core_EC_mc_n339) );
  XNOR2X1 U9657 ( .A(n1547), .B(top_core_EC_mc_n342), .Y(top_core_EC_mc_n338)
         );
  XNOR2X1 U9658 ( .A(n1547), .B(top_core_EC_mc_n344), .Y(top_core_EC_mc_n340)
         );
  OAI22X1 U9659 ( .A0(top_core_EC_mc_n249), .A1(n2527), .B0(n2382), .B1(
        top_core_EC_mc_n250), .Y(top_core_EC_mix_out_6_) );
  XOR2X1 U9660 ( .A(top_core_EC_mc_n251), .B(top_core_EC_mc_n252), .Y(
        top_core_EC_mc_n250) );
  XNOR2X1 U9661 ( .A(n1546), .B(top_core_EC_mc_n253), .Y(top_core_EC_mc_n249)
         );
  XNOR2X1 U9662 ( .A(n1546), .B(top_core_EC_mc_n255), .Y(top_core_EC_mc_n251)
         );
  OAI22X1 U9663 ( .A0(top_core_EC_mc_n184), .A1(n2427), .B0(n2383), .B1(
        top_core_EC_mc_n185), .Y(top_core_EC_mix_out_7_) );
  XOR2X1 U9664 ( .A(top_core_EC_mc_n186), .B(top_core_EC_mc_n187), .Y(
        top_core_EC_mc_n185) );
  XNOR2X1 U9665 ( .A(n1545), .B(top_core_EC_mc_n188), .Y(top_core_EC_mc_n184)
         );
  XNOR2X1 U9666 ( .A(n1545), .B(top_core_EC_mc_n190), .Y(top_core_EC_mc_n186)
         );
  OAI22X1 U9667 ( .A0(top_core_EC_mc_n95), .A1(n2458), .B0(n2384), .B1(
        top_core_EC_mc_n96), .Y(top_core_EC_mix_out_8_) );
  XOR2X1 U9668 ( .A(top_core_EC_mc_n97), .B(top_core_EC_mc_n98), .Y(
        top_core_EC_mc_n96) );
  XNOR2X1 U9669 ( .A(n1548), .B(top_core_EC_mc_n99), .Y(top_core_EC_mc_n95) );
  XNOR2X1 U9670 ( .A(n1548), .B(top_core_EC_mc_n101), .Y(top_core_EC_mc_n97)
         );
  OAI22X1 U9671 ( .A0(top_core_EC_mc_n845), .A1(n2465), .B0(n2376), .B1(
        top_core_EC_mc_n846), .Y(top_core_EC_mix_out_10_) );
  XOR2X1 U9672 ( .A(top_core_EC_mc_n847), .B(top_core_EC_mc_n848), .Y(
        top_core_EC_mc_n846) );
  XNOR2X1 U9673 ( .A(top_core_EC_mc_mix_in_2_10_), .B(top_core_EC_mc_n849), 
        .Y(top_core_EC_mc_n845) );
  XNOR2X1 U9674 ( .A(top_core_EC_mc_mix_in_2_10_), .B(top_core_EC_mc_n585), 
        .Y(top_core_EC_mc_n847) );
  OAI22X1 U9675 ( .A0(top_core_EC_mc_n698), .A1(n2463), .B0(n2378), .B1(
        top_core_EC_mc_n699), .Y(top_core_EC_mix_out_13_) );
  XOR2X1 U9676 ( .A(top_core_EC_mc_n700), .B(top_core_EC_mc_n701), .Y(
        top_core_EC_mc_n699) );
  XNOR2X1 U9677 ( .A(top_core_EC_mc_mix_in_8[15]), .B(top_core_EC_mc_n702), 
        .Y(top_core_EC_mc_n698) );
  XNOR2X1 U9678 ( .A(top_core_EC_mc_mix_in_8[15]), .B(top_core_EC_mc_n344), 
        .Y(top_core_EC_mc_n700) );
  OAI22X1 U9679 ( .A0(top_core_EC_mc_n691), .A1(n2422), .B0(n2378), .B1(
        top_core_EC_mc_n692), .Y(top_core_EC_mix_out_14_) );
  XOR2X1 U9680 ( .A(top_core_EC_mc_n693), .B(top_core_EC_mc_n694), .Y(
        top_core_EC_mc_n692) );
  XNOR2X1 U9681 ( .A(n1550), .B(top_core_EC_mc_n695), .Y(top_core_EC_mc_n691)
         );
  XNOR2X1 U9682 ( .A(n1550), .B(top_core_EC_mc_n255), .Y(top_core_EC_mc_n693)
         );
  OAI22X1 U9683 ( .A0(top_core_EC_mc_n684), .A1(n2403), .B0(n2378), .B1(
        top_core_EC_mc_n685), .Y(top_core_EC_mix_out_15_) );
  XOR2X1 U9684 ( .A(top_core_EC_mc_n686), .B(top_core_EC_mc_n687), .Y(
        top_core_EC_mc_n685) );
  XNOR2X1 U9685 ( .A(n1549), .B(top_core_EC_mc_n688), .Y(top_core_EC_mc_n684)
         );
  XNOR2X1 U9686 ( .A(n1549), .B(top_core_EC_mc_n190), .Y(top_core_EC_mc_n686)
         );
  OAI22X1 U9687 ( .A0(top_core_EC_mc_n678), .A1(n2404), .B0(n2378), .B1(
        top_core_EC_mc_n679), .Y(top_core_EC_mix_out_16_) );
  XOR2X1 U9688 ( .A(top_core_EC_mc_n624), .B(top_core_EC_mc_n680), .Y(
        top_core_EC_mc_n679) );
  XNOR2X1 U9689 ( .A(n1545), .B(top_core_EC_mc_n681), .Y(top_core_EC_mc_n678)
         );
  XOR2X1 U9690 ( .A(top_core_EC_mc_n681), .B(top_core_EC_mc_n682), .Y(
        top_core_EC_mc_n680) );
  OAI22X1 U9691 ( .A0(top_core_EC_mc_n665), .A1(n2470), .B0(n2378), .B1(
        top_core_EC_mc_n666), .Y(top_core_EC_mix_out_18_) );
  XOR2X1 U9692 ( .A(top_core_EC_mc_n611), .B(top_core_EC_mc_n667), .Y(
        top_core_EC_mc_n666) );
  XNOR2X1 U9693 ( .A(top_core_EC_mc_mix_in_2_26_), .B(top_core_EC_mc_n668), 
        .Y(top_core_EC_mc_n665) );
  XOR2X1 U9694 ( .A(top_core_EC_mc_n584), .B(top_core_EC_mc_n668), .Y(
        top_core_EC_mc_n667) );
  OAI22X1 U9695 ( .A0(top_core_EC_mc_n640), .A1(n2416), .B0(n2378), .B1(
        top_core_EC_mc_n641), .Y(top_core_EC_mix_out_21_) );
  XOR2X1 U9696 ( .A(top_core_EC_mc_n590), .B(top_core_EC_mc_n642), .Y(
        top_core_EC_mc_n641) );
  XNOR2X1 U9697 ( .A(top_core_EC_mc_mix_in_8[31]), .B(top_core_EC_mc_n643), 
        .Y(top_core_EC_mc_n640) );
  XOR2X1 U9698 ( .A(top_core_EC_mc_n343), .B(top_core_EC_mc_n643), .Y(
        top_core_EC_mc_n642) );
  OAI22X1 U9699 ( .A0(top_core_EC_mc_n634), .A1(n2438), .B0(n2378), .B1(
        top_core_EC_mc_n635), .Y(top_core_EC_mix_out_22_) );
  XOR2X1 U9700 ( .A(top_core_EC_mc_n574), .B(top_core_EC_mc_n636), .Y(
        top_core_EC_mc_n635) );
  XNOR2X1 U9701 ( .A(n1547), .B(top_core_EC_mc_n637), .Y(top_core_EC_mc_n634)
         );
  XOR2X1 U9702 ( .A(top_core_EC_mc_n254), .B(top_core_EC_mc_n637), .Y(
        top_core_EC_mc_n636) );
  OAI22X1 U9703 ( .A0(top_core_EC_mc_n628), .A1(n2476), .B0(n2378), .B1(
        top_core_EC_mc_n629), .Y(top_core_EC_mix_out_23_) );
  XOR2X1 U9704 ( .A(top_core_EC_mc_n567), .B(top_core_EC_mc_n630), .Y(
        top_core_EC_mc_n629) );
  XNOR2X1 U9705 ( .A(n1546), .B(top_core_EC_mc_n631), .Y(top_core_EC_mc_n628)
         );
  XOR2X1 U9706 ( .A(top_core_EC_mc_n189), .B(top_core_EC_mc_n631), .Y(
        top_core_EC_mc_n630) );
  OAI22X1 U9707 ( .A0(top_core_EC_mc_n622), .A1(n2477), .B0(n2378), .B1(
        top_core_EC_mc_n623), .Y(top_core_EC_mix_out_24_) );
  XOR2X1 U9708 ( .A(top_core_EC_mc_n624), .B(top_core_EC_mc_n625), .Y(
        top_core_EC_mc_n623) );
  XNOR2X1 U9709 ( .A(n1545), .B(top_core_EC_mc_n626), .Y(top_core_EC_mc_n622)
         );
  XOR2X1 U9710 ( .A(top_core_EC_mc_n100), .B(top_core_EC_mc_n626), .Y(
        top_core_EC_mc_n625) );
  OAI22X1 U9711 ( .A0(top_core_EC_mc_n609), .A1(n2477), .B0(n2379), .B1(
        top_core_EC_mc_n610), .Y(top_core_EC_mix_out_26_) );
  XOR2X1 U9712 ( .A(top_core_EC_mc_n611), .B(top_core_EC_mc_n612), .Y(
        top_core_EC_mc_n610) );
  XNOR2X1 U9713 ( .A(top_core_EC_mc_mix_in_2_26_), .B(top_core_EC_mc_n613), 
        .Y(top_core_EC_mc_n609) );
  XOR2X1 U9714 ( .A(top_core_EC_mc_n613), .B(top_core_EC_mc_n614), .Y(
        top_core_EC_mc_n612) );
  OAI22X1 U9715 ( .A0(top_core_EC_mc_n588), .A1(n2478), .B0(n2379), .B1(
        top_core_EC_mc_n589), .Y(top_core_EC_mix_out_29_) );
  XOR2X1 U9716 ( .A(top_core_EC_mc_n590), .B(top_core_EC_mc_n591), .Y(
        top_core_EC_mc_n589) );
  XNOR2X1 U9717 ( .A(top_core_EC_mc_mix_in_8[31]), .B(top_core_EC_mc_n592), 
        .Y(top_core_EC_mc_n588) );
  XOR2X1 U9718 ( .A(top_core_EC_mc_n592), .B(top_core_EC_mc_n593), .Y(
        top_core_EC_mc_n591) );
  OAI22X1 U9719 ( .A0(top_core_EC_mc_n572), .A1(n2479), .B0(n2379), .B1(
        top_core_EC_mc_n573), .Y(top_core_EC_mix_out_30_) );
  XOR2X1 U9720 ( .A(top_core_EC_mc_n574), .B(top_core_EC_mc_n575), .Y(
        top_core_EC_mc_n573) );
  XNOR2X1 U9721 ( .A(n1547), .B(top_core_EC_mc_n576), .Y(top_core_EC_mc_n572)
         );
  XOR2X1 U9722 ( .A(top_core_EC_mc_n576), .B(top_core_EC_mc_n577), .Y(
        top_core_EC_mc_n575) );
  OAI22X1 U9723 ( .A0(top_core_EC_mc_n565), .A1(n2479), .B0(n2379), .B1(
        top_core_EC_mc_n566), .Y(top_core_EC_mix_out_31_) );
  XOR2X1 U9724 ( .A(top_core_EC_mc_n567), .B(top_core_EC_mc_n568), .Y(
        top_core_EC_mc_n566) );
  XNOR2X1 U9725 ( .A(n1546), .B(top_core_EC_mc_n569), .Y(top_core_EC_mc_n565)
         );
  XOR2X1 U9726 ( .A(top_core_EC_mc_n569), .B(top_core_EC_mc_n570), .Y(
        top_core_EC_mc_n568) );
  OAI22X1 U9727 ( .A0(top_core_EC_mc_n557), .A1(n2480), .B0(n2379), .B1(
        top_core_EC_mc_n558), .Y(top_core_EC_mix_out_32_) );
  XOR2X1 U9728 ( .A(top_core_EC_mc_n559), .B(top_core_EC_mc_n560), .Y(
        top_core_EC_mc_n558) );
  XNOR2X1 U9729 ( .A(top_core_EC_mix_in[56]), .B(top_core_EC_mc_n561), .Y(
        top_core_EC_mc_n557) );
  XNOR2X1 U9730 ( .A(top_core_EC_mix_in[56]), .B(top_core_EC_mc_n449), .Y(
        top_core_EC_mc_n559) );
  OAI22X1 U9731 ( .A0(top_core_EC_mc_n549), .A1(n2480), .B0(n2379), .B1(
        top_core_EC_mc_n550), .Y(top_core_EC_mix_out_33_) );
  XOR2X1 U9732 ( .A(top_core_EC_mc_n551), .B(top_core_EC_mc_n552), .Y(
        top_core_EC_mc_n550) );
  XNOR2X1 U9733 ( .A(top_core_EC_mc_mix_in_2_58_), .B(top_core_EC_mc_n553), 
        .Y(top_core_EC_mc_n549) );
  XNOR2X1 U9734 ( .A(top_core_EC_mc_mix_in_2_58_), .B(top_core_EC_mc_n441), 
        .Y(top_core_EC_mc_n551) );
  OAI22X1 U9735 ( .A0(top_core_EC_mc_n487), .A1(n2483), .B0(n2375), .B1(
        top_core_EC_mc_n488), .Y(top_core_EC_mix_out_40_) );
  XOR2X1 U9736 ( .A(top_core_EC_mc_n489), .B(top_core_EC_mc_n490), .Y(
        top_core_EC_mc_n488) );
  XNOR2X1 U9737 ( .A(n1542), .B(top_core_EC_mc_n491), .Y(top_core_EC_mc_n487)
         );
  XNOR2X1 U9738 ( .A(n1542), .B(top_core_EC_mc_n449), .Y(top_core_EC_mc_n489)
         );
  OAI22X1 U9739 ( .A0(top_core_EC_mc_n477), .A1(n2483), .B0(n2380), .B1(
        top_core_EC_mc_n478), .Y(top_core_EC_mix_out_42_) );
  XOR2X1 U9740 ( .A(top_core_EC_mc_n479), .B(top_core_EC_mc_n480), .Y(
        top_core_EC_mc_n478) );
  XNOR2X1 U9741 ( .A(top_core_EC_mc_mix_in_2_42_), .B(top_core_EC_mc_n481), 
        .Y(top_core_EC_mc_n477) );
  XNOR2X1 U9742 ( .A(top_core_EC_mc_mix_in_2_42_), .B(top_core_EC_mc_n424), 
        .Y(top_core_EC_mc_n479) );
  OAI22X1 U9743 ( .A0(top_core_EC_mc_n462), .A1(n2484), .B0(n2380), .B1(
        top_core_EC_mc_n463), .Y(top_core_EC_mix_out_45_) );
  XOR2X1 U9744 ( .A(top_core_EC_mc_n464), .B(top_core_EC_mc_n465), .Y(
        top_core_EC_mc_n463) );
  XNOR2X1 U9745 ( .A(top_core_EC_mc_mix_in_8[47]), .B(top_core_EC_mc_n466), 
        .Y(top_core_EC_mc_n462) );
  XNOR2X1 U9746 ( .A(top_core_EC_mc_mix_in_8[47]), .B(top_core_EC_mc_n400), 
        .Y(top_core_EC_mc_n464) );
  OAI22X1 U9747 ( .A0(top_core_EC_mc_n457), .A1(n2472), .B0(n2380), .B1(
        top_core_EC_mc_n458), .Y(top_core_EC_mix_out_46_) );
  XOR2X1 U9748 ( .A(top_core_EC_mc_n459), .B(top_core_EC_mc_n460), .Y(
        top_core_EC_mc_n458) );
  XNOR2X1 U9749 ( .A(n1544), .B(top_core_EC_mc_n461), .Y(top_core_EC_mc_n457)
         );
  XNOR2X1 U9750 ( .A(n1544), .B(top_core_EC_mc_n392), .Y(top_core_EC_mc_n459)
         );
  OAI22X1 U9751 ( .A0(top_core_EC_mc_n452), .A1(n2471), .B0(n2380), .B1(
        top_core_EC_mc_n453), .Y(top_core_EC_mix_out_47_) );
  XOR2X1 U9752 ( .A(top_core_EC_mc_n454), .B(top_core_EC_mc_n455), .Y(
        top_core_EC_mc_n453) );
  XNOR2X1 U9753 ( .A(n1543), .B(top_core_EC_mc_n456), .Y(top_core_EC_mc_n452)
         );
  XNOR2X1 U9754 ( .A(n1543), .B(top_core_EC_mc_n384), .Y(top_core_EC_mc_n454)
         );
  OAI22X1 U9755 ( .A0(top_core_EC_mc_n436), .A1(n2463), .B0(n2380), .B1(
        top_core_EC_mc_n437), .Y(top_core_EC_mix_out_49_) );
  XOR2X1 U9756 ( .A(top_core_EC_mc_n365), .B(top_core_EC_mc_n438), .Y(
        top_core_EC_mc_n437) );
  XNOR2X1 U9757 ( .A(top_core_EC_mc_mix_in_4_58_), .B(top_core_EC_mc_n439), 
        .Y(top_core_EC_mc_n436) );
  XOR2X1 U9758 ( .A(top_core_EC_mc_n439), .B(top_core_EC_mc_n440), .Y(
        top_core_EC_mc_n438) );
  OAI22X1 U9759 ( .A0(top_core_EC_mc_n419), .A1(n2462), .B0(n2381), .B1(
        top_core_EC_mc_n420), .Y(top_core_EC_mix_out_50_) );
  XOR2X1 U9760 ( .A(top_core_EC_mc_n357), .B(top_core_EC_mc_n421), .Y(
        top_core_EC_mc_n420) );
  XNOR2X1 U9761 ( .A(top_core_EC_mc_mix_in_2_58_), .B(top_core_EC_mc_n422), 
        .Y(top_core_EC_mc_n419) );
  XOR2X1 U9762 ( .A(top_core_EC_mc_n422), .B(top_core_EC_mc_n423), .Y(
        top_core_EC_mc_n421) );
  OAI22X1 U9763 ( .A0(top_core_EC_mc_n411), .A1(n2447), .B0(n2381), .B1(
        top_core_EC_mc_n412), .Y(top_core_EC_mix_out_51_) );
  XOR2X1 U9764 ( .A(top_core_EC_mc_n349), .B(top_core_EC_mc_n413), .Y(
        top_core_EC_mc_n412) );
  XNOR2X1 U9765 ( .A(top_core_EC_mc_mix_in_2_59_), .B(top_core_EC_mc_n414), 
        .Y(top_core_EC_mc_n411) );
  XOR2X1 U9766 ( .A(top_core_EC_mc_n414), .B(top_core_EC_mc_n415), .Y(
        top_core_EC_mc_n413) );
  OAI22X1 U9767 ( .A0(top_core_EC_mc_n403), .A1(n2448), .B0(n2381), .B1(
        top_core_EC_mc_n404), .Y(top_core_EC_mix_out_52_) );
  XOR2X1 U9768 ( .A(top_core_EC_mc_n332), .B(top_core_EC_mc_n405), .Y(
        top_core_EC_mc_n404) );
  XNOR2X1 U9769 ( .A(top_core_EC_mc_mix_in_8[62]), .B(top_core_EC_mc_n406), 
        .Y(top_core_EC_mc_n403) );
  XOR2X1 U9770 ( .A(top_core_EC_mc_n406), .B(top_core_EC_mc_n407), .Y(
        top_core_EC_mc_n405) );
  OAI22X1 U9771 ( .A0(top_core_EC_mc_n363), .A1(n2484), .B0(n2381), .B1(
        top_core_EC_mc_n364), .Y(top_core_EC_mix_out_57_) );
  XOR2X1 U9772 ( .A(top_core_EC_mc_n365), .B(top_core_EC_mc_n366), .Y(
        top_core_EC_mc_n364) );
  XNOR2X1 U9773 ( .A(top_core_EC_mc_mix_in_4_58_), .B(top_core_EC_mc_n367), 
        .Y(top_core_EC_mc_n363) );
  XOR2X1 U9774 ( .A(top_core_EC_mc_n367), .B(top_core_EC_mc_n368), .Y(
        top_core_EC_mc_n366) );
  NAND2X1 U9775 ( .A(n338), .B(n1138), .Y(n13879) );
  NAND2X1 U9776 ( .A(n337), .B(n999), .Y(n17029) );
  NAND2X1 U9777 ( .A(n339), .B(n943), .Y(n18289) );
  NAND2X1 U9778 ( .A(n340), .B(n1083), .Y(n15139) );
  NAND2X1 U9779 ( .A(n341), .B(n1069), .Y(n15454) );
  NAND2X1 U9780 ( .A(n342), .B(n1013), .Y(n16714) );
  NAND2X1 U9781 ( .A(n343), .B(n929), .Y(n18604) );
  NAND2X1 U9782 ( .A(n344), .B(n1097), .Y(n14824) );
  NAND2X1 U9783 ( .A(n345), .B(n1027), .Y(n16399) );
  NAND2X1 U9784 ( .A(n346), .B(n957), .Y(n17974) );
  NAND2X1 U9785 ( .A(n347), .B(n1111), .Y(n14509) );
  NAND2X1 U9786 ( .A(n348), .B(n1041), .Y(n16084) );
  NAND2X1 U9787 ( .A(n349), .B(n971), .Y(n17659) );
  NAND2X1 U9788 ( .A(n350), .B(n1125), .Y(n14194) );
  NAND2X1 U9789 ( .A(n351), .B(n1055), .Y(n15769) );
  NAND2X1 U9790 ( .A(n352), .B(n985), .Y(n17344) );
  CLKINVX3 U9791 ( .A(n10068), .Y(n5384) );
  CLKINVX3 U9792 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n254), .Y(n6169) );
  CLKINVX3 U9793 ( .A(n11236), .Y(n5030) );
  CLKINVX3 U9794 ( .A(n8316), .Y(n5856) );
  CLKINVX3 U9795 ( .A(n10944), .Y(n5114) );
  CLKINVX3 U9796 ( .A(n9192), .Y(n5620) );
  CLKINVX3 U9797 ( .A(n7440), .Y(n6084) );
  CLKINVX3 U9798 ( .A(n10360), .Y(n5300) );
  CLKINVX3 U9799 ( .A(n9484), .Y(n5544) );
  CLKINVX3 U9800 ( .A(n8608), .Y(n5772) );
  CLKINVX3 U9801 ( .A(n7732), .Y(n6008) );
  CLKINVX3 U9802 ( .A(n11528), .Y(n4914) );
  CLKINVX3 U9803 ( .A(n10652), .Y(n5222) );
  CLKINVX3 U9804 ( .A(n9776), .Y(n5468) );
  CLKINVX3 U9805 ( .A(n8900), .Y(n5696) );
  CLKINVX3 U9806 ( .A(n8024), .Y(n5932) );
  NAND2X1 U9807 ( .A(n1191), .B(n1738), .Y(n12617) );
  NAND2X1 U9808 ( .A(n1200), .B(n1709), .Y(n12932) );
  NAND2X1 U9809 ( .A(n1151), .B(n1680), .Y(n13247) );
  NAND2X1 U9810 ( .A(n1160), .B(n1652), .Y(n13562) );
  AOI31X1 U9811 ( .A0(n11672), .A1(n11673), .A2(n11650), .B0(n11674), .Y(
        n11667) );
  AOI31X1 U9812 ( .A0(top_core_KE_sb1_n97), .A1(top_core_KE_sb1_n98), .A2(
        top_core_KE_sb1_n75), .B0(top_core_KE_sb1_n99), .Y(top_core_KE_sb1_n92) );
  AOI31X1 U9813 ( .A0(n11988), .A1(n11989), .A2(n11966), .B0(n11990), .Y(
        n11983) );
  AOI31X1 U9814 ( .A0(n12934), .A1(n12935), .A2(n12912), .B0(n12936), .Y(
        n12929) );
  AOI31X1 U9815 ( .A0(n13564), .A1(n13565), .A2(n13542), .B0(n13566), .Y(
        n13559) );
  AOI31X1 U9816 ( .A0(n12619), .A1(n12620), .A2(n12597), .B0(n12621), .Y(
        n12614) );
  CLKINVX2 U9817 ( .A(n106), .Y(n5363) );
  CLKINVX2 U9818 ( .A(n107), .Y(n6131) );
  CLKINVX2 U9819 ( .A(n108), .Y(n5009) );
  CLKINVX2 U9820 ( .A(n109), .Y(n5835) );
  CLKINVX2 U9821 ( .A(n110), .Y(n5751) );
  CLKINVX2 U9822 ( .A(n111), .Y(n4893) );
  CLKINVX2 U9823 ( .A(n112), .Y(n5447) );
  CLKINVX2 U9824 ( .A(n113), .Y(n5911) );
  CLKINVX2 U9825 ( .A(n114), .Y(n5523) );
  CLKINVX2 U9826 ( .A(n115), .Y(n5093) );
  CLKINVX2 U9827 ( .A(n116), .Y(n5987) );
  CLKINVX2 U9828 ( .A(n117), .Y(n5599) );
  CLKINVX2 U9829 ( .A(n118), .Y(n5201) );
  CLKINVX2 U9830 ( .A(n119), .Y(n6063) );
  CLKINVX2 U9831 ( .A(n120), .Y(n5675) );
  CLKINVX2 U9832 ( .A(n121), .Y(n5279) );
  OAI221XL U9833 ( .A0(n14095), .A1(n13847), .B0(n3448), .B1(n14096), .C0(
        n14097), .Y(n14094) );
  AOI211X1 U9834 ( .A0(n6118), .A1(n14100), .B0(n14101), .C0(n14102), .Y(
        n14096) );
  AOI211X1 U9835 ( .A0(n6151), .A1(n449), .B0(n14106), .C0(n14107), .Y(n14095)
         );
  OAI221XL U9836 ( .A0(n17245), .A1(n16997), .B0(n2847), .B1(n17246), .C0(
        n17247), .Y(n17244) );
  AOI211X1 U9837 ( .A0(n5335), .A1(n17250), .B0(n17251), .C0(n17252), .Y(
        n17246) );
  AOI211X1 U9838 ( .A0(n5380), .A1(n450), .B0(n17256), .C0(n17257), .Y(n17245)
         );
  OAI221XL U9839 ( .A0(n18505), .A1(n18257), .B0(n2605), .B1(n18506), .C0(
        n18507), .Y(n18504) );
  AOI211X1 U9840 ( .A0(n4981), .A1(n18510), .B0(n18511), .C0(n18512), .Y(
        n18506) );
  AOI211X1 U9841 ( .A0(n5026), .A1(n451), .B0(n18516), .C0(n18517), .Y(n18505)
         );
  OAI221XL U9842 ( .A0(n15355), .A1(n15107), .B0(n3207), .B1(n15356), .C0(
        n15357), .Y(n15354) );
  AOI211X1 U9843 ( .A0(n5807), .A1(n15360), .B0(n15361), .C0(n15362), .Y(
        n15356) );
  AOI211X1 U9844 ( .A0(n5852), .A1(n452), .B0(n15366), .C0(n15367), .Y(n15355)
         );
  OAI221XL U9845 ( .A0(n15670), .A1(n15422), .B0(n3146), .B1(n15671), .C0(
        n15672), .Y(n15669) );
  AOI211X1 U9846 ( .A0(n5723), .A1(n15675), .B0(n15676), .C0(n15677), .Y(
        n15671) );
  AOI211X1 U9847 ( .A0(n5768), .A1(n453), .B0(n15681), .C0(n15682), .Y(n15670)
         );
  OAI221XL U9848 ( .A0(n18820), .A1(n18572), .B0(n2544), .B1(n18821), .C0(
        n18822), .Y(n18819) );
  AOI211X1 U9849 ( .A0(n4865), .A1(n18825), .B0(n18826), .C0(n18827), .Y(
        n18821) );
  AOI211X1 U9850 ( .A0(n4910), .A1(n454), .B0(n18831), .C0(n18832), .Y(n18820)
         );
  OAI221XL U9851 ( .A0(n16930), .A1(n16682), .B0(n2908), .B1(n16931), .C0(
        n16932), .Y(n16929) );
  AOI211X1 U9852 ( .A0(n5419), .A1(n16935), .B0(n16936), .C0(n16937), .Y(
        n16931) );
  AOI211X1 U9853 ( .A0(n5464), .A1(n455), .B0(n16941), .C0(n16942), .Y(n16930)
         );
  OAI221XL U9854 ( .A0(n15040), .A1(n14792), .B0(n3268), .B1(n15041), .C0(
        n15042), .Y(n15039) );
  AOI211X1 U9855 ( .A0(n5883), .A1(n15045), .B0(n15046), .C0(n15047), .Y(
        n15041) );
  AOI211X1 U9856 ( .A0(n5928), .A1(n456), .B0(n15051), .C0(n15052), .Y(n15040)
         );
  OAI221XL U9857 ( .A0(n16615), .A1(n16367), .B0(n2969), .B1(n16616), .C0(
        n16617), .Y(n16614) );
  AOI211X1 U9858 ( .A0(n5495), .A1(n16620), .B0(n16621), .C0(n16622), .Y(
        n16616) );
  AOI211X1 U9859 ( .A0(n5540), .A1(n457), .B0(n16626), .C0(n16627), .Y(n16615)
         );
  OAI221XL U9860 ( .A0(n18190), .A1(n17942), .B0(n2666), .B1(n18191), .C0(
        n18192), .Y(n18189) );
  AOI211X1 U9861 ( .A0(n5065), .A1(n18195), .B0(n18196), .C0(n18197), .Y(
        n18191) );
  AOI211X1 U9862 ( .A0(n5110), .A1(n458), .B0(n18201), .C0(n18202), .Y(n18190)
         );
  OAI221XL U9863 ( .A0(n14725), .A1(n14477), .B0(n3329), .B1(n14726), .C0(
        n14727), .Y(n14724) );
  AOI211X1 U9864 ( .A0(n5959), .A1(n14730), .B0(n14731), .C0(n14732), .Y(
        n14726) );
  AOI211X1 U9865 ( .A0(n6004), .A1(n459), .B0(n14736), .C0(n14737), .Y(n14725)
         );
  OAI221XL U9866 ( .A0(n16300), .A1(n16052), .B0(n3027), .B1(n16301), .C0(
        n16302), .Y(n16299) );
  AOI211X1 U9867 ( .A0(n5571), .A1(n16305), .B0(n16306), .C0(n16307), .Y(
        n16301) );
  AOI211X1 U9868 ( .A0(n5616), .A1(n460), .B0(n16311), .C0(n16312), .Y(n16300)
         );
  OAI221XL U9869 ( .A0(n17875), .A1(n17627), .B0(n2726), .B1(n17876), .C0(
        n17877), .Y(n17874) );
  AOI211X1 U9870 ( .A0(n5173), .A1(n17880), .B0(n17881), .C0(n17882), .Y(
        n17876) );
  AOI211X1 U9871 ( .A0(n5218), .A1(n461), .B0(n17886), .C0(n17887), .Y(n17875)
         );
  OAI221XL U9872 ( .A0(n14410), .A1(n14162), .B0(n3387), .B1(n14411), .C0(
        n14412), .Y(n14409) );
  AOI211X1 U9873 ( .A0(n6035), .A1(n14415), .B0(n14416), .C0(n14417), .Y(
        n14411) );
  AOI211X1 U9874 ( .A0(n6080), .A1(n462), .B0(n14421), .C0(n14422), .Y(n14410)
         );
  OAI221XL U9875 ( .A0(n15985), .A1(n15737), .B0(n3088), .B1(n15986), .C0(
        n15987), .Y(n15984) );
  AOI211X1 U9876 ( .A0(n5647), .A1(n15990), .B0(n15991), .C0(n15992), .Y(
        n15986) );
  AOI211X1 U9877 ( .A0(n5692), .A1(n463), .B0(n15996), .C0(n15997), .Y(n15985)
         );
  OAI221XL U9878 ( .A0(n17560), .A1(n17312), .B0(n2787), .B1(n17561), .C0(
        n17562), .Y(n17559) );
  AOI211X1 U9879 ( .A0(n5251), .A1(n17565), .B0(n17566), .C0(n17567), .Y(
        n17561) );
  AOI211X1 U9880 ( .A0(n5296), .A1(n464), .B0(n17571), .C0(n17572), .Y(n17560)
         );
  XOR2X1 U9881 ( .A(top_core_EC_mc_mix_in_2_16_), .B(top_core_EC_mix_in[16]), 
        .Y(top_core_EC_mc_mix_in_4_18_) );
  XOR2X1 U9882 ( .A(top_core_EC_mc_mix_in_2_32_), .B(top_core_EC_mix_in[32]), 
        .Y(top_core_EC_mc_mix_in_4_34_) );
  XOR2X1 U9883 ( .A(top_core_EC_mc_mix_in_2_32_), .B(top_core_EC_mix_in[35]), 
        .Y(top_core_EC_mc_mix_in_8[38]) );
  AOI31X1 U9884 ( .A0(n12931), .A1(n12932), .A2(n12933), .B0(n1696), .Y(n12930) );
  AOI31X1 U9885 ( .A0(n12616), .A1(n12617), .A2(n12618), .B0(n1725), .Y(n12615) );
  XNOR2X1 U9886 ( .A(top_core_EC_mc_n927), .B(top_core_EC_mc_n928), .Y(
        top_core_EC_mc_n101) );
  XNOR2X1 U9887 ( .A(top_core_EC_mc_mix_in_8[16]), .B(
        top_core_EC_mc_mix_in_8[0]), .Y(top_core_EC_mc_n927) );
  XOR2X1 U9888 ( .A(n1550), .B(n1547), .Y(top_core_EC_mc_n928) );
  XNOR2X1 U9889 ( .A(top_core_EC_mc_n675), .B(top_core_EC_mc_n676), .Y(
        top_core_EC_mc_n8) );
  XNOR2X1 U9890 ( .A(top_core_EC_mc_mix_in_8[1]), .B(
        top_core_EC_mc_mix_in_8[17]), .Y(top_core_EC_mc_n675) );
  XOR2X1 U9891 ( .A(top_core_EC_mc_mix_in_8[9]), .B(
        top_core_EC_mc_mix_in_8[25]), .Y(top_core_EC_mc_n676) );
  XOR2X1 U9892 ( .A(top_core_EC_mc_mix_in_8[0]), .B(top_core_EC_mc_mix_in_4_0_), .Y(top_core_EC_mc_mix_in_8[1]) );
  XNOR2X1 U9893 ( .A(top_core_EC_mc_n777), .B(top_core_EC_mc_n778), .Y(
        top_core_EC_mc_n498) );
  XNOR2X1 U9894 ( .A(top_core_EC_mc_mix_in_8[19]), .B(
        top_core_EC_mc_mix_in_8[11]), .Y(top_core_EC_mc_n777) );
  XOR2X1 U9895 ( .A(top_core_EC_mc_mix_in_8[3]), .B(
        top_core_EC_mc_mix_in_8[27]), .Y(top_core_EC_mc_n778) );
  XOR2X1 U9896 ( .A(top_core_EC_mc_mix_in_8[16]), .B(
        top_core_EC_mc_mix_in_4_18_), .Y(top_core_EC_mc_mix_in_8[19]) );
  XNOR2X1 U9897 ( .A(top_core_EC_mc_n710), .B(top_core_EC_mc_n711), .Y(
        top_core_EC_mc_n433) );
  XNOR2X1 U9898 ( .A(top_core_EC_mc_mix_in_8[20]), .B(
        top_core_EC_mc_mix_in_8[12]), .Y(top_core_EC_mc_n710) );
  XOR2X1 U9899 ( .A(top_core_EC_mc_mix_in_8[4]), .B(
        top_core_EC_mc_mix_in_8[28]), .Y(top_core_EC_mc_n711) );
  XOR2X1 U9900 ( .A(top_core_EC_mc_mix_in_8[16]), .B(
        top_core_EC_mc_mix_in_4_19_), .Y(top_core_EC_mc_mix_in_8[20]) );
  XNOR2X1 U9901 ( .A(top_core_EC_mc_n689), .B(top_core_EC_mc_n690), .Y(
        top_core_EC_mc_n190) );
  XNOR2X1 U9902 ( .A(top_core_EC_mc_mix_in_8[23]), .B(
        top_core_EC_mc_mix_in_8[15]), .Y(top_core_EC_mc_n689) );
  XOR2X1 U9903 ( .A(top_core_EC_mc_mix_in_8[7]), .B(
        top_core_EC_mc_mix_in_8[31]), .Y(top_core_EC_mc_n690) );
  XNOR2X1 U9904 ( .A(top_core_EC_mc_n554), .B(top_core_EC_mc_n555), .Y(
        top_core_EC_mc_n441) );
  XNOR2X1 U9905 ( .A(top_core_EC_mc_mix_in_8[41]), .B(
        top_core_EC_mc_mix_in_8[33]), .Y(top_core_EC_mc_n554) );
  XOR2X1 U9906 ( .A(top_core_EC_mc_mix_in_8[57]), .B(
        top_core_EC_mc_mix_in_8[49]), .Y(top_core_EC_mc_n555) );
  XOR2X1 U9907 ( .A(n1544), .B(n1543), .Y(top_core_EC_mc_mix_in_8[41]) );
  XNOR2X1 U9908 ( .A(top_core_EC_mc_n546), .B(top_core_EC_mc_n547), .Y(
        top_core_EC_mc_n424) );
  XNOR2X1 U9909 ( .A(top_core_EC_mc_mix_in_8[42]), .B(
        top_core_EC_mc_mix_in_8[34]), .Y(top_core_EC_mc_n546) );
  XOR2X1 U9910 ( .A(top_core_EC_mc_mix_in_8[58]), .B(
        top_core_EC_mc_mix_in_8[50]), .Y(top_core_EC_mc_n547) );
  XNOR2X1 U9911 ( .A(top_core_EC_mc_n538), .B(top_core_EC_mc_n539), .Y(
        top_core_EC_mc_n416) );
  XNOR2X1 U9912 ( .A(top_core_EC_mc_mix_in_8[43]), .B(
        top_core_EC_mc_mix_in_8[35]), .Y(top_core_EC_mc_n538) );
  XOR2X1 U9913 ( .A(top_core_EC_mc_mix_in_8[59]), .B(
        top_core_EC_mc_mix_in_8[51]), .Y(top_core_EC_mc_n539) );
  XOR2X1 U9914 ( .A(n1544), .B(top_core_EC_mc_mix_in_4_42_), .Y(
        top_core_EC_mc_mix_in_8[43]) );
  XNOR2X1 U9915 ( .A(top_core_EC_mc_n530), .B(top_core_EC_mc_n531), .Y(
        top_core_EC_mc_n408) );
  XNOR2X1 U9916 ( .A(top_core_EC_mc_mix_in_8[44]), .B(
        top_core_EC_mc_mix_in_8[36]), .Y(top_core_EC_mc_n530) );
  XOR2X1 U9917 ( .A(top_core_EC_mc_mix_in_8[60]), .B(
        top_core_EC_mc_mix_in_8[52]), .Y(top_core_EC_mc_n531) );
  XOR2X1 U9918 ( .A(n1544), .B(top_core_EC_mc_mix_in_4_43_), .Y(
        top_core_EC_mc_mix_in_8[44]) );
  XNOR2X1 U9919 ( .A(top_core_EC_mc_n522), .B(top_core_EC_mc_n523), .Y(
        top_core_EC_mc_n400) );
  XNOR2X1 U9920 ( .A(top_core_EC_mc_mix_in_8[45]), .B(
        top_core_EC_mc_mix_in_8[37]), .Y(top_core_EC_mc_n522) );
  XOR2X1 U9921 ( .A(top_core_EC_mc_mix_in_8[61]), .B(
        top_core_EC_mc_mix_in_8[53]), .Y(top_core_EC_mc_n523) );
  XNOR2X1 U9922 ( .A(top_core_EC_mc_n514), .B(top_core_EC_mc_n515), .Y(
        top_core_EC_mc_n392) );
  XNOR2X1 U9923 ( .A(top_core_EC_mc_mix_in_8[46]), .B(
        top_core_EC_mc_mix_in_8[38]), .Y(top_core_EC_mc_n514) );
  XOR2X1 U9924 ( .A(top_core_EC_mc_mix_in_8[62]), .B(
        top_core_EC_mc_mix_in_8[54]), .Y(top_core_EC_mc_n515) );
  XNOR2X1 U9925 ( .A(top_core_EC_mc_n287), .B(top_core_EC_mc_n288), .Y(
        top_core_EC_mc_n165) );
  XNOR2X1 U9926 ( .A(top_core_EC_mc_mix_in_8[74]), .B(
        top_core_EC_mc_mix_in_8[66]), .Y(top_core_EC_mc_n287) );
  XOR2X1 U9927 ( .A(top_core_EC_mc_mix_in_8[90]), .B(
        top_core_EC_mc_mix_in_8[82]), .Y(top_core_EC_mc_n288) );
  XNOR2X1 U9928 ( .A(top_core_EC_mc_n263), .B(top_core_EC_mc_n264), .Y(
        top_core_EC_mc_n141) );
  XNOR2X1 U9929 ( .A(top_core_EC_mc_mix_in_8[77]), .B(
        top_core_EC_mc_mix_in_8[69]), .Y(top_core_EC_mc_n263) );
  XOR2X1 U9930 ( .A(top_core_EC_mc_mix_in_8[93]), .B(
        top_core_EC_mc_mix_in_8[85]), .Y(top_core_EC_mc_n264) );
  XNOR2X1 U9931 ( .A(top_core_EC_mc_n246), .B(top_core_EC_mc_n247), .Y(
        top_core_EC_mc_n133) );
  XNOR2X1 U9932 ( .A(top_core_EC_mc_mix_in_8[78]), .B(
        top_core_EC_mc_mix_in_8[70]), .Y(top_core_EC_mc_n246) );
  XOR2X1 U9933 ( .A(top_core_EC_mc_mix_in_8[94]), .B(
        top_core_EC_mc_mix_in_8[86]), .Y(top_core_EC_mc_n247) );
  XNOR2X1 U9934 ( .A(top_core_EC_mc_n874), .B(top_core_EC_mc_n875), .Y(
        top_core_EC_mc_n26) );
  XNOR2X1 U9935 ( .A(top_core_EC_mc_mix_in_8[114]), .B(
        top_core_EC_mc_mix_in_8[106]), .Y(top_core_EC_mc_n874) );
  XOR2X1 U9936 ( .A(top_core_EC_mc_mix_in_8[98]), .B(
        top_core_EC_mc_mix_in_8[122]), .Y(top_core_EC_mc_n875) );
  XNOR2X1 U9937 ( .A(top_core_EC_mc_n911), .B(top_core_EC_mc_n912), .Y(
        top_core_EC_mc_n800) );
  XNOR2X1 U9938 ( .A(top_core_EC_mc_mix_in_8[109]), .B(
        top_core_EC_mc_mix_in_8[101]), .Y(top_core_EC_mc_n911) );
  XOR2X1 U9939 ( .A(top_core_EC_mc_mix_in_8[125]), .B(
        top_core_EC_mc_mix_in_8[117]), .Y(top_core_EC_mc_n912) );
  XNOR2X1 U9940 ( .A(top_core_EC_mc_n903), .B(top_core_EC_mc_n904), .Y(
        top_core_EC_mc_n792) );
  XNOR2X1 U9941 ( .A(top_core_EC_mc_mix_in_8[110]), .B(
        top_core_EC_mc_mix_in_8[102]), .Y(top_core_EC_mc_n903) );
  XOR2X1 U9942 ( .A(top_core_EC_mc_mix_in_8[126]), .B(
        top_core_EC_mc_mix_in_8[118]), .Y(top_core_EC_mc_n904) );
  OAI221XL U9943 ( .A0(n2861), .A1(n10165), .B0(n10166), .B1(n2853), .C0(
        n10074), .Y(n10159) );
  NAND2XL U9944 ( .A(n9905), .B(n9888), .Y(n10168) );
  OAI221XL U9945 ( .A0(n3461), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n351), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n352), .B1(n3454), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n260), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n345) );
  NAND2XL U9946 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n88), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n70), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n354) );
  OAI221XL U9947 ( .A0(n3221), .A1(n8413), .B0(n8414), .B1(n3213), .C0(n8322), 
        .Y(n8407) );
  NAND2XL U9948 ( .A(n8153), .B(n8136), .Y(n8416) );
  OAI221XL U9949 ( .A0(n2621), .A1(n11333), .B0(n11334), .B1(n2611), .C0(
        n11242), .Y(n11327) );
  NAND2XL U9950 ( .A(n11073), .B(n11056), .Y(n11336) );
  OAI221XL U9951 ( .A0(n2680), .A1(n11041), .B0(n11042), .B1(n2672), .C0(
        n10950), .Y(n11035) );
  NAND2XL U9952 ( .A(n10781), .B(n10764), .Y(n11044) );
  OAI221XL U9953 ( .A0(n3403), .A1(n7537), .B0(n7538), .B1(n3393), .C0(n7446), 
        .Y(n7531) );
  NAND2XL U9954 ( .A(n7277), .B(n7260), .Y(n7540) );
  OAI221XL U9955 ( .A0(n3043), .A1(n9289), .B0(n9290), .B1(n3033), .C0(n9198), 
        .Y(n9283) );
  NAND2XL U9956 ( .A(n9029), .B(n9012), .Y(n9292) );
  OAI221XL U9957 ( .A0(n2803), .A1(n10457), .B0(n10458), .B1(n2793), .C0(
        n10366), .Y(n10451) );
  NAND2XL U9958 ( .A(n10197), .B(n10180), .Y(n10460) );
  OAI221XL U9959 ( .A0(n2985), .A1(n9581), .B0(n9582), .B1(n2975), .C0(n9490), 
        .Y(n9575) );
  NAND2XL U9960 ( .A(n9321), .B(n9304), .Y(n9584) );
  OAI221XL U9961 ( .A0(n3162), .A1(n8705), .B0(n8706), .B1(n3152), .C0(n8614), 
        .Y(n8699) );
  NAND2XL U9962 ( .A(n8445), .B(n8428), .Y(n8708) );
  OAI221XL U9963 ( .A0(n3345), .A1(n7829), .B0(n7830), .B1(n3335), .C0(n7738), 
        .Y(n7823) );
  NAND2XL U9964 ( .A(n7569), .B(n7552), .Y(n7832) );
  OAI221XL U9965 ( .A0(n2554), .A1(n11625), .B0(n11626), .B1(n2550), .C0(
        n11534), .Y(n11619) );
  NAND2XL U9966 ( .A(n11365), .B(n11348), .Y(n11628) );
  OAI221XL U9967 ( .A0(n2740), .A1(n10749), .B0(n10750), .B1(n2732), .C0(
        n10658), .Y(n10743) );
  NAND2XL U9968 ( .A(n10489), .B(n10472), .Y(n10752) );
  OAI221XL U9969 ( .A0(n2924), .A1(n9873), .B0(n9874), .B1(n2914), .C0(n9782), 
        .Y(n9867) );
  NAND2XL U9970 ( .A(n9613), .B(n9596), .Y(n9876) );
  OAI221XL U9971 ( .A0(n3102), .A1(n8997), .B0(n8998), .B1(n3094), .C0(n8906), 
        .Y(n8991) );
  NAND2XL U9972 ( .A(n8737), .B(n8720), .Y(n9000) );
  OAI221XL U9973 ( .A0(n3284), .A1(n8121), .B0(n8122), .B1(n3274), .C0(n8030), 
        .Y(n8115) );
  NAND2XL U9974 ( .A(n7861), .B(n7844), .Y(n8124) );
  OAI221XL U9975 ( .A0(n1222), .A1(n11675), .B0(n11651), .B1(n11883), .C0(
        n11676), .Y(n11882) );
  OAI221XL U9976 ( .A0(n1216), .A1(top_core_KE_sb1_n100), .B0(
        top_core_KE_sb1_n76), .B1(top_core_KE_sb1_n312), .C0(
        top_core_KE_sb1_n101), .Y(top_core_KE_sb1_n311) );
  OAI221XL U9977 ( .A0(n1181), .A1(n12306), .B0(n12283), .B1(n12514), .C0(
        n12307), .Y(n12513) );
  OAI221XL U9978 ( .A0(n1173), .A1(n13252), .B0(n13228), .B1(n13459), .C0(
        n13253), .Y(n13458) );
  OAI221XL U9979 ( .A0(n1176), .A1(n11991), .B0(n11967), .B1(n12199), .C0(
        n11992), .Y(n12198) );
  OAI221XL U9980 ( .A0(n1213), .A1(n12622), .B0(n12598), .B1(n12829), .C0(
        n12623), .Y(n12828) );
  OAI221XL U9981 ( .A0(n1178), .A1(n13567), .B0(n13543), .B1(n13774), .C0(
        n13568), .Y(n13773) );
  OAI221XL U9982 ( .A0(n1219), .A1(n12937), .B0(n12913), .B1(n13144), .C0(
        n12938), .Y(n13143) );
  XOR2X1 U9983 ( .A(top_core_EC_mc_mix_in_2_0_), .B(top_core_EC_mix_in[0]), 
        .Y(top_core_EC_mc_mix_in_4_2_) );
  XOR2X1 U9984 ( .A(top_core_EC_mc_mix_in_2_48_), .B(top_core_EC_mix_in[48]), 
        .Y(top_core_EC_mc_mix_in_4_50_) );
  XOR2X1 U9985 ( .A(top_core_EC_mc_mix_in_2_48_), .B(top_core_EC_mix_in[51]), 
        .Y(top_core_EC_mc_mix_in_8[54]) );
  AOI21X1 U9986 ( .A0(n5353), .A1(n529), .B0(n17161), .Y(n17160) );
  AOI21X1 U9987 ( .A0(n6121), .A1(n530), .B0(n14011), .Y(n14010) );
  AOI21X1 U9988 ( .A0(n4999), .A1(n531), .B0(n18421), .Y(n18420) );
  AOI21X1 U9989 ( .A0(n5825), .A1(n532), .B0(n15271), .Y(n15270) );
  AOI21X1 U9990 ( .A0(n5741), .A1(n538), .B0(n15586), .Y(n15585) );
  AOI21X1 U9991 ( .A0(n4883), .A1(n540), .B0(n18736), .Y(n18735) );
  AOI21X1 U9992 ( .A0(n5437), .A1(n542), .B0(n16846), .Y(n16845) );
  AOI21X1 U9993 ( .A0(n5901), .A1(n544), .B0(n14956), .Y(n14955) );
  AOI21X1 U9994 ( .A0(n5513), .A1(n537), .B0(n16531), .Y(n16530) );
  AOI21X1 U9995 ( .A0(n5083), .A1(n533), .B0(n18106), .Y(n18105) );
  AOI21X1 U9996 ( .A0(n5977), .A1(n539), .B0(n14641), .Y(n14640) );
  AOI21X1 U9997 ( .A0(n5589), .A1(n534), .B0(n16216), .Y(n16215) );
  AOI21X1 U9998 ( .A0(n5191), .A1(n541), .B0(n17791), .Y(n17790) );
  AOI21X1 U9999 ( .A0(n6053), .A1(n535), .B0(n14326), .Y(n14325) );
  AOI21X1 U10000 ( .A0(n5665), .A1(n543), .B0(n15901), .Y(n15900) );
  AOI21X1 U10001 ( .A0(n5269), .A1(n536), .B0(n17476), .Y(n17475) );
  XOR2X1 U10002 ( .A(top_core_EC_mc_mix_in_2_16_), .B(top_core_EC_mix_in[19]), 
        .Y(top_core_EC_mc_mix_in_8[22]) );
  OAI211X1 U10003 ( .A0(n9894), .A1(n9893), .B0(n5367), .C0(n10164), .Y(n10160) );
  INVX1 U10004 ( .A(n9902), .Y(n5367) );
  AOI21X1 U10005 ( .A0(n417), .A1(n9954), .B0(n5340), .Y(n10164) );
  OAI211X1 U10006 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n77), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n76), .B0(n6157), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n350), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n346) );
  INVX1 U10007 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n85), .Y(n6157) );
  AOI21X1 U10008 ( .A0(n418), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n139), 
        .B0(n6136), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n350) );
  OAI211X1 U10009 ( .A0(n8142), .A1(n8141), .B0(n5839), .C0(n8412), .Y(n8408)
         );
  INVX1 U10010 ( .A(n8150), .Y(n5839) );
  AOI21X1 U10011 ( .A0(n420), .A1(n8202), .B0(n5812), .Y(n8412) );
  OAI211X1 U10012 ( .A0(n11062), .A1(n11061), .B0(n5013), .C0(n11332), .Y(
        n11328) );
  INVX1 U10013 ( .A(n11070), .Y(n5013) );
  AOI21X1 U10014 ( .A0(n419), .A1(n11122), .B0(n4986), .Y(n11332) );
  OAI211X1 U10015 ( .A0(n10770), .A1(n10769), .B0(n5097), .C0(n11040), .Y(
        n11036) );
  INVX1 U10016 ( .A(n10778), .Y(n5097) );
  AOI21X1 U10017 ( .A0(n421), .A1(n10830), .B0(n5070), .Y(n11040) );
  OAI211X1 U10018 ( .A0(n7266), .A1(n7265), .B0(n6067), .C0(n7536), .Y(n7532)
         );
  INVX1 U10019 ( .A(n7274), .Y(n6067) );
  AOI21X1 U10020 ( .A0(n423), .A1(n7326), .B0(n6040), .Y(n7536) );
  OAI211X1 U10021 ( .A0(n9018), .A1(n9017), .B0(n5603), .C0(n9288), .Y(n9284)
         );
  INVX1 U10022 ( .A(n9026), .Y(n5603) );
  AOI21X1 U10023 ( .A0(n422), .A1(n9078), .B0(n5576), .Y(n9288) );
  OAI211X1 U10024 ( .A0(n10186), .A1(n10185), .B0(n5283), .C0(n10456), .Y(
        n10452) );
  INVX1 U10025 ( .A(n10194), .Y(n5283) );
  AOI21X1 U10026 ( .A0(n424), .A1(n10246), .B0(n5256), .Y(n10456) );
  OAI211X1 U10027 ( .A0(n9310), .A1(n9309), .B0(n5527), .C0(n9580), .Y(n9576)
         );
  INVX1 U10028 ( .A(n9318), .Y(n5527) );
  AOI21X1 U10029 ( .A0(n425), .A1(n9370), .B0(n5500), .Y(n9580) );
  OAI211X1 U10030 ( .A0(n8434), .A1(n8433), .B0(n5755), .C0(n8704), .Y(n8700)
         );
  INVX1 U10031 ( .A(n8442), .Y(n5755) );
  AOI21X1 U10032 ( .A0(n426), .A1(n8494), .B0(n5728), .Y(n8704) );
  OAI211X1 U10033 ( .A0(n7558), .A1(n7557), .B0(n5991), .C0(n7828), .Y(n7824)
         );
  INVX1 U10034 ( .A(n7566), .Y(n5991) );
  AOI21X1 U10035 ( .A0(n427), .A1(n7618), .B0(n5964), .Y(n7828) );
  OAI211X1 U10036 ( .A0(n11354), .A1(n11353), .B0(n4897), .C0(n11624), .Y(
        n11620) );
  INVX1 U10037 ( .A(n11362), .Y(n4897) );
  AOI21X1 U10038 ( .A0(n428), .A1(n11414), .B0(n4870), .Y(n11624) );
  OAI211X1 U10039 ( .A0(n10478), .A1(n10477), .B0(n5205), .C0(n10748), .Y(
        n10744) );
  INVX1 U10040 ( .A(n10486), .Y(n5205) );
  AOI21X1 U10041 ( .A0(n429), .A1(n10538), .B0(n5178), .Y(n10748) );
  OAI211X1 U10042 ( .A0(n9602), .A1(n9601), .B0(n5451), .C0(n9872), .Y(n9868)
         );
  INVX1 U10043 ( .A(n9610), .Y(n5451) );
  AOI21X1 U10044 ( .A0(n430), .A1(n9662), .B0(n5424), .Y(n9872) );
  OAI211X1 U10045 ( .A0(n8726), .A1(n8725), .B0(n5679), .C0(n8996), .Y(n8992)
         );
  INVX1 U10046 ( .A(n8734), .Y(n5679) );
  AOI21X1 U10047 ( .A0(n431), .A1(n8786), .B0(n5652), .Y(n8996) );
  OAI211X1 U10048 ( .A0(n7850), .A1(n7849), .B0(n5915), .C0(n8120), .Y(n8116)
         );
  INVX1 U10049 ( .A(n7858), .Y(n5915) );
  AOI21X1 U10050 ( .A0(n432), .A1(n7910), .B0(n5888), .Y(n8120) );
  XOR2X1 U10051 ( .A(top_core_EC_mc_mix_in_2_0_), .B(top_core_EC_mix_in[3]), 
        .Y(top_core_EC_mc_mix_in_8[6]) );
  NAND2X1 U10052 ( .A(n6597), .B(n13553), .Y(n13648) );
  AOI31XL U10053 ( .A0(n1003), .A1(n17126), .A2(n17008), .B0(n5332), .Y(n17276) );
  INVX1 U10054 ( .A(n17231), .Y(n5332) );
  AOI31XL U10055 ( .A0(n1142), .A1(n13976), .A2(n13858), .B0(n6116), .Y(n14126) );
  INVX1 U10056 ( .A(n14081), .Y(n6116) );
  AOI31XL U10057 ( .A0(n1087), .A1(n15236), .A2(n15118), .B0(n5804), .Y(n15386) );
  INVX1 U10058 ( .A(n15341), .Y(n5804) );
  AOI31XL U10059 ( .A0(n947), .A1(n18386), .A2(n18268), .B0(n4978), .Y(n18536)
         );
  INVX1 U10060 ( .A(n18491), .Y(n4978) );
  AOI31XL U10061 ( .A0(n1073), .A1(n15551), .A2(n15433), .B0(n5720), .Y(n15701) );
  INVX1 U10062 ( .A(n15656), .Y(n5720) );
  AOI31XL U10063 ( .A0(n1017), .A1(n16811), .A2(n16693), .B0(n5416), .Y(n16961) );
  INVX1 U10064 ( .A(n16916), .Y(n5416) );
  AOI31XL U10065 ( .A0(n933), .A1(n18701), .A2(n18583), .B0(n4862), .Y(n18851)
         );
  INVX1 U10066 ( .A(n18806), .Y(n4862) );
  AOI31XL U10067 ( .A0(n1101), .A1(n14921), .A2(n14803), .B0(n5880), .Y(n15071) );
  INVX1 U10068 ( .A(n15026), .Y(n5880) );
  AOI31XL U10069 ( .A0(n1031), .A1(n16496), .A2(n16378), .B0(n5492), .Y(n16646) );
  INVX1 U10070 ( .A(n16601), .Y(n5492) );
  AOI31XL U10071 ( .A0(n961), .A1(n18071), .A2(n17953), .B0(n5062), .Y(n18221)
         );
  INVX1 U10072 ( .A(n18176), .Y(n5062) );
  AOI31XL U10073 ( .A0(n1115), .A1(n14606), .A2(n14488), .B0(n5956), .Y(n14756) );
  INVX1 U10074 ( .A(n14711), .Y(n5956) );
  AOI31XL U10075 ( .A0(n1045), .A1(n16181), .A2(n16063), .B0(n5568), .Y(n16331) );
  INVX1 U10076 ( .A(n16286), .Y(n5568) );
  AOI31XL U10077 ( .A0(n975), .A1(n17756), .A2(n17638), .B0(n5170), .Y(n17906)
         );
  INVX1 U10078 ( .A(n17861), .Y(n5170) );
  AOI31XL U10079 ( .A0(n1129), .A1(n14291), .A2(n14173), .B0(n6032), .Y(n14441) );
  INVX1 U10080 ( .A(n14396), .Y(n6032) );
  AOI31XL U10081 ( .A0(n1059), .A1(n15866), .A2(n15748), .B0(n5644), .Y(n16016) );
  INVX1 U10082 ( .A(n15971), .Y(n5644) );
  AOI31XL U10083 ( .A0(n989), .A1(n17441), .A2(n17323), .B0(n5248), .Y(n17591)
         );
  INVX1 U10084 ( .A(n17546), .Y(n5248) );
  NAND2X1 U10085 ( .A(n1157), .B(n1651), .Y(n13549) );
  NAND2X1 U10086 ( .A(n1148), .B(n1680), .Y(n13234) );
  NAND2X1 U10087 ( .A(n1197), .B(n1709), .Y(n12919) );
  NAND2X1 U10088 ( .A(n1188), .B(n1738), .Y(n12604) );
  NOR2XL U10089 ( .A(n180), .B(n1687), .Y(n13455) );
  NOR2XL U10090 ( .A(n181), .B(n1745), .Y(n12825) );
  NOR2XL U10091 ( .A(n182), .B(n1716), .Y(n13140) );
  AOI22X1 U10092 ( .A0(n3481), .A1(n3479), .B0(n3472), .B1(n530), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n77) );
  AOI22X1 U10093 ( .A0(n2880), .A1(n2875), .B0(n2871), .B1(n529), .Y(n9894) );
  AOI22X1 U10094 ( .A0(n2638), .A1(n2633), .B0(n2629), .B1(n531), .Y(n11062)
         );
  AOI22X1 U10095 ( .A0(n3240), .A1(n3233), .B0(n3231), .B1(n532), .Y(n8142) );
  AOI22X1 U10096 ( .A0(n2699), .A1(n2696), .B0(n2690), .B1(n533), .Y(n10770)
         );
  AOI22X1 U10097 ( .A0(n3060), .A1(n3055), .B0(n3051), .B1(n534), .Y(n9018) );
  AOI22X1 U10098 ( .A0(n3420), .A1(n3417), .B0(n3411), .B1(n535), .Y(n7266) );
  AOI22X1 U10099 ( .A0(n3002), .A1(n2999), .B0(n2993), .B1(n537), .Y(n9310) );
  AOI22X1 U10100 ( .A0(n3179), .A1(n3172), .B0(n3170), .B1(n538), .Y(n8434) );
  AOI22X1 U10101 ( .A0(n3362), .A1(n3355), .B0(n3353), .B1(n539), .Y(n7558) );
  AOI22X1 U10102 ( .A0(n2577), .A1(n2572), .B0(n2568), .B1(n540), .Y(n11354)
         );
  AOI22X1 U10103 ( .A0(n2759), .A1(n2752), .B0(n2750), .B1(n541), .Y(n10478)
         );
  AOI22X1 U10104 ( .A0(n2941), .A1(n2938), .B0(n2932), .B1(n542), .Y(n9602) );
  AOI22X1 U10105 ( .A0(n3121), .A1(n3116), .B0(n3112), .B1(n543), .Y(n8726) );
  AOI22X1 U10106 ( .A0(n3301), .A1(top_core_EC_ss_in[26]), .B0(n3292), .B1(
        n544), .Y(n7850) );
  AOI22X1 U10107 ( .A0(n2820), .A1(top_core_EC_ss_in[90]), .B0(n2811), .B1(
        n536), .Y(n10186) );
  AOI22XL U10108 ( .A0(n1680), .A1(n6549), .B0(n1275), .B1(n1148), .Y(n13440)
         );
  AOI22XL U10109 ( .A0(n1738), .A1(n6844), .B0(n1269), .B1(n1188), .Y(n12810)
         );
  AOI22XL U10110 ( .A0(n1651), .A1(n6597), .B0(n1278), .B1(n1157), .Y(n13755)
         );
  AOI22XL U10111 ( .A0(n1709), .A1(n6890), .B0(n1272), .B1(n1197), .Y(n13125)
         );
  AOI21X1 U10112 ( .A0(n3484), .A1(n1138), .B0(n1137), .Y(n13934) );
  AOI21X1 U10113 ( .A0(n3182), .A1(n1069), .B0(n1068), .Y(n15509) );
  AOI21X1 U10114 ( .A0(n2884), .A1(n999), .B0(n998), .Y(n17084) );
  AOI21X1 U10115 ( .A0(n2580), .A1(n929), .B0(n928), .Y(n18659) );
  AOI21X1 U10116 ( .A0(n2951), .A1(n1013), .B0(n1012), .Y(n16769) );
  AOI21X1 U10117 ( .A0(n2643), .A1(n943), .B0(n942), .Y(n18344) );
  AOI21X1 U10118 ( .A0(n3243), .A1(n1083), .B0(n1082), .Y(n15194) );
  AOI21X1 U10119 ( .A0(n3304), .A1(n1097), .B0(n1096), .Y(n14879) );
  AOI21X1 U10120 ( .A0(n3005), .A1(n1027), .B0(n1026), .Y(n16454) );
  AOI21X1 U10121 ( .A0(n2702), .A1(n957), .B0(n956), .Y(n18029) );
  AOI21X1 U10122 ( .A0(n3365), .A1(n1111), .B0(n1110), .Y(n14564) );
  AOI21X1 U10123 ( .A0(n3070), .A1(n1041), .B0(n1040), .Y(n16139) );
  AOI21X1 U10124 ( .A0(n2762), .A1(n971), .B0(n970), .Y(n17714) );
  AOI21X1 U10125 ( .A0(n3425), .A1(n1125), .B0(n1124), .Y(n14249) );
  AOI21X1 U10126 ( .A0(n3124), .A1(n1055), .B0(n1054), .Y(n15824) );
  AOI21X1 U10127 ( .A0(n2830), .A1(n985), .B0(n984), .Y(n17399) );
  INVX1 U10128 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n76), .Y(n6144) );
  INVX1 U10129 ( .A(n8141), .Y(n5820) );
  INVX1 U10130 ( .A(n9893), .Y(n5348) );
  INVX1 U10131 ( .A(n11061), .Y(n4994) );
  INVX1 U10132 ( .A(n10769), .Y(n5078) );
  INVX1 U10133 ( .A(n9017), .Y(n5584) );
  INVX1 U10134 ( .A(n7265), .Y(n6048) );
  INVX1 U10135 ( .A(n10185), .Y(n5264) );
  INVX1 U10136 ( .A(n9309), .Y(n5508) );
  INVX1 U10137 ( .A(n8433), .Y(n5736) );
  INVX1 U10138 ( .A(n7557), .Y(n5972) );
  INVX1 U10139 ( .A(n11353), .Y(n4878) );
  INVX1 U10140 ( .A(n10477), .Y(n5186) );
  INVX1 U10141 ( .A(n9601), .Y(n5432) );
  INVX1 U10142 ( .A(n8725), .Y(n5660) );
  INVX1 U10143 ( .A(n7849), .Y(n5896) );
  OAI211X1 U10144 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n107), .A1(n3454), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n108), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n109), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n92) );
  AOI211X1 U10145 ( .A0(n6165), .A1(n466), .B0(n6163), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n114), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n107) );
  AOI22X1 U10146 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n110), .A1(n3452), 
        .B0(n723), .B1(n6119), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n109) );
  INVX1 U10147 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n115), .Y(n6163) );
  OAI211X1 U10148 ( .A0(n9922), .A1(n2853), .B0(n9923), .C0(n9924), .Y(n9908)
         );
  AOI211X1 U10149 ( .A0(n5375), .A1(n465), .B0(n5373), .C0(n9929), .Y(n9922)
         );
  AOI22X1 U10150 ( .A0(n9925), .A1(n2851), .B0(n722), .B1(n5333), .Y(n9924) );
  INVX1 U10151 ( .A(n9930), .Y(n5373) );
  OAI211X1 U10152 ( .A0(n11090), .A1(n2611), .B0(n11091), .C0(n11092), .Y(
        n11076) );
  AOI211X1 U10153 ( .A0(n5021), .A1(n467), .B0(n5019), .C0(n11097), .Y(n11090)
         );
  AOI22X1 U10154 ( .A0(n11093), .A1(n2609), .B0(n724), .B1(n4979), .Y(n11092)
         );
  INVX1 U10155 ( .A(n11098), .Y(n5019) );
  OAI211X1 U10156 ( .A0(n8170), .A1(n3213), .B0(n8171), .C0(n8172), .Y(n8156)
         );
  AOI211X1 U10157 ( .A0(n5847), .A1(n468), .B0(n5845), .C0(n8177), .Y(n8170)
         );
  AOI22X1 U10158 ( .A0(n8173), .A1(n3211), .B0(n725), .B1(n5805), .Y(n8172) );
  INVX1 U10159 ( .A(n8178), .Y(n5845) );
  OAI211X1 U10160 ( .A0(n10798), .A1(n2672), .B0(n10799), .C0(n10800), .Y(
        n10784) );
  AOI211X1 U10161 ( .A0(n5105), .A1(n474), .B0(n5103), .C0(n10805), .Y(n10798)
         );
  AOI22X1 U10162 ( .A0(n10801), .A1(n2670), .B0(n731), .B1(n5063), .Y(n10800)
         );
  INVX1 U10163 ( .A(n10806), .Y(n5103) );
  OAI211X1 U10164 ( .A0(n9046), .A1(n3033), .B0(n9047), .C0(n9048), .Y(n9032)
         );
  AOI211X1 U10165 ( .A0(n5611), .A1(n476), .B0(n5609), .C0(n9053), .Y(n9046)
         );
  AOI22X1 U10166 ( .A0(n9049), .A1(n3031), .B0(n733), .B1(n5569), .Y(n9048) );
  INVX1 U10167 ( .A(n9054), .Y(n5609) );
  OAI211X1 U10168 ( .A0(n7294), .A1(n3393), .B0(n7295), .C0(n7296), .Y(n7280)
         );
  AOI211X1 U10169 ( .A0(n6075), .A1(n478), .B0(n6073), .C0(n7301), .Y(n7294)
         );
  AOI22X1 U10170 ( .A0(n7297), .A1(n3391), .B0(n735), .B1(n6033), .Y(n7296) );
  INVX1 U10171 ( .A(n7302), .Y(n6073) );
  OAI211X1 U10172 ( .A0(n10214), .A1(n2793), .B0(n10215), .C0(n10216), .Y(
        n10200) );
  AOI211X1 U10173 ( .A0(n5291), .A1(n480), .B0(n5289), .C0(n10221), .Y(n10214)
         );
  AOI22X1 U10174 ( .A0(n10217), .A1(n2791), .B0(n737), .B1(n5249), .Y(n10216)
         );
  INVX1 U10175 ( .A(n10222), .Y(n5289) );
  OAI211X1 U10176 ( .A0(n9338), .A1(n2975), .B0(n9339), .C0(n9340), .Y(n9324)
         );
  AOI211X1 U10177 ( .A0(n5535), .A1(n473), .B0(n5533), .C0(n9345), .Y(n9338)
         );
  AOI22X1 U10178 ( .A0(n9341), .A1(n2973), .B0(n730), .B1(n5493), .Y(n9340) );
  INVX1 U10179 ( .A(n9346), .Y(n5533) );
  OAI211X1 U10180 ( .A0(n8462), .A1(n3152), .B0(n8463), .C0(n8464), .Y(n8448)
         );
  AOI211X1 U10181 ( .A0(n5763), .A1(n469), .B0(n5761), .C0(n8469), .Y(n8462)
         );
  AOI22X1 U10182 ( .A0(n8465), .A1(n3150), .B0(n726), .B1(n5721), .Y(n8464) );
  INVX1 U10183 ( .A(n8470), .Y(n5761) );
  OAI211X1 U10184 ( .A0(n7586), .A1(n3335), .B0(n7587), .C0(n7588), .Y(n7572)
         );
  AOI211X1 U10185 ( .A0(n5999), .A1(n475), .B0(n5997), .C0(n7593), .Y(n7586)
         );
  AOI22X1 U10186 ( .A0(n7589), .A1(n3333), .B0(n732), .B1(n5957), .Y(n7588) );
  INVX1 U10187 ( .A(n7594), .Y(n5997) );
  OAI211X1 U10188 ( .A0(n11382), .A1(n2550), .B0(n11383), .C0(n11384), .Y(
        n11368) );
  AOI211X1 U10189 ( .A0(n4905), .A1(n471), .B0(n4903), .C0(n11389), .Y(n11382)
         );
  AOI22X1 U10190 ( .A0(n11385), .A1(n2548), .B0(n728), .B1(n4863), .Y(n11384)
         );
  INVX1 U10191 ( .A(n11390), .Y(n4903) );
  OAI211X1 U10192 ( .A0(n10506), .A1(n2732), .B0(n10507), .C0(n10508), .Y(
        n10492) );
  AOI211X1 U10193 ( .A0(n5213), .A1(n477), .B0(n5211), .C0(n10513), .Y(n10506)
         );
  AOI22X1 U10194 ( .A0(n10509), .A1(n2730), .B0(n734), .B1(n5171), .Y(n10508)
         );
  INVX1 U10195 ( .A(n10514), .Y(n5211) );
  OAI211X1 U10196 ( .A0(n9630), .A1(n2914), .B0(n9631), .C0(n9632), .Y(n9616)
         );
  AOI211X1 U10197 ( .A0(n5459), .A1(n470), .B0(n5457), .C0(n9637), .Y(n9630)
         );
  AOI22X1 U10198 ( .A0(n9633), .A1(n2912), .B0(n727), .B1(n5417), .Y(n9632) );
  INVX1 U10199 ( .A(n9638), .Y(n5457) );
  OAI211X1 U10200 ( .A0(n8754), .A1(n3094), .B0(n8755), .C0(n8756), .Y(n8740)
         );
  AOI211X1 U10201 ( .A0(n5687), .A1(n479), .B0(n5685), .C0(n8761), .Y(n8754)
         );
  AOI22X1 U10202 ( .A0(n8757), .A1(n3092), .B0(n736), .B1(n5645), .Y(n8756) );
  INVX1 U10203 ( .A(n8762), .Y(n5685) );
  OAI211X1 U10204 ( .A0(n7878), .A1(n3274), .B0(n7879), .C0(n7880), .Y(n7864)
         );
  AOI211X1 U10205 ( .A0(n5923), .A1(n472), .B0(n5921), .C0(n7885), .Y(n7878)
         );
  AOI22X1 U10206 ( .A0(n7881), .A1(n3272), .B0(n729), .B1(n5881), .Y(n7880) );
  INVX1 U10207 ( .A(n7886), .Y(n5921) );
  OAI211XL U10208 ( .A0(n17007), .A1(n106), .B0(n17042), .C0(n17004), .Y(
        n17106) );
  OAI211XL U10209 ( .A0(n13857), .A1(n107), .B0(n13892), .C0(n13854), .Y(
        n13956) );
  OAI211XL U10210 ( .A0(n18267), .A1(n108), .B0(n18302), .C0(n18264), .Y(
        n18366) );
  OAI211XL U10211 ( .A0(n15117), .A1(n109), .B0(n15152), .C0(n15114), .Y(
        n15216) );
  OAI211XL U10212 ( .A0(n15432), .A1(n110), .B0(n15467), .C0(n15429), .Y(
        n15531) );
  OAI211XL U10213 ( .A0(n18582), .A1(n111), .B0(n18617), .C0(n18579), .Y(
        n18681) );
  OAI211XL U10214 ( .A0(n16692), .A1(n112), .B0(n16727), .C0(n16689), .Y(
        n16791) );
  OAI211XL U10215 ( .A0(n14802), .A1(n113), .B0(n14837), .C0(n14799), .Y(
        n14901) );
  OAI211XL U10216 ( .A0(n16377), .A1(n114), .B0(n16412), .C0(n16374), .Y(
        n16476) );
  OAI211XL U10217 ( .A0(n17952), .A1(n115), .B0(n17987), .C0(n17949), .Y(
        n18051) );
  OAI211XL U10218 ( .A0(n14487), .A1(n116), .B0(n14522), .C0(n14484), .Y(
        n14586) );
  OAI211XL U10219 ( .A0(n16062), .A1(n117), .B0(n16097), .C0(n16059), .Y(
        n16161) );
  OAI211XL U10220 ( .A0(n17637), .A1(n118), .B0(n17672), .C0(n17634), .Y(
        n17736) );
  OAI211XL U10221 ( .A0(n14172), .A1(n119), .B0(n14207), .C0(n14169), .Y(
        n14271) );
  OAI211XL U10222 ( .A0(n15747), .A1(n120), .B0(n15782), .C0(n15744), .Y(
        n15846) );
  OAI211XL U10223 ( .A0(n17322), .A1(n121), .B0(n17357), .C0(n17319), .Y(
        n17421) );
  OAI211XL U10224 ( .A0(n1681), .A1(n3), .B0(n13311), .C0(n13440), .Y(n13456)
         );
  OAI211XL U10225 ( .A0(n1739), .A1(n4), .B0(n12681), .C0(n12810), .Y(n12826)
         );
  OAI211XL U10226 ( .A0(n1710), .A1(n5), .B0(n12996), .C0(n13125), .Y(n13141)
         );
  OAI211XL U10227 ( .A0(n17007), .A1(n30), .B0(n17045), .C0(n17233), .Y(n17228) );
  NOR3X1 U10228 ( .A(n2869), .B(n1005), .C(n17205), .Y(n17234) );
  OAI211XL U10229 ( .A0(n13857), .A1(n31), .B0(n13895), .C0(n14083), .Y(n14078) );
  NOR3X1 U10230 ( .A(n3469), .B(n1144), .C(n14055), .Y(n14084) );
  OAI211XL U10231 ( .A0(n15117), .A1(n33), .B0(n15155), .C0(n15343), .Y(n15338) );
  NOR3X1 U10232 ( .A(n3229), .B(n1089), .C(n15315), .Y(n15344) );
  OAI211XL U10233 ( .A0(n18267), .A1(n32), .B0(n18305), .C0(n18493), .Y(n18488) );
  NOR3X1 U10234 ( .A(n2627), .B(n949), .C(n18465), .Y(n18494) );
  OAI211XL U10235 ( .A0(n15432), .A1(n34), .B0(n15470), .C0(n15658), .Y(n15653) );
  NOR3X1 U10236 ( .A(n3168), .B(n1075), .C(n15630), .Y(n15659) );
  OAI211XL U10237 ( .A0(n16692), .A1(n36), .B0(n16730), .C0(n16918), .Y(n16913) );
  NOR3X1 U10238 ( .A(n2930), .B(n1019), .C(n16890), .Y(n16919) );
  OAI211XL U10239 ( .A0(n18582), .A1(n35), .B0(n18620), .C0(n18808), .Y(n18803) );
  NOR3X1 U10240 ( .A(n2566), .B(n935), .C(n18780), .Y(n18809) );
  OAI211XL U10241 ( .A0(n14802), .A1(n37), .B0(n14840), .C0(n15028), .Y(n15023) );
  NOR3X1 U10242 ( .A(n3290), .B(n1103), .C(n15000), .Y(n15029) );
  OAI211XL U10243 ( .A0(n16377), .A1(n38), .B0(n16415), .C0(n16603), .Y(n16598) );
  NOR3X1 U10244 ( .A(n2991), .B(n1033), .C(n16575), .Y(n16604) );
  OAI211XL U10245 ( .A0(n17952), .A1(n39), .B0(n17990), .C0(n18178), .Y(n18173) );
  NOR3X1 U10246 ( .A(n2687), .B(n963), .C(n18150), .Y(n18179) );
  OAI211XL U10247 ( .A0(n14487), .A1(n40), .B0(n14525), .C0(n14713), .Y(n14708) );
  NOR3X1 U10248 ( .A(n3351), .B(n1117), .C(n14685), .Y(n14714) );
  OAI211XL U10249 ( .A0(n16062), .A1(n41), .B0(n16100), .C0(n16288), .Y(n16283) );
  NOR3X1 U10250 ( .A(n3049), .B(n1047), .C(n16260), .Y(n16289) );
  OAI211XL U10251 ( .A0(n17637), .A1(n42), .B0(n17675), .C0(n17863), .Y(n17858) );
  NOR3X1 U10252 ( .A(n2748), .B(n977), .C(n17835), .Y(n17864) );
  OAI211XL U10253 ( .A0(n14172), .A1(n43), .B0(n14210), .C0(n14398), .Y(n14393) );
  NOR3X1 U10254 ( .A(n3409), .B(n1131), .C(n14370), .Y(n14399) );
  OAI211XL U10255 ( .A0(n15747), .A1(n44), .B0(n15785), .C0(n15973), .Y(n15968) );
  NOR3X1 U10256 ( .A(n3110), .B(n1061), .C(n15945), .Y(n15974) );
  OAI211XL U10257 ( .A0(n17322), .A1(n45), .B0(n17360), .C0(n17548), .Y(n17543) );
  NOR3X1 U10258 ( .A(n2809), .B(n991), .C(n17520), .Y(n17549) );
  NAND2X1 U10259 ( .A(n673), .B(n6915), .Y(n11680) );
  NAND2X1 U10260 ( .A(n674), .B(n6869), .Y(top_core_KE_sb1_n105) );
  NAND2X1 U10261 ( .A(n675), .B(n6622), .Y(n12311) );
  NAND2X1 U10262 ( .A(n677), .B(n6550), .Y(n13257) );
  NAND2X1 U10263 ( .A(n676), .B(n6575), .Y(n11996) );
  NAND2X1 U10264 ( .A(n678), .B(n6845), .Y(n12627) );
  NAND2X1 U10265 ( .A(n679), .B(n6598), .Y(n13572) );
  NAND2X1 U10266 ( .A(n680), .B(n6891), .Y(n12942) );
  NAND2X1 U10267 ( .A(n685), .B(n6597), .Y(n13664) );
  NAND2X1 U10268 ( .A(n995), .B(n2893), .Y(n17130) );
  NAND2X1 U10269 ( .A(n1134), .B(n3494), .Y(n13980) );
  NAND2X1 U10270 ( .A(n1079), .B(n3253), .Y(n15240) );
  NAND2X1 U10271 ( .A(n939), .B(n2650), .Y(n18390) );
  NAND2X1 U10272 ( .A(n1065), .B(n3192), .Y(n15555) );
  NAND2X1 U10273 ( .A(n1009), .B(n2954), .Y(n16815) );
  NAND2X1 U10274 ( .A(n925), .B(top_core_EC_ss_in[120]), .Y(n18705) );
  NAND2X1 U10275 ( .A(n1093), .B(n3314), .Y(n14925) );
  NAND2X1 U10276 ( .A(n1023), .B(n3015), .Y(n16500) );
  NAND2X1 U10277 ( .A(n953), .B(n2711), .Y(n18075) );
  NAND2X1 U10278 ( .A(n1107), .B(n3375), .Y(n14610) );
  NAND2X1 U10279 ( .A(n1037), .B(n3072), .Y(n16185) );
  NAND2X1 U10280 ( .A(n967), .B(n2772), .Y(n17760) );
  NAND2X1 U10281 ( .A(n1121), .B(n3433), .Y(n14295) );
  NAND2X1 U10282 ( .A(n1051), .B(n3134), .Y(n15870) );
  NAND2X1 U10283 ( .A(n981), .B(n2833), .Y(n17445) );
  NAND2X1 U10284 ( .A(n1134), .B(n3486), .Y(n13878) );
  NAND2X1 U10285 ( .A(n995), .B(n2891), .Y(n17028) );
  NAND2X1 U10286 ( .A(n939), .B(n2649), .Y(n18288) );
  NAND2X1 U10287 ( .A(n1079), .B(n3251), .Y(n15138) );
  NAND2X1 U10288 ( .A(n1065), .B(n3184), .Y(n15453) );
  NAND2X1 U10289 ( .A(n925), .B(n2582), .Y(n18603) );
  NAND2X1 U10290 ( .A(n1009), .B(n2952), .Y(n16713) );
  NAND2X1 U10291 ( .A(n1093), .B(n3312), .Y(n14823) );
  NAND2X1 U10292 ( .A(n1023), .B(n3013), .Y(n16398) );
  NAND2X1 U10293 ( .A(n953), .B(n2704), .Y(n17973) );
  NAND2X1 U10294 ( .A(n1107), .B(n3367), .Y(n14508) );
  NAND2X1 U10295 ( .A(n1037), .B(n3071), .Y(n16083) );
  NAND2X1 U10296 ( .A(n967), .B(n2764), .Y(n17658) );
  NAND2X1 U10297 ( .A(n1121), .B(n3431), .Y(n14193) );
  NAND2X1 U10298 ( .A(n1051), .B(n3126), .Y(n15768) );
  NAND2X1 U10299 ( .A(n981), .B(n2831), .Y(n17343) );
  NOR4BBX1 U10300 ( .AN(n17131), .BN(n17132), .C(n17009), .D(n16999), .Y(
        n17102) );
  AOI222X1 U10301 ( .A0(n2863), .A1(n17133), .B0(n17134), .B1(n2865), .C0(n386), .C1(n5328), .Y(n17132) );
  OAI21XL U10302 ( .A0(n17135), .A1(n1310), .B0(n17046), .Y(n17134) );
  NOR4BBX1 U10303 ( .AN(n13981), .BN(n13982), .C(n13859), .D(n13849), .Y(
        n13952) );
  AOI222X1 U10304 ( .A0(n3460), .A1(n13983), .B0(n13984), .B1(n3466), .C0(n385), .C1(n6112), .Y(n13982) );
  OAI21XL U10305 ( .A0(n13985), .A1(n1280), .B0(n13896), .Y(n13984) );
  NOR4BBX1 U10306 ( .AN(n18391), .BN(n18392), .C(n18269), .D(n18259), .Y(
        n18362) );
  AOI222X1 U10307 ( .A0(n2620), .A1(n18393), .B0(n18394), .B1(n2609), .C0(n387), .C1(n4974), .Y(n18392) );
  OAI21XL U10308 ( .A0(n18395), .A1(n1322), .B0(n18306), .Y(n18394) );
  NOR4BBX1 U10309 ( .AN(n15241), .BN(n15242), .C(n15119), .D(n15109), .Y(
        n15212) );
  AOI222X1 U10310 ( .A0(n3223), .A1(n15243), .B0(n15244), .B1(n3225), .C0(n388), .C1(n5800), .Y(n15242) );
  OAI21XL U10311 ( .A0(n15245), .A1(n1292), .B0(n15156), .Y(n15244) );
  NOR4BBX1 U10312 ( .AN(n15556), .BN(n15557), .C(n15434), .D(n15424), .Y(
        n15527) );
  AOI222X1 U10313 ( .A0(n3161), .A1(n15558), .B0(n15559), .B1(n3164), .C0(n389), .C1(n5716), .Y(n15557) );
  OAI21XL U10314 ( .A0(n15560), .A1(n1295), .B0(n15471), .Y(n15559) );
  NOR4BBX1 U10315 ( .AN(n18706), .BN(n18707), .C(n18584), .D(n18574), .Y(
        n18677) );
  AOI222X1 U10316 ( .A0(n2558), .A1(n18708), .B0(n18709), .B1(n2562), .C0(n390), .C1(n4858), .Y(n18707) );
  OAI21XL U10317 ( .A0(n18710), .A1(n1325), .B0(n18621), .Y(n18709) );
  NOR4BBX1 U10318 ( .AN(n16816), .BN(n16817), .C(n16694), .D(n16684), .Y(
        n16787) );
  AOI222X1 U10319 ( .A0(n2923), .A1(n16818), .B0(n16819), .B1(n2926), .C0(n391), .C1(n5412), .Y(n16817) );
  OAI21XL U10320 ( .A0(n16820), .A1(n1307), .B0(n16731), .Y(n16819) );
  NOR4BBX1 U10321 ( .AN(n14926), .BN(n14927), .C(n14804), .D(n14794), .Y(
        n14897) );
  AOI222X1 U10322 ( .A0(n3283), .A1(n14928), .B0(n14929), .B1(n3286), .C0(n392), .C1(n5876), .Y(n14927) );
  OAI21XL U10323 ( .A0(n14930), .A1(n1289), .B0(n14841), .Y(n14929) );
  NOR4BBX1 U10324 ( .AN(n16501), .BN(n16502), .C(n16379), .D(n16369), .Y(
        n16472) );
  AOI222X1 U10325 ( .A0(n2984), .A1(n16503), .B0(n16504), .B1(n2987), .C0(n393), .C1(n5488), .Y(n16502) );
  OAI21XL U10326 ( .A0(n16505), .A1(n1304), .B0(n16416), .Y(n16504) );
  NOR4BBX1 U10327 ( .AN(n18076), .BN(n18077), .C(n17954), .D(n17944), .Y(
        n18047) );
  AOI222X1 U10328 ( .A0(n2682), .A1(n18078), .B0(n18079), .B1(n2684), .C0(n394), .C1(n5058), .Y(n18077) );
  OAI21XL U10329 ( .A0(n18080), .A1(n1319), .B0(n17991), .Y(n18079) );
  NOR4BBX1 U10330 ( .AN(n14611), .BN(n14612), .C(n14489), .D(n14479), .Y(
        n14582) );
  AOI222X1 U10331 ( .A0(n3344), .A1(n14613), .B0(n14614), .B1(n3333), .C0(n395), .C1(n5952), .Y(n14612) );
  OAI21XL U10332 ( .A0(n14615), .A1(n1286), .B0(n14526), .Y(n14614) );
  NOR4BBX1 U10333 ( .AN(n16186), .BN(n16187), .C(n16064), .D(n16054), .Y(
        n16157) );
  AOI222X1 U10334 ( .A0(n3042), .A1(n16188), .B0(n16189), .B1(n3031), .C0(n396), .C1(n5564), .Y(n16187) );
  OAI21XL U10335 ( .A0(n16190), .A1(n1301), .B0(n16101), .Y(n16189) );
  NOR4BBX1 U10336 ( .AN(n17761), .BN(n17762), .C(n17639), .D(n17629), .Y(
        n17732) );
  AOI222X1 U10337 ( .A0(n2742), .A1(n17763), .B0(n17764), .B1(n2744), .C0(n397), .C1(n5166), .Y(n17762) );
  OAI21XL U10338 ( .A0(n17765), .A1(n1316), .B0(n17676), .Y(n17764) );
  NOR4BBX1 U10339 ( .AN(n14296), .BN(n14297), .C(n14174), .D(n14164), .Y(
        n14267) );
  AOI222X1 U10340 ( .A0(n3402), .A1(n14298), .B0(n14299), .B1(n3391), .C0(n398), .C1(n6028), .Y(n14297) );
  OAI21XL U10341 ( .A0(n14300), .A1(n1283), .B0(n14211), .Y(n14299) );
  NOR4BBX1 U10342 ( .AN(n15871), .BN(n15872), .C(n15749), .D(n15739), .Y(
        n15842) );
  AOI222X1 U10343 ( .A0(n3104), .A1(n15873), .B0(n15874), .B1(n3106), .C0(n399), .C1(n5640), .Y(n15872) );
  OAI21XL U10344 ( .A0(n15875), .A1(n1298), .B0(n15786), .Y(n15874) );
  NOR4BBX1 U10345 ( .AN(n17446), .BN(n17447), .C(n17324), .D(n17314), .Y(
        n17417) );
  AOI222X1 U10346 ( .A0(n2802), .A1(n17448), .B0(n17449), .B1(n2805), .C0(n400), .C1(n5244), .Y(n17447) );
  OAI21XL U10347 ( .A0(n17450), .A1(n1313), .B0(n17361), .Y(n17449) );
  NAND2X1 U10348 ( .A(n5330), .B(n999), .Y(n17275) );
  NAND2X1 U10349 ( .A(n6114), .B(n1138), .Y(n14125) );
  NAND2X1 U10350 ( .A(n5802), .B(n1083), .Y(n15385) );
  NAND2X1 U10351 ( .A(n4976), .B(n943), .Y(n18535) );
  NAND2X1 U10352 ( .A(n5718), .B(n1069), .Y(n15700) );
  NAND2X1 U10353 ( .A(n5414), .B(n1013), .Y(n16960) );
  NAND2X1 U10354 ( .A(n4860), .B(n929), .Y(n18850) );
  NAND2X1 U10355 ( .A(n5878), .B(n1097), .Y(n15070) );
  NAND2X1 U10356 ( .A(n5490), .B(n1027), .Y(n16645) );
  NAND2X1 U10357 ( .A(n5060), .B(n957), .Y(n18220) );
  NAND2X1 U10358 ( .A(n5954), .B(n1111), .Y(n14755) );
  NAND2X1 U10359 ( .A(n5566), .B(n1041), .Y(n16330) );
  NAND2X1 U10360 ( .A(n5168), .B(n971), .Y(n17905) );
  NAND2X1 U10361 ( .A(n6030), .B(n1125), .Y(n14440) );
  NAND2X1 U10362 ( .A(n5642), .B(n1055), .Y(n16015) );
  NAND2X1 U10363 ( .A(n5246), .B(n985), .Y(n17590) );
  NOR4X1 U10364 ( .A(n13242), .B(n13243), .C(n13244), .D(n13245), .Y(n13208)
         );
  OAI21XL U10365 ( .A0(n1680), .A1(n13252), .B0(n13253), .Y(n13243) );
  AOI31X1 U10366 ( .A0(n13249), .A1(n13250), .A2(n13227), .B0(n13251), .Y(
        n13244) );
  NAND2X1 U10367 ( .A(n1157), .B(n1180), .Y(n13540) );
  NAND2X1 U10368 ( .A(n1180), .B(n6597), .Y(n13563) );
  NAND3XL U10369 ( .A(n9970), .B(n2872), .C(n17126), .Y(n17240) );
  NAND3XL U10370 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .B(n3473), .C(
        n13976), .Y(n14090) );
  NAND3XL U10371 ( .A(n8218), .B(n3232), .C(n15236), .Y(n15350) );
  NAND3XL U10372 ( .A(n11138), .B(n2630), .C(n18386), .Y(n18500) );
  NAND3XL U10373 ( .A(n8510), .B(n3171), .C(n15551), .Y(n15665) );
  NAND3XL U10374 ( .A(n9678), .B(n2933), .C(n16811), .Y(n16925) );
  NAND3XL U10375 ( .A(n11430), .B(n2569), .C(n18701), .Y(n18815) );
  NAND3XL U10376 ( .A(n7926), .B(n3293), .C(n14921), .Y(n15035) );
  NAND3XL U10377 ( .A(n9386), .B(n2994), .C(n16496), .Y(n16610) );
  NAND3XL U10378 ( .A(n10846), .B(n2691), .C(n18071), .Y(n18185) );
  NAND3XL U10379 ( .A(n7634), .B(n3354), .C(n14606), .Y(n14720) );
  NAND3XL U10380 ( .A(n9094), .B(n3052), .C(n16181), .Y(n16295) );
  NAND3XL U10381 ( .A(n10554), .B(n2751), .C(n17756), .Y(n17870) );
  NAND3XL U10382 ( .A(n7342), .B(n3412), .C(n14291), .Y(n14405) );
  NAND3XL U10383 ( .A(n8802), .B(n3113), .C(n15866), .Y(n15980) );
  NAND3XL U10384 ( .A(n10262), .B(n2812), .C(n17441), .Y(n17555) );
  AOI21XL U10385 ( .A0(n1274), .A1(n6549), .B0(n13455), .Y(n13266) );
  AOI21XL U10386 ( .A0(n1268), .A1(n6844), .B0(n12825), .Y(n12636) );
  AOI21XL U10387 ( .A0(n1277), .A1(n6597), .B0(n13770), .Y(n13581) );
  AOI21XL U10388 ( .A0(n1271), .A1(n6890), .B0(n13140), .Y(n12951) );
  NOR2XL U10389 ( .A(n73), .B(n1666), .Y(n13233) );
  NOR2XL U10390 ( .A(n75), .B(n1695), .Y(n12918) );
  NOR2XL U10391 ( .A(n74), .B(n1724), .Y(n12603) );
  INVX1 U10392 ( .A(n12626), .Y(n6780) );
  INVX1 U10393 ( .A(n12941), .Y(n6819) );
  INVX1 U10394 ( .A(n13256), .Y(n6477) );
  CLKINVX3 U10395 ( .A(n3947), .Y(n3714) );
  CLKINVX3 U10396 ( .A(n3947), .Y(n3712) );
  CLKINVX3 U10397 ( .A(n3929), .Y(n3711) );
  CLKINVX3 U10398 ( .A(n3908), .Y(n3710) );
  CLKINVX3 U10399 ( .A(n3930), .Y(n3709) );
  CLKINVX3 U10400 ( .A(n3947), .Y(n3713) );
  NOR2XL U10401 ( .A(n13223), .B(n1673), .Y(n13280) );
  NOR2XL U10402 ( .A(n12593), .B(n1731), .Y(n12650) );
  NOR2XL U10403 ( .A(n12908), .B(n1702), .Y(n12965) );
  CLKINVX3 U10404 ( .A(n3907), .Y(n3904) );
  CLKINVX3 U10405 ( .A(n3907), .Y(n3905) );
  XOR2X1 U10406 ( .A(top_core_EC_mc_mix_in_4_32_), .B(
        top_core_EC_mc_mix_in_2_34_), .Y(top_core_EC_mc_mix_in_4_35_) );
  XOR2X1 U10407 ( .A(top_core_EC_mc_mix_in_8[32]), .B(
        top_core_EC_mc_mix_in_8[48]), .Y(top_core_EC_mc_n329) );
  XOR2X1 U10408 ( .A(top_core_EC_mc_mix_in_4_32_), .B(
        top_core_EC_mc_mix_in_4_48_), .Y(top_core_EC_mc_n321) );
  XOR2X1 U10409 ( .A(top_core_EC_mc_mix_in_4_32_), .B(
        top_core_EC_mc_mix_in_2_32_), .Y(top_core_EC_mc_mix_in_8[34]) );
  XOR2X1 U10410 ( .A(top_core_EC_mc_mix_in_4_32_), .B(
        top_core_EC_mc_mix_in_2_35_), .Y(top_core_EC_mc_mix_in_8[37]) );
  XOR2X1 U10411 ( .A(top_core_EC_mc_mix_in_4_16_), .B(
        top_core_EC_mc_mix_in_2_18_), .Y(top_core_EC_mc_mix_in_4_19_) );
  CLKINVX3 U10412 ( .A(n11706), .Y(n6920) );
  CLKINVX3 U10413 ( .A(top_core_KE_sb1_n131), .Y(n6874) );
  CLKINVX3 U10414 ( .A(n12022), .Y(n6580) );
  CLKINVX3 U10415 ( .A(n13283), .Y(n6556) );
  CLKINVX3 U10416 ( .A(n12968), .Y(n6897) );
  CLKINVX3 U10417 ( .A(n13598), .Y(n6604) );
  CLKINVX3 U10418 ( .A(n12653), .Y(n6851) );
  XOR2X1 U10419 ( .A(top_core_EC_mc_mix_in_2_0_), .B(top_core_EC_mix_in[2]), 
        .Y(top_core_EC_mc_mix_in_2_3_) );
  XOR2X1 U10420 ( .A(top_core_EC_mc_mix_in_2_48_), .B(top_core_EC_mix_in[50]), 
        .Y(top_core_EC_mc_mix_in_2_51_) );
  XOR2X1 U10421 ( .A(top_core_EC_mc_mix_in_8[15]), .B(
        top_core_EC_mc_mix_in_8[6]), .Y(top_core_EC_mc_n435) );
  XOR2X1 U10422 ( .A(top_core_EC_mc_mix_in_2_16_), .B(top_core_EC_mix_in[18]), 
        .Y(top_core_EC_mc_mix_in_2_19_) );
  XOR2X1 U10423 ( .A(top_core_EC_mc_mix_in_2_32_), .B(top_core_EC_mix_in[34]), 
        .Y(top_core_EC_mc_mix_in_2_35_) );
  XOR2X1 U10424 ( .A(top_core_EC_mc_mix_in_2_32_), .B(
        top_core_EC_mc_mix_in_2_48_), .Y(top_core_EC_mc_n313) );
  XOR2X1 U10425 ( .A(top_core_EC_mc_mix_in_2_26_), .B(
        top_core_EC_mc_mix_in_4_18_), .Y(top_core_EC_mc_n10) );
  XOR2X1 U10426 ( .A(n1548), .B(top_core_EC_mc_mix_in_4_0_), .Y(
        top_core_EC_mc_n192) );
  XOR2X1 U10427 ( .A(n1549), .B(top_core_EC_mc_mix_in_8[0]), .Y(
        top_core_EC_mc_n257) );
  XOR2X1 U10428 ( .A(top_core_EC_mc_mix_in_8[39]), .B(
        top_core_EC_mc_mix_in_8[55]), .Y(top_core_EC_mc_n337) );
  XOR2X1 U10429 ( .A(top_core_EC_mix_in[24]), .B(top_core_EC_mc_mix_in_2_16_), 
        .Y(top_core_EC_mc_n103) );
  XOR2X1 U10430 ( .A(top_core_EC_mc_mix_in_2_34_), .B(
        top_core_EC_mc_mix_in_2_50_), .Y(top_core_EC_mc_n370) );
  XOR2X1 U10431 ( .A(n1549), .B(top_core_EC_mc_mix_in_2_10_), .Y(
        top_core_EC_mc_mix_in_4_11_) );
  XOR2X1 U10432 ( .A(n1543), .B(top_core_EC_mc_mix_in_2_42_), .Y(
        top_core_EC_mc_mix_in_4_43_) );
  XOR2X1 U10433 ( .A(top_core_EC_mix_in[32]), .B(top_core_EC_mix_in[48]), .Y(
        top_core_EC_mc_n378) );
  XOR2X1 U10434 ( .A(top_core_EC_mix_in[34]), .B(top_core_EC_mix_in[50]), .Y(
        top_core_EC_mc_n362) );
  XOR2X1 U10435 ( .A(top_core_EC_mix_in[35]), .B(top_core_EC_mix_in[51]), .Y(
        top_core_EC_mc_n354) );
  NAND2X1 U10436 ( .A(n1001), .B(n722), .Y(n10079) );
  NAND2X1 U10437 ( .A(n1143), .B(n723), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n265) );
  NAND2X1 U10438 ( .A(n945), .B(n724), .Y(n11247) );
  NAND2X1 U10439 ( .A(n1085), .B(n725), .Y(n8327) );
  NAND2X1 U10440 ( .A(n959), .B(n731), .Y(n10955) );
  NAND2X1 U10441 ( .A(n1127), .B(n735), .Y(n7451) );
  NAND2X1 U10442 ( .A(n1043), .B(n733), .Y(n9203) );
  NAND2X1 U10443 ( .A(n987), .B(n737), .Y(n10371) );
  NAND2X1 U10444 ( .A(n1029), .B(n730), .Y(n9495) );
  NAND2X1 U10445 ( .A(n1071), .B(n726), .Y(n8619) );
  NAND2X1 U10446 ( .A(n1113), .B(n732), .Y(n7743) );
  NAND2X1 U10447 ( .A(n931), .B(n728), .Y(n11539) );
  NAND2X1 U10448 ( .A(n973), .B(n734), .Y(n10663) );
  NAND2X1 U10449 ( .A(n1015), .B(n727), .Y(n9787) );
  NAND2X1 U10450 ( .A(n1057), .B(n736), .Y(n8911) );
  NAND2X1 U10451 ( .A(n1099), .B(n729), .Y(n8035) );
  XOR2X1 U10452 ( .A(top_core_EC_mix_in[10]), .B(top_core_EC_mc_mix_in_2_2_), 
        .Y(top_core_EC_mc_n587) );
  XOR2X1 U10453 ( .A(top_core_EC_mix_in[11]), .B(top_core_EC_mc_mix_in_2_3_), 
        .Y(top_core_EC_mc_n500) );
  XOR2X1 U10454 ( .A(n1550), .B(top_core_EC_mc_mix_in_8[7]), .Y(
        top_core_EC_mc_n346) );
  XOR2X1 U10455 ( .A(top_core_EC_mc_n410), .B(top_core_EC_mc_n337), .Y(
        top_core_EC_mc_n471) );
  XOR2X1 U10456 ( .A(top_core_EC_mc_n175), .B(top_core_EC_mc_n111), .Y(
        top_core_EC_mc_n227) );
  XOR2X1 U10457 ( .A(top_core_EC_mc_n151), .B(top_core_EC_mc_n78), .Y(
        top_core_EC_mc_n212) );
  XOR2X1 U10458 ( .A(top_core_EC_mc_n828), .B(top_core_EC_mc_n764), .Y(
        top_core_EC_mc_n880) );
  XOR2X1 U10459 ( .A(top_core_EC_mc_n810), .B(top_core_EC_mc_n743), .Y(
        top_core_EC_mc_n861) );
  XOR2X1 U10460 ( .A(top_core_EC_mc_n394), .B(top_core_EC_mc_n321), .Y(
        top_core_EC_mc_n461) );
  XOR2X1 U10461 ( .A(top_core_EC_mc_n386), .B(top_core_EC_mc_n313), .Y(
        top_core_EC_mc_n456) );
  XOR2X1 U10462 ( .A(top_core_EC_mc_n135), .B(top_core_EC_mc_n62), .Y(
        top_core_EC_mc_n202) );
  XOR2X1 U10463 ( .A(top_core_EC_mc_n127), .B(top_core_EC_mc_n54), .Y(
        top_core_EC_mc_n197) );
  XOR2X1 U10464 ( .A(top_core_EC_mc_n794), .B(top_core_EC_mc_n727), .Y(
        top_core_EC_mc_n844) );
  XOR2X1 U10465 ( .A(top_core_EC_mc_n786), .B(top_core_EC_mc_n719), .Y(
        top_core_EC_mc_n839) );
  XOR2X1 U10466 ( .A(top_core_EC_mc_n426), .B(top_core_EC_mc_n362), .Y(
        top_core_EC_mc_n481) );
  XOR2X1 U10467 ( .A(top_core_EC_mc_n418), .B(top_core_EC_mc_n354), .Y(
        top_core_EC_mc_n476) );
  XOR2X1 U10468 ( .A(top_core_EC_mc_n183), .B(top_core_EC_mc_n119), .Y(
        top_core_EC_mc_n232) );
  XOR2X1 U10469 ( .A(top_core_EC_mc_n402), .B(top_core_EC_mc_n329), .Y(
        top_core_EC_mc_n466) );
  XOR2X1 U10470 ( .A(top_core_EC_mc_n167), .B(top_core_EC_mc_n94), .Y(
        top_core_EC_mc_n222) );
  XOR2X1 U10471 ( .A(top_core_EC_mc_n159), .B(top_core_EC_mc_n86), .Y(
        top_core_EC_mc_n217) );
  XOR2X1 U10472 ( .A(top_core_EC_mc_n834), .B(top_core_EC_mc_n771), .Y(
        top_core_EC_mc_n887) );
  XOR2X1 U10473 ( .A(top_core_EC_mc_n143), .B(top_core_EC_mc_n70), .Y(
        top_core_EC_mc_n207) );
  XOR2X1 U10474 ( .A(top_core_EC_mc_n822), .B(top_core_EC_mc_n757), .Y(
        top_core_EC_mc_n873) );
  XOR2X1 U10475 ( .A(top_core_EC_mc_n816), .B(top_core_EC_mc_n750), .Y(
        top_core_EC_mc_n866) );
  XOR2X1 U10476 ( .A(top_core_EC_mc_n802), .B(top_core_EC_mc_n735), .Y(
        top_core_EC_mc_n856) );
  XNOR2X1 U10477 ( .A(top_core_EC_mc_n929), .B(top_core_EC_mc_n627), .Y(
        top_core_EC_mc_n926) );
  XNOR2X1 U10478 ( .A(top_core_EC_mix_in[16]), .B(n1548), .Y(
        top_core_EC_mc_n929) );
  XNOR2X1 U10479 ( .A(top_core_EC_mc_n677), .B(top_core_EC_mc_n10), .Y(
        top_core_EC_mc_n674) );
  XNOR2X1 U10480 ( .A(top_core_EC_mc_mix_in_2_2_), .B(
        top_core_EC_mc_mix_in_2_10_), .Y(top_core_EC_mc_n677) );
  XNOR2X1 U10481 ( .A(top_core_EC_mc_n669), .B(top_core_EC_mc_n670), .Y(
        top_core_EC_mc_n668) );
  XNOR2X1 U10482 ( .A(top_core_EC_mix_in[10]), .B(top_core_EC_mix_in[2]), .Y(
        top_core_EC_mc_n669) );
  XNOR2X1 U10483 ( .A(top_core_EC_mc_n663), .B(top_core_EC_mc_n664), .Y(
        top_core_EC_mc_n662) );
  XNOR2X1 U10484 ( .A(top_core_EC_mix_in[11]), .B(top_core_EC_mix_in[3]), .Y(
        top_core_EC_mc_n663) );
  XNOR2X1 U10485 ( .A(top_core_EC_mc_n650), .B(top_core_EC_mc_n651), .Y(
        top_core_EC_mc_n649) );
  XNOR2X1 U10486 ( .A(top_core_EC_mc_mix_in_8[15]), .B(
        top_core_EC_mc_mix_in_8[7]), .Y(top_core_EC_mc_n650) );
  XNOR2X1 U10487 ( .A(top_core_EC_mc_n644), .B(top_core_EC_mc_n645), .Y(
        top_core_EC_mc_n643) );
  XNOR2X1 U10488 ( .A(n1550), .B(top_core_EC_mc_mix_in_8[0]), .Y(
        top_core_EC_mc_n644) );
  XNOR2X1 U10489 ( .A(top_core_EC_mc_n638), .B(top_core_EC_mc_n639), .Y(
        top_core_EC_mc_n637) );
  XNOR2X1 U10490 ( .A(n1549), .B(top_core_EC_mc_mix_in_4_0_), .Y(
        top_core_EC_mc_n638) );
  XNOR2X1 U10491 ( .A(top_core_EC_mc_n632), .B(top_core_EC_mc_n633), .Y(
        top_core_EC_mc_n631) );
  XNOR2X1 U10492 ( .A(n1548), .B(top_core_EC_mc_mix_in_2_0_), .Y(
        top_core_EC_mc_n632) );
  XNOR2X1 U10493 ( .A(top_core_EC_mc_n564), .B(top_core_EC_mc_n377), .Y(
        top_core_EC_mc_n561) );
  XNOR2X1 U10494 ( .A(top_core_EC_mix_in[48]), .B(n1542), .Y(
        top_core_EC_mc_n564) );
  XNOR2X1 U10495 ( .A(top_core_EC_mc_n556), .B(top_core_EC_mc_n369), .Y(
        top_core_EC_mc_n553) );
  XNOR2X1 U10496 ( .A(top_core_EC_mc_mix_in_2_50_), .B(
        top_core_EC_mc_mix_in_4_42_), .Y(top_core_EC_mc_n556) );
  XNOR2X1 U10497 ( .A(top_core_EC_mc_n548), .B(top_core_EC_mc_n361), .Y(
        top_core_EC_mc_n545) );
  XNOR2X1 U10498 ( .A(top_core_EC_mix_in[50]), .B(top_core_EC_mc_mix_in_2_42_), 
        .Y(top_core_EC_mc_n548) );
  XNOR2X1 U10499 ( .A(top_core_EC_mc_n540), .B(top_core_EC_mc_n353), .Y(
        top_core_EC_mc_n537) );
  XNOR2X1 U10500 ( .A(top_core_EC_mix_in[51]), .B(top_core_EC_mc_mix_in_2_43_), 
        .Y(top_core_EC_mc_n540) );
  XNOR2X1 U10501 ( .A(top_core_EC_mc_n532), .B(top_core_EC_mc_n336), .Y(
        top_core_EC_mc_n529) );
  XNOR2X1 U10502 ( .A(top_core_EC_mc_mix_in_8[55]), .B(
        top_core_EC_mc_mix_in_8[46]), .Y(top_core_EC_mc_n532) );
  XNOR2X1 U10503 ( .A(top_core_EC_mc_n524), .B(top_core_EC_mc_n328), .Y(
        top_core_EC_mc_n521) );
  XNOR2X1 U10504 ( .A(top_core_EC_mc_mix_in_8[48]), .B(
        top_core_EC_mc_mix_in_8[47]), .Y(top_core_EC_mc_n524) );
  XNOR2X1 U10505 ( .A(top_core_EC_mc_n516), .B(top_core_EC_mc_n320), .Y(
        top_core_EC_mc_n513) );
  XNOR2X1 U10506 ( .A(top_core_EC_mc_mix_in_4_48_), .B(n1544), .Y(
        top_core_EC_mc_n516) );
  XNOR2X1 U10507 ( .A(top_core_EC_mc_n508), .B(top_core_EC_mc_n312), .Y(
        top_core_EC_mc_n505) );
  XNOR2X1 U10508 ( .A(top_core_EC_mc_mix_in_2_48_), .B(n1543), .Y(
        top_core_EC_mc_n508) );
  XOR2X1 U10509 ( .A(n1546), .B(n1545), .Y(top_core_EC_mc_mix_in_8[26]) );
  XOR2X1 U10510 ( .A(n1549), .B(top_core_EC_mc_mix_in_2_11_), .Y(
        top_core_EC_mc_mix_in_8[13]) );
  XOR2X1 U10511 ( .A(top_core_EC_mc_mix_in_4_0_), .B(
        top_core_EC_mc_mix_in_2_2_), .Y(top_core_EC_mc_mix_in_4_3_) );
  XOR2X1 U10512 ( .A(top_core_EC_mc_mix_in_8[0]), .B(
        top_core_EC_mc_mix_in_8[16]), .Y(top_core_EC_mc_n189) );
  XOR2X1 U10513 ( .A(top_core_EC_mc_mix_in_4_48_), .B(
        top_core_EC_mc_mix_in_2_50_), .Y(top_core_EC_mc_mix_in_4_51_) );
  XOR2X1 U10514 ( .A(top_core_EC_mc_mix_in_4_48_), .B(
        top_core_EC_mc_mix_in_2_48_), .Y(top_core_EC_mc_mix_in_8[50]) );
  XOR2X1 U10515 ( .A(top_core_EC_mc_mix_in_4_48_), .B(
        top_core_EC_mc_mix_in_2_51_), .Y(top_core_EC_mc_mix_in_8[53]) );
  XOR2X1 U10516 ( .A(top_core_EC_mc_mix_in_4_48_), .B(
        top_core_EC_mc_mix_in_4_32_), .Y(top_core_EC_mc_n448) );
  XOR2X1 U10517 ( .A(top_core_EC_mc_mix_in_8[48]), .B(
        top_core_EC_mc_mix_in_8[32]), .Y(top_core_EC_mc_n383) );
  XOR2X1 U10518 ( .A(top_core_EC_mc_mix_in_4_16_), .B(
        top_core_EC_mc_mix_in_4_0_), .Y(top_core_EC_mc_n682) );
  XOR2X1 U10519 ( .A(top_core_EC_mc_mix_in_4_16_), .B(
        top_core_EC_mc_mix_in_4_0_), .Y(top_core_EC_mc_n578) );
  XOR2X1 U10520 ( .A(top_core_EC_mc_mix_in_8[16]), .B(
        top_core_EC_mc_mix_in_8[0]), .Y(top_core_EC_mc_n594) );
  XOR2X1 U10521 ( .A(top_core_EC_mc_mix_in_8[31]), .B(
        top_core_EC_mc_mix_in_8[15]), .Y(top_core_EC_mc_n577) );
  XOR2X1 U10522 ( .A(top_core_EC_mc_mix_in_8[31]), .B(
        top_core_EC_mc_mix_in_8[22]), .Y(top_core_EC_mc_n651) );
  XOR2X1 U10523 ( .A(top_core_EC_mc_mix_in_8[47]), .B(
        top_core_EC_mc_mix_in_8[38]), .Y(top_core_EC_mc_n336) );
  XOR2X1 U10524 ( .A(top_core_EC_mc_mix_in_4_16_), .B(
        top_core_EC_mc_mix_in_2_16_), .Y(top_core_EC_mc_mix_in_8[18]) );
  XOR2X1 U10525 ( .A(top_core_EC_mc_mix_in_4_16_), .B(
        top_core_EC_mc_mix_in_2_19_), .Y(top_core_EC_mc_mix_in_8[21]) );
  XOR2X1 U10526 ( .A(top_core_EC_mc_mix_in_2_16_), .B(
        top_core_EC_mc_mix_in_2_0_), .Y(top_core_EC_mc_n571) );
  XOR2X1 U10527 ( .A(top_core_EC_mc_mix_in_2_58_), .B(
        top_core_EC_mc_mix_in_4_50_), .Y(top_core_EC_mc_n443) );
  AOI22X1 U10528 ( .A0(n722), .A1(n5392), .B0(n353), .B1(n993), .Y(n10048) );
  AOI22X1 U10529 ( .A0(n723), .A1(n6176), .B0(n354), .B1(n1135), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n234) );
  AOI22X1 U10530 ( .A0(n724), .A1(n5038), .B0(n356), .B1(n937), .Y(n11216) );
  AOI22X1 U10531 ( .A0(n725), .A1(n5864), .B0(n355), .B1(n1077), .Y(n8296) );
  AOI22X1 U10532 ( .A0(n731), .A1(n5122), .B0(n357), .B1(n951), .Y(n10924) );
  AOI22X1 U10533 ( .A0(n733), .A1(n5628), .B0(n359), .B1(n1035), .Y(n9172) );
  AOI22X1 U10534 ( .A0(n735), .A1(n6092), .B0(n358), .B1(n1119), .Y(n7420) );
  AOI22X1 U10535 ( .A0(n737), .A1(n5308), .B0(n360), .B1(n979), .Y(n10340) );
  AOI22X1 U10536 ( .A0(n730), .A1(n5552), .B0(n361), .B1(n1021), .Y(n9464) );
  AOI22X1 U10537 ( .A0(n726), .A1(n5780), .B0(n362), .B1(n1063), .Y(n8588) );
  AOI22X1 U10538 ( .A0(n732), .A1(n6016), .B0(n363), .B1(n1105), .Y(n7712) );
  AOI22X1 U10539 ( .A0(n728), .A1(n4922), .B0(n364), .B1(n923), .Y(n11508) );
  AOI22X1 U10540 ( .A0(n734), .A1(n5230), .B0(n365), .B1(n965), .Y(n10632) );
  AOI22X1 U10541 ( .A0(n727), .A1(n5476), .B0(n366), .B1(n1007), .Y(n9756) );
  AOI22X1 U10542 ( .A0(n736), .A1(n5704), .B0(n367), .B1(n1049), .Y(n8880) );
  AOI22X1 U10543 ( .A0(n729), .A1(n5940), .B0(n368), .B1(n1091), .Y(n8004) );
  XOR2X1 U10544 ( .A(top_core_EC_mc_mix_in_2_10_), .B(
        top_core_EC_mc_mix_in_4_2_), .Y(top_core_EC_mc_n621) );
  XOR2X1 U10545 ( .A(top_core_EC_mc_mix_in_2_42_), .B(
        top_core_EC_mc_mix_in_4_34_), .Y(top_core_EC_mc_n369) );
  AOI22X1 U10546 ( .A0(n417), .A1(n5376), .B0(n698), .B1(n2880), .Y(n9968) );
  AOI22X1 U10547 ( .A0(n418), .A1(n6166), .B0(n699), .B1(n3481), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n154) );
  AOI22X1 U10548 ( .A0(n419), .A1(n5022), .B0(n700), .B1(n2638), .Y(n11136) );
  AOI22X1 U10549 ( .A0(n420), .A1(n5848), .B0(n701), .B1(n3240), .Y(n8216) );
  AOI22X1 U10550 ( .A0(n421), .A1(n5106), .B0(n707), .B1(n2699), .Y(n10844) );
  AOI22X1 U10551 ( .A0(n422), .A1(n5612), .B0(n709), .B1(n3060), .Y(n9092) );
  AOI22X1 U10552 ( .A0(n423), .A1(n6076), .B0(n711), .B1(n3420), .Y(n7340) );
  AOI22X1 U10553 ( .A0(n424), .A1(n5292), .B0(n713), .B1(n2820), .Y(n10260) );
  AOI22X1 U10554 ( .A0(n425), .A1(n5536), .B0(n706), .B1(n3002), .Y(n9384) );
  AOI22X1 U10555 ( .A0(n426), .A1(n5764), .B0(n702), .B1(n3179), .Y(n8508) );
  AOI22X1 U10556 ( .A0(n427), .A1(n6000), .B0(n708), .B1(n3362), .Y(n7632) );
  AOI22X1 U10557 ( .A0(n428), .A1(n4906), .B0(n704), .B1(n2577), .Y(n11428) );
  AOI22X1 U10558 ( .A0(n429), .A1(n5214), .B0(n710), .B1(n2759), .Y(n10552) );
  AOI22X1 U10559 ( .A0(n430), .A1(n5460), .B0(n703), .B1(n2941), .Y(n9676) );
  AOI22X1 U10560 ( .A0(n431), .A1(n5688), .B0(n712), .B1(n3121), .Y(n8800) );
  AOI22X1 U10561 ( .A0(n432), .A1(n5924), .B0(n705), .B1(n3301), .Y(n7924) );
  XOR2X1 U10562 ( .A(n1543), .B(top_core_EC_mc_mix_in_8[32]), .Y(
        top_core_EC_mc_n320) );
  XOR2X1 U10563 ( .A(n1542), .B(top_core_EC_mc_mix_in_4_32_), .Y(
        top_core_EC_mc_n312) );
  NAND2X1 U10564 ( .A(n6915), .B(n6826), .Y(n11677) );
  NAND2X1 U10565 ( .A(n6869), .B(n6804), .Y(top_core_KE_sb1_n102) );
  NAND2X1 U10566 ( .A(n6622), .B(n6530), .Y(n12308) );
  NAND2X1 U10567 ( .A(n6550), .B(n6472), .Y(n13254) );
  NAND2X1 U10568 ( .A(n6575), .B(n6507), .Y(n11993) );
  NAND2X1 U10569 ( .A(n6845), .B(n6775), .Y(n12624) );
  NAND2X1 U10570 ( .A(n6598), .B(n6519), .Y(n13569) );
  NAND2X1 U10571 ( .A(n6891), .B(n6815), .Y(n12939) );
  XOR2X1 U10572 ( .A(n1545), .B(top_core_EC_mc_mix_in_4_16_), .Y(
        top_core_EC_mc_n633) );
  XOR2X1 U10573 ( .A(n1546), .B(top_core_EC_mc_mix_in_8[16]), .Y(
        top_core_EC_mc_n639) );
  XOR2X1 U10574 ( .A(top_core_EC_mc_mix_in_8[7]), .B(
        top_core_EC_mc_mix_in_8[23]), .Y(top_core_EC_mc_n254) );
  XOR2X1 U10575 ( .A(top_core_EC_mc_mix_in_8[55]), .B(
        top_core_EC_mc_mix_in_8[39]), .Y(top_core_EC_mc_n391) );
  XOR2X1 U10576 ( .A(top_core_EC_mc_mix_in_8[23]), .B(
        top_core_EC_mc_mix_in_8[7]), .Y(top_core_EC_mc_n601) );
  XOR2X1 U10577 ( .A(top_core_EC_mix_in[8]), .B(top_core_EC_mc_mix_in_2_0_), 
        .Y(top_core_EC_mc_n627) );
  XOR2X1 U10578 ( .A(top_core_EC_mix_in[56]), .B(top_core_EC_mc_mix_in_2_48_), 
        .Y(top_core_EC_mc_n451) );
  XOR2X1 U10579 ( .A(top_core_EC_mix_in[40]), .B(top_core_EC_mc_mix_in_2_32_), 
        .Y(top_core_EC_mc_n377) );
  XOR2X1 U10580 ( .A(n1546), .B(top_core_EC_mc_mix_in_2_26_), .Y(
        top_core_EC_mc_mix_in_4_27_) );
  XOR2X1 U10581 ( .A(top_core_EC_mc_mix_in_2_18_), .B(
        top_core_EC_mc_mix_in_2_2_), .Y(top_core_EC_mc_n9) );
  XOR2X1 U10582 ( .A(top_core_EC_mix_in[26]), .B(top_core_EC_mc_mix_in_2_18_), 
        .Y(top_core_EC_mc_n670) );
  XOR2X1 U10583 ( .A(top_core_EC_mix_in[27]), .B(top_core_EC_mc_mix_in_2_19_), 
        .Y(top_core_EC_mc_n664) );
  XOR2X1 U10584 ( .A(top_core_EC_mix_in[42]), .B(top_core_EC_mc_mix_in_2_34_), 
        .Y(top_core_EC_mc_n361) );
  XOR2X1 U10585 ( .A(top_core_EC_mix_in[43]), .B(top_core_EC_mc_mix_in_2_35_), 
        .Y(top_core_EC_mc_n353) );
  XOR2X1 U10586 ( .A(top_core_EC_mix_in[0]), .B(top_core_EC_mix_in[16]), .Y(
        top_core_EC_mc_n102) );
  XOR2X1 U10587 ( .A(top_core_EC_mix_in[18]), .B(top_core_EC_mix_in[2]), .Y(
        top_core_EC_mc_n615) );
  XOR2X1 U10588 ( .A(top_core_EC_mix_in[19]), .B(top_core_EC_mix_in[3]), .Y(
        top_core_EC_mc_n608) );
  XOR2X1 U10589 ( .A(top_core_EC_mc_mix_in_4_58_), .B(
        top_core_EC_mc_mix_in_4_42_), .Y(top_core_EC_mc_n360) );
  XOR2X1 U10590 ( .A(top_core_EC_mc_mix_in_4_90_), .B(
        top_core_EC_mc_mix_in_4_74_), .Y(top_core_EC_mc_n92) );
  XOR2X1 U10591 ( .A(top_core_EC_mc_mix_in_4_122_), .B(
        top_core_EC_mc_mix_in_4_106_), .Y(top_core_EC_mc_n756) );
  XOR2X1 U10592 ( .A(top_core_EC_mc_mix_in_8[62]), .B(
        top_core_EC_mc_mix_in_8[46]), .Y(top_core_EC_mc_n327) );
  XOR2X1 U10593 ( .A(top_core_EC_mc_mix_in_8[94]), .B(
        top_core_EC_mc_mix_in_8[78]), .Y(top_core_EC_mc_n68) );
  XOR2X1 U10594 ( .A(top_core_EC_mc_mix_in_8[126]), .B(
        top_core_EC_mc_mix_in_8[110]), .Y(top_core_EC_mc_n733) );
  XOR2X1 U10595 ( .A(n1544), .B(top_core_EC_mc_mix_in_8[39]), .Y(
        top_core_EC_mc_n328) );
  XOR2X1 U10596 ( .A(n1547), .B(top_core_EC_mc_mix_in_8[23]), .Y(
        top_core_EC_mc_n645) );
  XOR2X1 U10597 ( .A(top_core_EC_mc_mix_in_4_82_), .B(
        top_core_EC_mc_mix_in_4_66_), .Y(top_core_EC_mc_n164) );
  XOR2X1 U10598 ( .A(top_core_EC_mc_mix_in_8[86]), .B(
        top_core_EC_mc_mix_in_8[70]), .Y(top_core_EC_mc_n140) );
  XOR2X1 U10599 ( .A(top_core_EC_mc_mix_in_4_98_), .B(
        top_core_EC_mc_mix_in_4_114_), .Y(top_core_EC_mc_n25) );
  XOR2X1 U10600 ( .A(top_core_EC_mc_mix_in_8[118]), .B(
        top_core_EC_mc_mix_in_8[102]), .Y(top_core_EC_mc_n799) );
  XOR2X1 U10601 ( .A(top_core_EC_mc_mix_in_8[82]), .B(
        top_core_EC_mc_mix_in_8[66]), .Y(top_core_EC_mc_n172) );
  XOR2X1 U10602 ( .A(top_core_EC_mc_mix_in_4_83_), .B(
        top_core_EC_mc_mix_in_4_67_), .Y(top_core_EC_mc_n156) );
  XOR2X1 U10603 ( .A(top_core_EC_mc_mix_in_8[85]), .B(
        top_core_EC_mc_mix_in_8[69]), .Y(top_core_EC_mc_n148) );
  XOR2X1 U10604 ( .A(top_core_EC_mc_mix_in_4_99_), .B(
        top_core_EC_mc_mix_in_4_115_), .Y(top_core_EC_mc_n16) );
  XOR2X1 U10605 ( .A(top_core_EC_mc_mix_in_8[117]), .B(
        top_core_EC_mc_mix_in_8[101]), .Y(top_core_EC_mc_n807) );
  XOR2X1 U10606 ( .A(top_core_EC_mc_mix_in_4_59_), .B(
        top_core_EC_mc_mix_in_4_43_), .Y(top_core_EC_mc_n352) );
  XOR2X1 U10607 ( .A(top_core_EC_mc_mix_in_4_91_), .B(
        top_core_EC_mc_mix_in_4_75_), .Y(top_core_EC_mc_n84) );
  XOR2X1 U10608 ( .A(top_core_EC_mc_mix_in_4_123_), .B(
        top_core_EC_mc_mix_in_4_107_), .Y(top_core_EC_mc_n749) );
  XOR2X1 U10609 ( .A(top_core_EC_mc_mix_in_8[122]), .B(
        top_core_EC_mc_mix_in_8[106]), .Y(top_core_EC_mc_n763) );
  XOR2X1 U10610 ( .A(top_core_EC_mc_n77), .B(top_core_EC_mc_n78), .Y(
        top_core_EC_mc_n75) );
  XOR2X1 U10611 ( .A(top_core_EC_mc_n742), .B(top_core_EC_mc_n743), .Y(
        top_core_EC_mc_n740) );
  XOR2X1 U10612 ( .A(top_core_EC_mc_n110), .B(top_core_EC_mc_n111), .Y(
        top_core_EC_mc_n108) );
  XOR2X1 U10613 ( .A(top_core_EC_mc_n61), .B(top_core_EC_mc_n62), .Y(
        top_core_EC_mc_n59) );
  XOR2X1 U10614 ( .A(top_core_EC_mc_n53), .B(top_core_EC_mc_n54), .Y(
        top_core_EC_mc_n51) );
  XOR2X1 U10615 ( .A(top_core_EC_mc_n726), .B(top_core_EC_mc_n727), .Y(
        top_core_EC_mc_n724) );
  XOR2X1 U10616 ( .A(top_core_EC_mc_n718), .B(top_core_EC_mc_n719), .Y(
        top_core_EC_mc_n716) );
  XOR2X1 U10617 ( .A(top_core_EC_mc_n118), .B(top_core_EC_mc_n119), .Y(
        top_core_EC_mc_n116) );
  XOR2X1 U10618 ( .A(top_core_EC_mc_n93), .B(top_core_EC_mc_n94), .Y(
        top_core_EC_mc_n91) );
  XOR2X1 U10619 ( .A(top_core_EC_mc_n85), .B(top_core_EC_mc_n86), .Y(
        top_core_EC_mc_n83) );
  XOR2X1 U10620 ( .A(top_core_EC_mc_n69), .B(top_core_EC_mc_n70), .Y(
        top_core_EC_mc_n67) );
  XOR2X1 U10621 ( .A(top_core_EC_mc_n771), .B(top_core_EC_mc_n46), .Y(
        top_core_EC_mc_n769) );
  XOR2X1 U10622 ( .A(top_core_EC_mc_n764), .B(top_core_EC_mc_n37), .Y(
        top_core_EC_mc_n762) );
  XOR2X1 U10623 ( .A(top_core_EC_mc_n757), .B(top_core_EC_mc_n28), .Y(
        top_core_EC_mc_n755) );
  XOR2X1 U10624 ( .A(top_core_EC_mc_n750), .B(top_core_EC_mc_n19), .Y(
        top_core_EC_mc_n748) );
  XOR2X1 U10625 ( .A(top_core_EC_mc_n734), .B(top_core_EC_mc_n735), .Y(
        top_core_EC_mc_n732) );
  XOR2X1 U10626 ( .A(top_core_EC_mc_mix_in_8[98]), .B(
        top_core_EC_mc_mix_in_8[114]), .Y(top_core_EC_mc_n34) );
  XOR2X1 U10627 ( .A(top_core_EC_mc_mix_in_8[58]), .B(
        top_core_EC_mc_mix_in_8[42]), .Y(top_core_EC_mc_n368) );
  XOR2X1 U10628 ( .A(top_core_EC_mc_mix_in_8[61]), .B(
        top_core_EC_mc_mix_in_8[45]), .Y(top_core_EC_mc_n335) );
  XOR2X1 U10629 ( .A(top_core_EC_mc_mix_in_8[90]), .B(
        top_core_EC_mc_mix_in_8[74]), .Y(top_core_EC_mc_n109) );
  XOR2X1 U10630 ( .A(top_core_EC_mc_mix_in_8[93]), .B(
        top_core_EC_mc_mix_in_8[77]), .Y(top_core_EC_mc_n76) );
  XOR2X1 U10631 ( .A(top_core_EC_mc_mix_in_8[125]), .B(
        top_core_EC_mc_mix_in_8[109]), .Y(top_core_EC_mc_n741) );
  XNOR2X1 U10632 ( .A(top_core_EC_mc_n658), .B(top_core_EC_mc_n621), .Y(
        top_core_EC_mc_n656) );
  XNOR2X1 U10633 ( .A(top_core_EC_mc_mix_in_2_18_), .B(
        top_core_EC_mc_mix_in_4_10_), .Y(top_core_EC_mc_n658) );
  XNOR2X1 U10634 ( .A(top_core_EC_mc_n586), .B(top_core_EC_mc_n587), .Y(
        top_core_EC_mc_n583) );
  XNOR2X1 U10635 ( .A(top_core_EC_mix_in[18]), .B(top_core_EC_mc_mix_in_2_10_), 
        .Y(top_core_EC_mc_n586) );
  XNOR2X1 U10636 ( .A(top_core_EC_mc_n499), .B(top_core_EC_mc_n500), .Y(
        top_core_EC_mc_n496) );
  XNOR2X1 U10637 ( .A(top_core_EC_mix_in[19]), .B(top_core_EC_mc_mix_in_2_11_), 
        .Y(top_core_EC_mc_n499) );
  XNOR2X1 U10638 ( .A(top_core_EC_mc_n434), .B(top_core_EC_mc_n435), .Y(
        top_core_EC_mc_n431) );
  XNOR2X1 U10639 ( .A(top_core_EC_mc_mix_in_8[23]), .B(
        top_core_EC_mc_mix_in_8[14]), .Y(top_core_EC_mc_n434) );
  XNOR2X1 U10640 ( .A(top_core_EC_mc_n345), .B(top_core_EC_mc_n346), .Y(
        top_core_EC_mc_n342) );
  XNOR2X1 U10641 ( .A(top_core_EC_mc_mix_in_8[16]), .B(
        top_core_EC_mc_mix_in_8[15]), .Y(top_core_EC_mc_n345) );
  XNOR2X1 U10642 ( .A(top_core_EC_mc_n256), .B(top_core_EC_mc_n257), .Y(
        top_core_EC_mc_n253) );
  XNOR2X1 U10643 ( .A(top_core_EC_mc_mix_in_4_16_), .B(n1550), .Y(
        top_core_EC_mc_n256) );
  XNOR2X1 U10644 ( .A(top_core_EC_mc_n191), .B(top_core_EC_mc_n192), .Y(
        top_core_EC_mc_n188) );
  XNOR2X1 U10645 ( .A(top_core_EC_mc_mix_in_2_16_), .B(n1549), .Y(
        top_core_EC_mc_n191) );
  XNOR2X1 U10646 ( .A(top_core_EC_mc_n683), .B(top_core_EC_mc_n103), .Y(
        top_core_EC_mc_n681) );
  XNOR2X1 U10647 ( .A(top_core_EC_mix_in[0]), .B(top_core_EC_mix_in[8]), .Y(
        top_core_EC_mc_n683) );
  XNOR2X1 U10648 ( .A(top_core_EC_mc_n450), .B(top_core_EC_mc_n451), .Y(
        top_core_EC_mc_n447) );
  XNOR2X1 U10649 ( .A(top_core_EC_mix_in[32]), .B(top_core_EC_mix_in[40]), .Y(
        top_core_EC_mc_n450) );
  XNOR2X1 U10650 ( .A(top_core_EC_mc_n442), .B(top_core_EC_mc_n443), .Y(
        top_core_EC_mc_n439) );
  XNOR2X1 U10651 ( .A(top_core_EC_mc_mix_in_2_34_), .B(
        top_core_EC_mc_mix_in_2_42_), .Y(top_core_EC_mc_n442) );
  XNOR2X1 U10652 ( .A(top_core_EC_mc_n425), .B(top_core_EC_mc_n426), .Y(
        top_core_EC_mc_n422) );
  XNOR2X1 U10653 ( .A(top_core_EC_mix_in[34]), .B(top_core_EC_mix_in[42]), .Y(
        top_core_EC_mc_n425) );
  XNOR2X1 U10654 ( .A(top_core_EC_mc_n417), .B(top_core_EC_mc_n418), .Y(
        top_core_EC_mc_n414) );
  XNOR2X1 U10655 ( .A(top_core_EC_mix_in[35]), .B(top_core_EC_mix_in[43]), .Y(
        top_core_EC_mc_n417) );
  XNOR2X1 U10656 ( .A(top_core_EC_mc_n409), .B(top_core_EC_mc_n410), .Y(
        top_core_EC_mc_n406) );
  XNOR2X1 U10657 ( .A(top_core_EC_mc_mix_in_8[39]), .B(
        top_core_EC_mc_mix_in_8[47]), .Y(top_core_EC_mc_n409) );
  XNOR2X1 U10658 ( .A(top_core_EC_mc_n401), .B(top_core_EC_mc_n402), .Y(
        top_core_EC_mc_n398) );
  XNOR2X1 U10659 ( .A(top_core_EC_mc_mix_in_8[32]), .B(n1544), .Y(
        top_core_EC_mc_n401) );
  XNOR2X1 U10660 ( .A(top_core_EC_mc_n393), .B(top_core_EC_mc_n394), .Y(
        top_core_EC_mc_n390) );
  XNOR2X1 U10661 ( .A(top_core_EC_mc_mix_in_4_32_), .B(n1543), .Y(
        top_core_EC_mc_n393) );
  XNOR2X1 U10662 ( .A(top_core_EC_mc_n385), .B(top_core_EC_mc_n386), .Y(
        top_core_EC_mc_n382) );
  XNOR2X1 U10663 ( .A(top_core_EC_mc_mix_in_2_32_), .B(n1542), .Y(
        top_core_EC_mc_n385) );
  XOR2X1 U10664 ( .A(n1546), .B(top_core_EC_mc_mix_in_2_27_), .Y(
        top_core_EC_mc_mix_in_8[29]) );
  XOR2X1 U10665 ( .A(n1547), .B(n1550), .Y(top_core_EC_mc_n570) );
  XOR2X1 U10666 ( .A(n1549), .B(n1546), .Y(top_core_EC_mc_n100) );
  XOR2X1 U10667 ( .A(n1549), .B(n1548), .Y(top_core_EC_mc_mix_in_8[10]) );
  XOR2X1 U10668 ( .A(n1543), .B(n1542), .Y(top_core_EC_mc_mix_in_8[42]) );
  XOR2X1 U10669 ( .A(n1543), .B(top_core_EC_mc_mix_in_2_43_), .Y(
        top_core_EC_mc_mix_in_8[45]) );
  NAND2X1 U10670 ( .A(n995), .B(n5335), .Y(n17239) );
  NAND2X1 U10671 ( .A(n1134), .B(n6118), .Y(n14089) );
  NAND2X1 U10672 ( .A(n1079), .B(n5807), .Y(n15349) );
  NAND2X1 U10673 ( .A(n939), .B(n4981), .Y(n18499) );
  NAND2X1 U10674 ( .A(n1065), .B(n5723), .Y(n15664) );
  NAND2X1 U10675 ( .A(n1009), .B(n5419), .Y(n16924) );
  NAND2X1 U10676 ( .A(n925), .B(n4865), .Y(n18814) );
  NAND2X1 U10677 ( .A(n1093), .B(n5883), .Y(n15034) );
  NAND2X1 U10678 ( .A(n1023), .B(n5495), .Y(n16609) );
  NAND2X1 U10679 ( .A(n953), .B(n5065), .Y(n18184) );
  NAND2X1 U10680 ( .A(n1107), .B(n5959), .Y(n14719) );
  NAND2X1 U10681 ( .A(n1037), .B(n5571), .Y(n16294) );
  NAND2X1 U10682 ( .A(n967), .B(n5173), .Y(n17869) );
  NAND2X1 U10683 ( .A(n1121), .B(n6035), .Y(n14404) );
  NAND2X1 U10684 ( .A(n1051), .B(n5647), .Y(n15979) );
  NAND2X1 U10685 ( .A(n981), .B(n5251), .Y(n17554) );
  INVX1 U10686 ( .A(n13770), .Y(n6606) );
  XOR2X1 U10687 ( .A(top_core_EC_mc_mix_in_4_0_), .B(
        top_core_EC_mc_mix_in_2_0_), .Y(top_core_EC_mc_mix_in_8[2]) );
  XOR2X1 U10688 ( .A(top_core_EC_mc_mix_in_4_0_), .B(
        top_core_EC_mc_mix_in_2_3_), .Y(top_core_EC_mc_mix_in_8[5]) );
  NAND2X1 U10689 ( .A(n3481), .B(n13918), .Y(n13882) );
  NAND2X1 U10690 ( .A(n2880), .B(n17068), .Y(n17032) );
  NAND2X1 U10691 ( .A(n2638), .B(n18328), .Y(n18292) );
  NAND2X1 U10692 ( .A(n3240), .B(n15178), .Y(n15142) );
  NAND2X1 U10693 ( .A(n3179), .B(n15493), .Y(n15457) );
  NAND2X1 U10694 ( .A(n2941), .B(n16753), .Y(n16717) );
  NAND2X1 U10695 ( .A(n2577), .B(n18643), .Y(n18607) );
  NAND2X1 U10696 ( .A(n3301), .B(n14863), .Y(n14827) );
  NAND2X1 U10697 ( .A(n3002), .B(n16438), .Y(n16402) );
  NAND2X1 U10698 ( .A(n2699), .B(n18013), .Y(n17977) );
  NAND2X1 U10699 ( .A(n3362), .B(n14548), .Y(n14512) );
  NAND2X1 U10700 ( .A(n3060), .B(n16123), .Y(n16087) );
  NAND2X1 U10701 ( .A(n2759), .B(n17698), .Y(n17662) );
  NAND2X1 U10702 ( .A(n3420), .B(n14233), .Y(n14197) );
  NAND2X1 U10703 ( .A(n3121), .B(n15808), .Y(n15772) );
  NAND2X1 U10704 ( .A(n2820), .B(n17383), .Y(n17347) );
  NAND2X1 U10705 ( .A(n6597), .B(n1178), .Y(n13617) );
  CLKINVX3 U10706 ( .A(n11658), .Y(n6909) );
  CLKINVX3 U10707 ( .A(top_core_KE_sb1_n83), .Y(n6863) );
  CLKINVX3 U10708 ( .A(n13235), .Y(n6544) );
  CLKINVX3 U10709 ( .A(n11974), .Y(n6569) );
  CLKINVX3 U10710 ( .A(n12920), .Y(n6885) );
  CLKINVX3 U10711 ( .A(n13550), .Y(n6592) );
  CLKINVX3 U10712 ( .A(n12605), .Y(n6839) );
  AOI22X1 U10713 ( .A0(n17195), .A1(n529), .B0(n17010), .B1(n995), .Y(n17190)
         );
  AOI22X1 U10714 ( .A0(n14045), .A1(n530), .B0(n13860), .B1(n1134), .Y(n14040)
         );
  AOI22X1 U10715 ( .A0(n18455), .A1(n531), .B0(n18270), .B1(n939), .Y(n18450)
         );
  AOI22X1 U10716 ( .A0(n15305), .A1(n532), .B0(n15120), .B1(n1079), .Y(n15300)
         );
  AOI22X1 U10717 ( .A0(n15620), .A1(n538), .B0(n15435), .B1(n1065), .Y(n15615)
         );
  AOI22X1 U10718 ( .A0(n16880), .A1(n542), .B0(n16695), .B1(n1009), .Y(n16875)
         );
  AOI22X1 U10719 ( .A0(n18770), .A1(n540), .B0(n18585), .B1(n925), .Y(n18765)
         );
  AOI22X1 U10720 ( .A0(n14990), .A1(n544), .B0(n14805), .B1(n1093), .Y(n14985)
         );
  AOI22X1 U10721 ( .A0(n16565), .A1(n537), .B0(n16380), .B1(n1023), .Y(n16560)
         );
  AOI22X1 U10722 ( .A0(n18140), .A1(n533), .B0(n17955), .B1(n953), .Y(n18135)
         );
  AOI22X1 U10723 ( .A0(n14675), .A1(n539), .B0(n14490), .B1(n1107), .Y(n14670)
         );
  AOI22X1 U10724 ( .A0(n16250), .A1(n534), .B0(n16065), .B1(n1037), .Y(n16245)
         );
  AOI22X1 U10725 ( .A0(n17825), .A1(n541), .B0(n17640), .B1(n967), .Y(n17820)
         );
  AOI22X1 U10726 ( .A0(n14360), .A1(n535), .B0(n14175), .B1(n1121), .Y(n14355)
         );
  AOI22X1 U10727 ( .A0(n15935), .A1(n543), .B0(n15750), .B1(n1051), .Y(n15930)
         );
  AOI22X1 U10728 ( .A0(n17510), .A1(n536), .B0(n17325), .B1(n981), .Y(n17505)
         );
  AOI22XL U10729 ( .A0(n17065), .A1(n106), .B0(n5357), .B1(n401), .Y(n17063)
         );
  AOI22XL U10730 ( .A0(n13915), .A1(n107), .B0(n6125), .B1(n402), .Y(n13913)
         );
  AOI22XL U10731 ( .A0(n18325), .A1(n108), .B0(n5003), .B1(n403), .Y(n18323)
         );
  AOI22XL U10732 ( .A0(n15175), .A1(n109), .B0(n5829), .B1(n404), .Y(n15173)
         );
  AOI22XL U10733 ( .A0(n15490), .A1(n110), .B0(n5745), .B1(n410), .Y(n15488)
         );
  AOI22XL U10734 ( .A0(n18640), .A1(n111), .B0(n4887), .B1(n412), .Y(n18638)
         );
  AOI22XL U10735 ( .A0(n16750), .A1(n112), .B0(n5441), .B1(n414), .Y(n16748)
         );
  AOI22XL U10736 ( .A0(n14860), .A1(n113), .B0(n5905), .B1(n416), .Y(n14858)
         );
  AOI22XL U10737 ( .A0(n16435), .A1(n114), .B0(n5517), .B1(n409), .Y(n16433)
         );
  AOI22XL U10738 ( .A0(n18010), .A1(n115), .B0(n5087), .B1(n405), .Y(n18008)
         );
  AOI22XL U10739 ( .A0(n14545), .A1(n116), .B0(n5981), .B1(n411), .Y(n14543)
         );
  AOI22XL U10740 ( .A0(n16120), .A1(n117), .B0(n5593), .B1(n406), .Y(n16118)
         );
  AOI22XL U10741 ( .A0(n17695), .A1(n118), .B0(n5195), .B1(n413), .Y(n17693)
         );
  AOI22XL U10742 ( .A0(n14230), .A1(n119), .B0(n6057), .B1(n407), .Y(n14228)
         );
  AOI22XL U10743 ( .A0(n15805), .A1(n120), .B0(n5669), .B1(n415), .Y(n15803)
         );
  AOI22XL U10744 ( .A0(n17380), .A1(n121), .B0(n5273), .B1(n408), .Y(n17378)
         );
  XNOR2X1 U10745 ( .A(top_core_EC_mc_mix_in_8[31]), .B(top_core_EC_mc_n344), 
        .Y(top_core_EC_mc_n590) );
  AOI22X1 U10746 ( .A0(n2846), .A1(n17273), .B0(n17274), .B1(n2848), .Y(n17272) );
  OAI211X1 U10747 ( .A0(n1003), .A1(n17275), .B0(n17276), .C0(n17277), .Y(
        n17274) );
  OAI211X1 U10748 ( .A0(n2897), .A1(n17275), .B0(n17281), .C0(n17282), .Y(
        n17273) );
  AOI22X1 U10749 ( .A0(n3447), .A1(n14123), .B0(n14124), .B1(n3450), .Y(n14122) );
  OAI211X1 U10750 ( .A0(n1142), .A1(n14125), .B0(n14126), .C0(n14127), .Y(
        n14124) );
  OAI211X1 U10751 ( .A0(n3498), .A1(n14125), .B0(n14131), .C0(n14132), .Y(
        n14123) );
  AOI22X1 U10752 ( .A0(n3206), .A1(n15383), .B0(n15384), .B1(n3208), .Y(n15382) );
  OAI211X1 U10753 ( .A0(n1087), .A1(n15385), .B0(n15386), .C0(n15387), .Y(
        n15384) );
  OAI211X1 U10754 ( .A0(n3257), .A1(n15385), .B0(n15391), .C0(n15392), .Y(
        n15383) );
  AOI22X1 U10755 ( .A0(n2604), .A1(n18533), .B0(n18534), .B1(n2606), .Y(n18532) );
  OAI211X1 U10756 ( .A0(n947), .A1(n18535), .B0(n18536), .C0(n18537), .Y(
        n18534) );
  OAI211X1 U10757 ( .A0(n2654), .A1(n18535), .B0(n18541), .C0(n18542), .Y(
        n18533) );
  AOI22X1 U10758 ( .A0(n3145), .A1(n15698), .B0(n15699), .B1(n3147), .Y(n15697) );
  OAI211X1 U10759 ( .A0(n1073), .A1(n15700), .B0(n15701), .C0(n15702), .Y(
        n15699) );
  OAI211X1 U10760 ( .A0(n3196), .A1(n15700), .B0(n15706), .C0(n15707), .Y(
        n15698) );
  AOI22X1 U10761 ( .A0(n2907), .A1(n16958), .B0(n16959), .B1(n2909), .Y(n16957) );
  OAI211X1 U10762 ( .A0(n1017), .A1(n16960), .B0(n16961), .C0(n16962), .Y(
        n16959) );
  OAI211X1 U10763 ( .A0(n2958), .A1(n16960), .B0(n16966), .C0(n16967), .Y(
        n16958) );
  AOI22X1 U10764 ( .A0(n2543), .A1(n18848), .B0(n18849), .B1(n2545), .Y(n18847) );
  OAI211X1 U10765 ( .A0(n933), .A1(n18850), .B0(n18851), .C0(n18852), .Y(
        n18849) );
  OAI211X1 U10766 ( .A0(n2593), .A1(n18850), .B0(n18856), .C0(n18857), .Y(
        n18848) );
  AOI22X1 U10767 ( .A0(n3267), .A1(n15068), .B0(n15069), .B1(n3269), .Y(n15067) );
  OAI211X1 U10768 ( .A0(n1101), .A1(n15070), .B0(n15071), .C0(n15072), .Y(
        n15069) );
  OAI211X1 U10769 ( .A0(n3320), .A1(n15070), .B0(n15076), .C0(n15077), .Y(
        n15068) );
  AOI22X1 U10770 ( .A0(n2968), .A1(n16643), .B0(n16644), .B1(n2970), .Y(n16642) );
  OAI211X1 U10771 ( .A0(n1031), .A1(n16645), .B0(n16646), .C0(n16647), .Y(
        n16644) );
  OAI211X1 U10772 ( .A0(n3021), .A1(n16645), .B0(n16651), .C0(n16652), .Y(
        n16643) );
  AOI22X1 U10773 ( .A0(n2665), .A1(n18218), .B0(n18219), .B1(n2667), .Y(n18217) );
  OAI211X1 U10774 ( .A0(n961), .A1(n18220), .B0(n18221), .C0(n18222), .Y(
        n18219) );
  OAI211X1 U10775 ( .A0(n2715), .A1(n18220), .B0(n18226), .C0(n18227), .Y(
        n18218) );
  AOI22X1 U10776 ( .A0(n3328), .A1(n14753), .B0(n14754), .B1(n3330), .Y(n14752) );
  OAI211X1 U10777 ( .A0(n1115), .A1(n14755), .B0(n14756), .C0(n14757), .Y(
        n14754) );
  OAI211X1 U10778 ( .A0(n3381), .A1(n14755), .B0(n14761), .C0(n14762), .Y(
        n14753) );
  AOI22X1 U10779 ( .A0(n3026), .A1(n16328), .B0(n16329), .B1(n3028), .Y(n16327) );
  OAI211X1 U10780 ( .A0(n1045), .A1(n16330), .B0(n16331), .C0(n16332), .Y(
        n16329) );
  OAI211X1 U10781 ( .A0(n3076), .A1(n16330), .B0(n16336), .C0(n16337), .Y(
        n16328) );
  AOI22X1 U10782 ( .A0(n2725), .A1(n17903), .B0(n17904), .B1(n2727), .Y(n17902) );
  OAI211X1 U10783 ( .A0(n975), .A1(n17905), .B0(n17906), .C0(n17907), .Y(
        n17904) );
  OAI211X1 U10784 ( .A0(n2780), .A1(n17905), .B0(n17911), .C0(n17912), .Y(
        n17903) );
  AOI22X1 U10785 ( .A0(n3386), .A1(n14438), .B0(n14439), .B1(n3388), .Y(n14437) );
  OAI211X1 U10786 ( .A0(n1129), .A1(n14440), .B0(n14441), .C0(n14442), .Y(
        n14439) );
  OAI211X1 U10787 ( .A0(n3437), .A1(n14440), .B0(n14446), .C0(n14447), .Y(
        n14438) );
  AOI22X1 U10788 ( .A0(n3087), .A1(n16013), .B0(n16014), .B1(n3089), .Y(n16012) );
  OAI211X1 U10789 ( .A0(n1059), .A1(n16015), .B0(n16016), .C0(n16017), .Y(
        n16014) );
  OAI211X1 U10790 ( .A0(n3140), .A1(n16015), .B0(n16021), .C0(n16022), .Y(
        n16013) );
  AOI22X1 U10791 ( .A0(n2786), .A1(n17588), .B0(n17589), .B1(n2788), .Y(n17587) );
  OAI211X1 U10792 ( .A0(n989), .A1(n17590), .B0(n17591), .C0(n17592), .Y(
        n17589) );
  OAI211X1 U10793 ( .A0(n2840), .A1(n17590), .B0(n17596), .C0(n17597), .Y(
        n17588) );
  XNOR2X1 U10794 ( .A(top_core_EC_mc_mix_in_2_26_), .B(top_core_EC_mc_n585), 
        .Y(top_core_EC_mc_n611) );
  XNOR2X1 U10795 ( .A(top_core_EC_mc_mix_in_2_58_), .B(top_core_EC_mc_n424), 
        .Y(top_core_EC_mc_n357) );
  NAND4BBX1 U10796 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n111), .BN(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n112), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n113), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n101), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n110) );
  NAND4BBX1 U10797 ( .AN(n9926), .BN(n9927), .C(n9928), .D(n9917), .Y(n9925)
         );
  NAND4BBX1 U10798 ( .AN(n11094), .BN(n11095), .C(n11096), .D(n11085), .Y(
        n11093) );
  NAND4BBX1 U10799 ( .AN(n8174), .BN(n8175), .C(n8176), .D(n8165), .Y(n8173)
         );
  NAND4BBX1 U10800 ( .AN(n10802), .BN(n10803), .C(n10804), .D(n10793), .Y(
        n10801) );
  NAND4BBX1 U10801 ( .AN(n9050), .BN(n9051), .C(n9052), .D(n9041), .Y(n9049)
         );
  NAND4BBX1 U10802 ( .AN(n7298), .BN(n7299), .C(n7300), .D(n7289), .Y(n7297)
         );
  NAND4BBX1 U10803 ( .AN(n10218), .BN(n10219), .C(n10220), .D(n10209), .Y(
        n10217) );
  NAND4BBX1 U10804 ( .AN(n9342), .BN(n9343), .C(n9344), .D(n9333), .Y(n9341)
         );
  NAND4BBX1 U10805 ( .AN(n8466), .BN(n8467), .C(n8468), .D(n8457), .Y(n8465)
         );
  NAND4BBX1 U10806 ( .AN(n7590), .BN(n7591), .C(n7592), .D(n7581), .Y(n7589)
         );
  NAND4BBX1 U10807 ( .AN(n11386), .BN(n11387), .C(n11388), .D(n11377), .Y(
        n11385) );
  NAND4BBX1 U10808 ( .AN(n10510), .BN(n10511), .C(n10512), .D(n10501), .Y(
        n10509) );
  NAND4BBX1 U10809 ( .AN(n9634), .BN(n9635), .C(n9636), .D(n9625), .Y(n9633)
         );
  NAND4BBX1 U10810 ( .AN(n8758), .BN(n8759), .C(n8760), .D(n8749), .Y(n8757)
         );
  NAND4BBX1 U10811 ( .AN(n7882), .BN(n7883), .C(n7884), .D(n7873), .Y(n7881)
         );
  XNOR2X1 U10812 ( .A(top_core_EC_mc_mix_in_4_58_), .B(top_core_EC_mc_n441), 
        .Y(top_core_EC_mc_n365) );
  XNOR2X1 U10813 ( .A(top_core_EC_mc_mix_in_4_90_), .B(top_core_EC_mc_n173), 
        .Y(top_core_EC_mc_n106) );
  XNOR2X1 U10814 ( .A(top_core_EC_mc_mix_in_4_122_), .B(top_core_EC_mc_n35), 
        .Y(top_core_EC_mc_n760) );
  XNOR2X1 U10815 ( .A(top_core_EC_mc_mix_in_8[62]), .B(top_core_EC_mc_n408), 
        .Y(top_core_EC_mc_n332) );
  XNOR2X1 U10816 ( .A(top_core_EC_mc_mix_in_8[94]), .B(top_core_EC_mc_n149), 
        .Y(top_core_EC_mc_n73) );
  XNOR2X1 U10817 ( .A(top_core_EC_mc_mix_in_8[126]), .B(top_core_EC_mc_n808), 
        .Y(top_core_EC_mc_n738) );
  XNOR2X1 U10818 ( .A(top_core_EC_mc_mix_in_2_59_), .B(top_core_EC_mc_n416), 
        .Y(top_core_EC_mc_n349) );
  XNOR2X1 U10819 ( .A(top_core_EC_mc_mix_in_2_91_), .B(top_core_EC_mc_n157), 
        .Y(top_core_EC_mc_n81) );
  XNOR2X1 U10820 ( .A(top_core_EC_mc_mix_in_2_123_), .B(top_core_EC_mc_n17), 
        .Y(top_core_EC_mc_n746) );
  OAI22X1 U10821 ( .A0(n17119), .A1(n2851), .B0(n2854), .B1(n17120), .Y(n17117) );
  AOI21X1 U10822 ( .A0(n17060), .A1(n2905), .B0(n998), .Y(n17119) );
  OAI22X1 U10823 ( .A0(n13969), .A1(n3452), .B0(n3455), .B1(n13970), .Y(n13967) );
  AOI21X1 U10824 ( .A0(n13910), .A1(n3499), .B0(n1137), .Y(n13969) );
  OAI22X1 U10825 ( .A0(n18379), .A1(n2609), .B0(n2612), .B1(n18380), .Y(n18377) );
  AOI21X1 U10826 ( .A0(n18320), .A1(n2654), .B0(n942), .Y(n18379) );
  OAI22X1 U10827 ( .A0(n15229), .A1(n3211), .B0(n3214), .B1(n15230), .Y(n15227) );
  AOI21X1 U10828 ( .A0(n15170), .A1(n3265), .B0(n1082), .Y(n15229) );
  OAI22X1 U10829 ( .A0(n15544), .A1(n3150), .B0(n3153), .B1(n15545), .Y(n15542) );
  AOI21X1 U10830 ( .A0(n15485), .A1(n3204), .B0(n1068), .Y(n15544) );
  OAI22X1 U10831 ( .A0(n18694), .A1(n2548), .B0(n2551), .B1(n18695), .Y(n18692) );
  AOI21X1 U10832 ( .A0(n18635), .A1(n2593), .B0(n928), .Y(n18694) );
  OAI22X1 U10833 ( .A0(n16804), .A1(n2912), .B0(n2915), .B1(n16805), .Y(n16802) );
  AOI21X1 U10834 ( .A0(n16745), .A1(n2966), .B0(n1012), .Y(n16804) );
  OAI22X1 U10835 ( .A0(n14914), .A1(n3272), .B0(n3275), .B1(n14915), .Y(n14912) );
  AOI21X1 U10836 ( .A0(n14855), .A1(n3316), .B0(n1096), .Y(n14914) );
  OAI22X1 U10837 ( .A0(n16489), .A1(n2973), .B0(n2976), .B1(n16490), .Y(n16487) );
  AOI21X1 U10838 ( .A0(n16430), .A1(n3017), .B0(n1026), .Y(n16489) );
  OAI22X1 U10839 ( .A0(n18064), .A1(n2670), .B0(n2673), .B1(n18065), .Y(n18062) );
  AOI21X1 U10840 ( .A0(n18005), .A1(n2712), .B0(n956), .Y(n18064) );
  OAI22X1 U10841 ( .A0(n14599), .A1(n3333), .B0(n3336), .B1(n14600), .Y(n14597) );
  AOI21X1 U10842 ( .A0(n14540), .A1(n3377), .B0(n1110), .Y(n14599) );
  OAI22X1 U10843 ( .A0(n16174), .A1(n3031), .B0(n3034), .B1(n16175), .Y(n16172) );
  AOI21X1 U10844 ( .A0(n16115), .A1(n3076), .B0(n1040), .Y(n16174) );
  OAI22X1 U10845 ( .A0(n17749), .A1(n2730), .B0(n2733), .B1(n17750), .Y(n17747) );
  AOI21X1 U10846 ( .A0(n17690), .A1(n2775), .B0(n970), .Y(n17749) );
  OAI22X1 U10847 ( .A0(n14284), .A1(n3391), .B0(n3394), .B1(n14285), .Y(n14282) );
  AOI21X1 U10848 ( .A0(n14225), .A1(n3434), .B0(n1124), .Y(n14284) );
  OAI22X1 U10849 ( .A0(n15859), .A1(n3092), .B0(n3095), .B1(n15860), .Y(n15857) );
  AOI21X1 U10850 ( .A0(n15800), .A1(n3136), .B0(n1054), .Y(n15859) );
  OAI22X1 U10851 ( .A0(n17434), .A1(n2791), .B0(n2794), .B1(n17435), .Y(n17432) );
  AOI21X1 U10852 ( .A0(n17375), .A1(n2836), .B0(n984), .Y(n17434) );
  XNOR2X1 U10853 ( .A(n1545), .B(top_core_EC_mc_n101), .Y(top_core_EC_mc_n624)
         );
  XNOR2X1 U10854 ( .A(n1547), .B(top_core_EC_mc_n255), .Y(top_core_EC_mc_n574)
         );
  XNOR2X1 U10855 ( .A(n1546), .B(top_core_EC_mc_n190), .Y(top_core_EC_mc_n567)
         );
  NAND2XL U10856 ( .A(n73), .B(n13382), .Y(n13218) );
  NAND2XL U10857 ( .A(n75), .B(n13067), .Y(n12903) );
  NAND2XL U10858 ( .A(n74), .B(n12752), .Y(n12588) );
  AOI21X1 U10859 ( .A0(n13250), .A1(n13350), .B0(n13251), .Y(n13357) );
  CLKINVX3 U10860 ( .A(n11674), .Y(n6826) );
  CLKINVX3 U10861 ( .A(top_core_KE_sb1_n99), .Y(n6804) );
  CLKINVX3 U10862 ( .A(n13251), .Y(n6472) );
  CLKINVX3 U10863 ( .A(n11990), .Y(n6507) );
  CLKINVX3 U10864 ( .A(n12621), .Y(n6775) );
  CLKINVX3 U10865 ( .A(n13566), .Y(n6519) );
  CLKINVX3 U10866 ( .A(n12936), .Y(n6815) );
  AOI22X1 U10867 ( .A0(n1143), .A1(n561), .B0(n6174), .B1(n3498), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n323) );
  AOI22X1 U10868 ( .A0(n1001), .A1(n562), .B0(n5387), .B1(n2894), .Y(n10137)
         );
  AOI22X1 U10869 ( .A0(n945), .A1(n563), .B0(n5033), .B1(n2657), .Y(n11305) );
  AOI22X1 U10870 ( .A0(n1085), .A1(n564), .B0(n5859), .B1(n3254), .Y(n8385) );
  AOI22X1 U10871 ( .A0(n959), .A1(n565), .B0(n5117), .B1(n2713), .Y(n11013) );
  AOI22X1 U10872 ( .A0(n1043), .A1(n566), .B0(n5623), .B1(n3079), .Y(n9261) );
  AOI22X1 U10873 ( .A0(n1127), .A1(n567), .B0(n6087), .B1(n3435), .Y(n7509) );
  AOI22X1 U10874 ( .A0(n987), .A1(n568), .B0(n5303), .B1(n2837), .Y(n10429) );
  AOI22X1 U10875 ( .A0(n1029), .A1(n569), .B0(n5547), .B1(n3018), .Y(n9553) );
  AOI22X1 U10876 ( .A0(n1071), .A1(n570), .B0(n5775), .B1(n3193), .Y(n8677) );
  AOI22X1 U10877 ( .A0(n1113), .A1(n571), .B0(n6011), .B1(n3378), .Y(n7801) );
  AOI22X1 U10878 ( .A0(n931), .A1(n572), .B0(n4917), .B1(n2596), .Y(n11597) );
  AOI22X1 U10879 ( .A0(n973), .A1(n573), .B0(n5225), .B1(n2776), .Y(n10721) );
  AOI22X1 U10880 ( .A0(n1015), .A1(n574), .B0(n5471), .B1(n2955), .Y(n9845) );
  AOI22X1 U10881 ( .A0(n1057), .A1(n575), .B0(n5699), .B1(n3137), .Y(n8969) );
  AOI22X1 U10882 ( .A0(n1099), .A1(n576), .B0(n5935), .B1(n3317), .Y(n8093) );
  OAI21XL U10883 ( .A0(n1802), .A1(n11675), .B0(n11676), .Y(n11666) );
  OAI21XL U10884 ( .A0(n1823), .A1(top_core_KE_sb1_n100), .B0(
        top_core_KE_sb1_n101), .Y(top_core_KE_sb1_n91) );
  OAI21XL U10885 ( .A0(n1760), .A1(n12306), .B0(n12307), .Y(n12297) );
  OAI21XL U10886 ( .A0(n1781), .A1(n11991), .B0(n11992), .Y(n11982) );
  OAI21XL U10887 ( .A0(n1709), .A1(n12937), .B0(n12938), .Y(n12928) );
  OAI21XL U10888 ( .A0(n1651), .A1(n13567), .B0(n13568), .Y(n13558) );
  OAI21XL U10889 ( .A0(n1738), .A1(n12622), .B0(n12623), .Y(n12613) );
  AOI22X1 U10890 ( .A0(n5334), .A1(n1005), .B0(n498), .B1(n17068), .Y(n17067)
         );
  AOI22X1 U10891 ( .A0(n6117), .A1(n1144), .B0(n497), .B1(n13918), .Y(n13917)
         );
  AOI22X1 U10892 ( .A0(n4980), .A1(n949), .B0(n501), .B1(n18328), .Y(n18327)
         );
  AOI22X1 U10893 ( .A0(n5806), .A1(n1089), .B0(n500), .B1(n15178), .Y(n15177)
         );
  AOI22X1 U10894 ( .A0(n5722), .A1(n1075), .B0(n499), .B1(n15493), .Y(n15492)
         );
  AOI22X1 U10895 ( .A0(n4864), .A1(n935), .B0(n502), .B1(n18643), .Y(n18642)
         );
  AOI22X1 U10896 ( .A0(n5418), .A1(n1019), .B0(n503), .B1(n16753), .Y(n16752)
         );
  AOI22X1 U10897 ( .A0(n5882), .A1(n1103), .B0(n504), .B1(n14863), .Y(n14862)
         );
  AOI22X1 U10898 ( .A0(n5494), .A1(n1033), .B0(n505), .B1(n16438), .Y(n16437)
         );
  AOI22X1 U10899 ( .A0(n5064), .A1(n963), .B0(n506), .B1(n18013), .Y(n18012)
         );
  AOI22X1 U10900 ( .A0(n5958), .A1(n1117), .B0(n507), .B1(n14548), .Y(n14547)
         );
  AOI22X1 U10901 ( .A0(n5570), .A1(n1047), .B0(n508), .B1(n16123), .Y(n16122)
         );
  AOI22X1 U10902 ( .A0(n5172), .A1(n977), .B0(n509), .B1(n17698), .Y(n17697)
         );
  AOI22X1 U10903 ( .A0(n6034), .A1(n1131), .B0(n510), .B1(n14233), .Y(n14232)
         );
  AOI22X1 U10904 ( .A0(n5646), .A1(n1061), .B0(n511), .B1(n15808), .Y(n15807)
         );
  AOI22X1 U10905 ( .A0(n5250), .A1(n991), .B0(n512), .B1(n17383), .Y(n17382)
         );
  AOI22X1 U10906 ( .A0(n5347), .A1(n498), .B0(n481), .B1(n5387), .Y(n9983) );
  AOI22X1 U10907 ( .A0(n6143), .A1(n497), .B0(n482), .B1(n6174), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n169) );
  AOI22X1 U10908 ( .A0(n4993), .A1(n501), .B0(n483), .B1(n5033), .Y(n11151) );
  AOI22X1 U10909 ( .A0(n5819), .A1(n500), .B0(n484), .B1(n5859), .Y(n8231) );
  AOI22X1 U10910 ( .A0(n5077), .A1(n506), .B0(n485), .B1(n5117), .Y(n10859) );
  AOI22X1 U10911 ( .A0(n5583), .A1(n508), .B0(n486), .B1(n5623), .Y(n9107) );
  AOI22X1 U10912 ( .A0(n6047), .A1(n510), .B0(n487), .B1(n6087), .Y(n7355) );
  AOI22X1 U10913 ( .A0(n5263), .A1(n512), .B0(n488), .B1(n5303), .Y(n10275) );
  AOI22X1 U10914 ( .A0(n5507), .A1(n505), .B0(n489), .B1(n5547), .Y(n9399) );
  AOI22X1 U10915 ( .A0(n5735), .A1(n499), .B0(n490), .B1(n5775), .Y(n8523) );
  AOI22X1 U10916 ( .A0(n5971), .A1(n507), .B0(n491), .B1(n6011), .Y(n7647) );
  AOI22X1 U10917 ( .A0(n4877), .A1(n502), .B0(n492), .B1(n4917), .Y(n11443) );
  AOI22X1 U10918 ( .A0(n5185), .A1(n509), .B0(n493), .B1(n5225), .Y(n10567) );
  AOI22X1 U10919 ( .A0(n5431), .A1(n503), .B0(n494), .B1(n5471), .Y(n9691) );
  AOI22X1 U10920 ( .A0(n5659), .A1(n511), .B0(n495), .B1(n5699), .Y(n8815) );
  AOI22X1 U10921 ( .A0(n5895), .A1(n504), .B0(n496), .B1(n5935), .Y(n7939) );
  AOI22X1 U10922 ( .A0(n2846), .A1(n17111), .B0(n17112), .B1(n2849), .Y(n17103) );
  NAND4X1 U10923 ( .A(n17113), .B(n17114), .C(n17115), .D(n17116), .Y(n17112)
         );
  OAI221XL U10924 ( .A0(n17123), .A1(n17030), .B0(n17124), .B1(n2853), .C0(
        n17125), .Y(n17111) );
  AOI22X1 U10925 ( .A0(n3447), .A1(n13961), .B0(n13962), .B1(n3449), .Y(n13953) );
  NAND4X1 U10926 ( .A(n13963), .B(n13964), .C(n13965), .D(n13966), .Y(n13962)
         );
  OAI221XL U10927 ( .A0(n13973), .A1(n13880), .B0(n13974), .B1(n3454), .C0(
        n13975), .Y(n13961) );
  AOI22X1 U10928 ( .A0(n2604), .A1(n18371), .B0(n18372), .B1(n2607), .Y(n18363) );
  NAND4X1 U10929 ( .A(n18373), .B(n18374), .C(n18375), .D(n18376), .Y(n18372)
         );
  OAI221XL U10930 ( .A0(n18383), .A1(n18290), .B0(n18384), .B1(n2611), .C0(
        n18385), .Y(n18371) );
  AOI22X1 U10931 ( .A0(n3206), .A1(n15221), .B0(n15222), .B1(n3209), .Y(n15213) );
  NAND4X1 U10932 ( .A(n15223), .B(n15224), .C(n15225), .D(n15226), .Y(n15222)
         );
  OAI221XL U10933 ( .A0(n15233), .A1(n15140), .B0(n15234), .B1(n3213), .C0(
        n15235), .Y(n15221) );
  AOI22X1 U10934 ( .A0(n3145), .A1(n15536), .B0(n15537), .B1(n3148), .Y(n15528) );
  NAND4X1 U10935 ( .A(n15538), .B(n15539), .C(n15540), .D(n15541), .Y(n15537)
         );
  OAI221XL U10936 ( .A0(n15548), .A1(n15455), .B0(n15549), .B1(n3152), .C0(
        n15550), .Y(n15536) );
  AOI22X1 U10937 ( .A0(n2543), .A1(n18686), .B0(n18687), .B1(n2546), .Y(n18678) );
  NAND4X1 U10938 ( .A(n18688), .B(n18689), .C(n18690), .D(n18691), .Y(n18687)
         );
  OAI221XL U10939 ( .A0(n18698), .A1(n18605), .B0(n18699), .B1(n2550), .C0(
        n18700), .Y(n18686) );
  AOI22X1 U10940 ( .A0(n2907), .A1(n16796), .B0(n16797), .B1(n2910), .Y(n16788) );
  NAND4X1 U10941 ( .A(n16798), .B(n16799), .C(n16800), .D(n16801), .Y(n16797)
         );
  OAI221XL U10942 ( .A0(n16808), .A1(n16715), .B0(n16809), .B1(n2914), .C0(
        n16810), .Y(n16796) );
  AOI22X1 U10943 ( .A0(n3267), .A1(n14906), .B0(n14907), .B1(n3270), .Y(n14898) );
  NAND4X1 U10944 ( .A(n14908), .B(n14909), .C(n14910), .D(n14911), .Y(n14907)
         );
  OAI221XL U10945 ( .A0(n14918), .A1(n14825), .B0(n14919), .B1(n3274), .C0(
        n14920), .Y(n14906) );
  AOI22X1 U10946 ( .A0(n2968), .A1(n16481), .B0(n16482), .B1(n2971), .Y(n16473) );
  NAND4X1 U10947 ( .A(n16483), .B(n16484), .C(n16485), .D(n16486), .Y(n16482)
         );
  OAI221XL U10948 ( .A0(n16493), .A1(n16400), .B0(n16494), .B1(n2975), .C0(
        n16495), .Y(n16481) );
  AOI22X1 U10949 ( .A0(n2665), .A1(n18056), .B0(n18057), .B1(n2668), .Y(n18048) );
  NAND4X1 U10950 ( .A(n18058), .B(n18059), .C(n18060), .D(n18061), .Y(n18057)
         );
  OAI221XL U10951 ( .A0(n18068), .A1(n17975), .B0(n18069), .B1(n2672), .C0(
        n18070), .Y(n18056) );
  AOI22X1 U10952 ( .A0(n3328), .A1(n14591), .B0(n14592), .B1(n3331), .Y(n14583) );
  NAND4X1 U10953 ( .A(n14593), .B(n14594), .C(n14595), .D(n14596), .Y(n14592)
         );
  OAI221XL U10954 ( .A0(n14603), .A1(n14510), .B0(n14604), .B1(n3335), .C0(
        n14605), .Y(n14591) );
  AOI22X1 U10955 ( .A0(n3026), .A1(n16166), .B0(n16167), .B1(n3029), .Y(n16158) );
  NAND4X1 U10956 ( .A(n16168), .B(n16169), .C(n16170), .D(n16171), .Y(n16167)
         );
  OAI221XL U10957 ( .A0(n16178), .A1(n16085), .B0(n16179), .B1(n3033), .C0(
        n16180), .Y(n16166) );
  AOI22X1 U10958 ( .A0(n2725), .A1(n17741), .B0(n17742), .B1(n2728), .Y(n17733) );
  NAND4X1 U10959 ( .A(n17743), .B(n17744), .C(n17745), .D(n17746), .Y(n17742)
         );
  OAI221XL U10960 ( .A0(n17753), .A1(n17660), .B0(n17754), .B1(n2732), .C0(
        n17755), .Y(n17741) );
  AOI22X1 U10961 ( .A0(n3386), .A1(n14276), .B0(n14277), .B1(n3389), .Y(n14268) );
  NAND4X1 U10962 ( .A(n14278), .B(n14279), .C(n14280), .D(n14281), .Y(n14277)
         );
  OAI221XL U10963 ( .A0(n14288), .A1(n14195), .B0(n14289), .B1(n3393), .C0(
        n14290), .Y(n14276) );
  AOI22X1 U10964 ( .A0(n3087), .A1(n15851), .B0(n15852), .B1(n3090), .Y(n15843) );
  NAND4X1 U10965 ( .A(n15853), .B(n15854), .C(n15855), .D(n15856), .Y(n15852)
         );
  OAI221XL U10966 ( .A0(n15863), .A1(n15770), .B0(n15864), .B1(n3094), .C0(
        n15865), .Y(n15851) );
  AOI22X1 U10967 ( .A0(n2786), .A1(n17426), .B0(n17427), .B1(n2789), .Y(n17418) );
  NAND4X1 U10968 ( .A(n17428), .B(n17429), .C(n17430), .D(n17431), .Y(n17427)
         );
  OAI221XL U10969 ( .A0(n17438), .A1(n17345), .B0(n17439), .B1(n2793), .C0(
        n17440), .Y(n17426) );
  AOI21XL U10970 ( .A0(n11705), .A1(n6920), .B0(n11741), .Y(n11863) );
  AOI21XL U10971 ( .A0(top_core_KE_sb1_n130), .A1(n6874), .B0(
        top_core_KE_sb1_n168), .Y(top_core_KE_sb1_n292) );
  AOI21XL U10972 ( .A0(n12336), .A1(n6627), .B0(n12372), .Y(n12494) );
  AOI21XL U10973 ( .A0(n12021), .A1(n6580), .B0(n12057), .Y(n12179) );
  AOI21XL U10974 ( .A0(n12652), .A1(n6851), .B0(n12688), .Y(n12809) );
  AOI21XL U10975 ( .A0(n13597), .A1(n6604), .B0(n13633), .Y(n13754) );
  AOI21XL U10976 ( .A0(n12967), .A1(n6897), .B0(n13003), .Y(n13124) );
  OAI21XL U10977 ( .A0(n9941), .A1(n9942), .B0(n2852), .Y(n9940) );
  NAND4X1 U10978 ( .A(n9947), .B(n9948), .C(n9949), .D(n9950), .Y(n9941) );
  OAI222XL U10979 ( .A0(n9943), .A1(n9891), .B0(n2899), .B1(n9944), .C0(n9945), 
        .C1(n9946), .Y(n9942) );
  OAI21XL U10980 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n126), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n127), .B0(n3453), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n125) );
  NAND4X1 U10981 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n132), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n133), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n134), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n135), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n126) );
  OAI222XL U10982 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n128), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n74), .B0(n3500), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n129), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n130), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n131), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n127) );
  OAI21XL U10983 ( .A0(n11109), .A1(n11110), .B0(n2610), .Y(n11108) );
  NAND4X1 U10984 ( .A(n11115), .B(n11116), .C(n11117), .D(n11118), .Y(n11109)
         );
  OAI222XL U10985 ( .A0(n11111), .A1(n11059), .B0(n2656), .B1(n11112), .C0(
        n11113), .C1(n11114), .Y(n11110) );
  OAI21XL U10986 ( .A0(n8189), .A1(n8190), .B0(n3212), .Y(n8188) );
  NAND4X1 U10987 ( .A(n8195), .B(n8196), .C(n8197), .D(n8198), .Y(n8189) );
  OAI222XL U10988 ( .A0(n8191), .A1(n8139), .B0(n3259), .B1(n8192), .C0(n8193), 
        .C1(n8194), .Y(n8190) );
  OAI21XL U10989 ( .A0(n10817), .A1(n10818), .B0(n2671), .Y(n10816) );
  NAND4X1 U10990 ( .A(n10823), .B(n10824), .C(n10825), .D(n10826), .Y(n10817)
         );
  OAI222XL U10991 ( .A0(n10819), .A1(n10767), .B0(n2717), .B1(n10820), .C0(
        n10821), .C1(n10822), .Y(n10818) );
  OAI21XL U10992 ( .A0(n9065), .A1(n9066), .B0(n3032), .Y(n9064) );
  NAND4X1 U10993 ( .A(n9071), .B(n9072), .C(n9073), .D(n9074), .Y(n9065) );
  OAI222XL U10994 ( .A0(n9067), .A1(n9015), .B0(n3078), .B1(n9068), .C0(n9069), 
        .C1(n9070), .Y(n9066) );
  OAI21XL U10995 ( .A0(n7313), .A1(n7314), .B0(n3392), .Y(n7312) );
  NAND4X1 U10996 ( .A(n7319), .B(n7320), .C(n7321), .D(n7322), .Y(n7313) );
  OAI222XL U10997 ( .A0(n7315), .A1(n7263), .B0(n3439), .B1(n7316), .C0(n7317), 
        .C1(n7318), .Y(n7314) );
  OAI21XL U10998 ( .A0(n10233), .A1(n10234), .B0(n2792), .Y(n10232) );
  NAND4X1 U10999 ( .A(n10239), .B(n10240), .C(n10241), .D(n10242), .Y(n10233)
         );
  OAI222XL U11000 ( .A0(n10235), .A1(n10183), .B0(n2842), .B1(n10236), .C0(
        n10237), .C1(n10238), .Y(n10234) );
  OAI21XL U11001 ( .A0(n9357), .A1(n9358), .B0(n2974), .Y(n9356) );
  NAND4X1 U11002 ( .A(n9363), .B(n9364), .C(n9365), .D(n9366), .Y(n9357) );
  OAI222XL U11003 ( .A0(n9359), .A1(n9307), .B0(n3019), .B1(n9360), .C0(n9361), 
        .C1(n9362), .Y(n9358) );
  OAI21XL U11004 ( .A0(n8481), .A1(n8482), .B0(n3151), .Y(n8480) );
  NAND4X1 U11005 ( .A(n8487), .B(n8488), .C(n8489), .D(n8490), .Y(n8481) );
  OAI222XL U11006 ( .A0(n8483), .A1(n8431), .B0(n3198), .B1(n8484), .C0(n8485), 
        .C1(n8486), .Y(n8482) );
  OAI21XL U11007 ( .A0(n7605), .A1(n7606), .B0(n3334), .Y(n7604) );
  NAND4X1 U11008 ( .A(n7611), .B(n7612), .C(n7613), .D(n7614), .Y(n7605) );
  OAI222XL U11009 ( .A0(n7607), .A1(n7555), .B0(n3379), .B1(n7608), .C0(n7609), 
        .C1(n7610), .Y(n7606) );
  OAI21XL U11010 ( .A0(n11401), .A1(n11402), .B0(n2549), .Y(n11400) );
  NAND4X1 U11011 ( .A(n11407), .B(n11408), .C(n11409), .D(n11410), .Y(n11401)
         );
  OAI222XL U11012 ( .A0(n11403), .A1(n11351), .B0(n2595), .B1(n11404), .C0(
        n11405), .C1(n11406), .Y(n11402) );
  OAI21XL U11013 ( .A0(n10525), .A1(n10526), .B0(n2731), .Y(n10524) );
  NAND4X1 U11014 ( .A(n10531), .B(n10532), .C(n10533), .D(n10534), .Y(n10525)
         );
  OAI222XL U11015 ( .A0(n10527), .A1(n10475), .B0(n2774), .B1(n10528), .C0(
        n10529), .C1(n10530), .Y(n10526) );
  OAI21XL U11016 ( .A0(n9649), .A1(n9650), .B0(n2913), .Y(n9648) );
  NAND4X1 U11017 ( .A(n9655), .B(n9656), .C(n9657), .D(n9658), .Y(n9649) );
  OAI222XL U11018 ( .A0(n9651), .A1(n9599), .B0(n2960), .B1(n9652), .C0(n9653), 
        .C1(n9654), .Y(n9650) );
  OAI21XL U11019 ( .A0(n8773), .A1(n8774), .B0(n3093), .Y(n8772) );
  NAND4X1 U11020 ( .A(n8779), .B(n8780), .C(n8781), .D(n8782), .Y(n8773) );
  OAI222XL U11021 ( .A0(n8775), .A1(n8723), .B0(n3138), .B1(n8776), .C0(n8777), 
        .C1(n8778), .Y(n8774) );
  OAI21XL U11022 ( .A0(n7897), .A1(n7898), .B0(n3273), .Y(n7896) );
  NAND4X1 U11023 ( .A(n7903), .B(n7904), .C(n7905), .D(n7906), .Y(n7897) );
  OAI222XL U11024 ( .A0(n7899), .A1(n7847), .B0(n3322), .B1(n7900), .C0(n7901), 
        .C1(n7902), .Y(n7898) );
  AOI21X1 U11025 ( .A0(n3447), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n61), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n62), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n60) );
  AOI31X1 U11026 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n63), .A1(n6158), 
        .A2(top_core_EC_ss_gen_tbox_0__sboxs_r_n64), .B0(n3448), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n62) );
  OAI222XL U11027 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n78), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n80), .B1(n3454), .C0(n3461), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n81), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n61) );
  INVX1 U11028 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n75), .Y(n6158) );
  AOI21X1 U11029 ( .A0(n2846), .A1(n9879), .B0(n9880), .Y(n9878) );
  AOI31X1 U11030 ( .A0(n9881), .A1(n5368), .A2(n9882), .B0(n2847), .Y(n9880)
         );
  OAI222XL U11031 ( .A0(n9895), .A1(n9896), .B0(n9897), .B1(n2853), .C0(n2860), 
        .C1(n9898), .Y(n9879) );
  INVX1 U11032 ( .A(n9892), .Y(n5368) );
  AOI21X1 U11033 ( .A0(n2604), .A1(n11047), .B0(n11048), .Y(n11046) );
  AOI31X1 U11034 ( .A0(n11049), .A1(n5014), .A2(n11050), .B0(n2605), .Y(n11048) );
  OAI222XL U11035 ( .A0(n11063), .A1(n11064), .B0(n11065), .B1(n2611), .C0(
        n2618), .C1(n11066), .Y(n11047) );
  INVX1 U11036 ( .A(n11060), .Y(n5014) );
  AOI21X1 U11037 ( .A0(n3206), .A1(n8127), .B0(n8128), .Y(n8126) );
  AOI31X1 U11038 ( .A0(n8129), .A1(n5840), .A2(n8130), .B0(n3207), .Y(n8128)
         );
  OAI222XL U11039 ( .A0(n8143), .A1(n8144), .B0(n8145), .B1(n3213), .C0(n3220), 
        .C1(n8146), .Y(n8127) );
  INVX1 U11040 ( .A(n8140), .Y(n5840) );
  AOI21X1 U11041 ( .A0(n2665), .A1(n10755), .B0(n10756), .Y(n10754) );
  AOI31X1 U11042 ( .A0(n10757), .A1(n5098), .A2(n10758), .B0(n2666), .Y(n10756) );
  OAI222XL U11043 ( .A0(n10771), .A1(n10772), .B0(n10773), .B1(n2672), .C0(
        n2679), .C1(n10774), .Y(n10755) );
  INVX1 U11044 ( .A(n10768), .Y(n5098) );
  AOI21X1 U11045 ( .A0(n3026), .A1(n9003), .B0(n9004), .Y(n9002) );
  AOI31X1 U11046 ( .A0(n9005), .A1(n5604), .A2(n9006), .B0(n3027), .Y(n9004)
         );
  OAI222XL U11047 ( .A0(n9019), .A1(n9020), .B0(n9021), .B1(n3033), .C0(n3040), 
        .C1(n9022), .Y(n9003) );
  INVX1 U11048 ( .A(n9016), .Y(n5604) );
  AOI21X1 U11049 ( .A0(n3386), .A1(n7251), .B0(n7252), .Y(n7250) );
  AOI31X1 U11050 ( .A0(n7253), .A1(n6068), .A2(n7254), .B0(n3387), .Y(n7252)
         );
  OAI222XL U11051 ( .A0(n7267), .A1(n7268), .B0(n7269), .B1(n3393), .C0(n3400), 
        .C1(n7270), .Y(n7251) );
  INVX1 U11052 ( .A(n7264), .Y(n6068) );
  AOI21X1 U11053 ( .A0(n2786), .A1(n10171), .B0(n10172), .Y(n10170) );
  AOI31X1 U11054 ( .A0(n10173), .A1(n5284), .A2(n10174), .B0(n2787), .Y(n10172) );
  OAI222XL U11055 ( .A0(n10187), .A1(n10188), .B0(n10189), .B1(n2793), .C0(
        n2800), .C1(n10190), .Y(n10171) );
  INVX1 U11056 ( .A(n10184), .Y(n5284) );
  AOI21X1 U11057 ( .A0(n2968), .A1(n9295), .B0(n9296), .Y(n9294) );
  AOI31X1 U11058 ( .A0(n9297), .A1(n5528), .A2(n9298), .B0(n2969), .Y(n9296)
         );
  OAI222XL U11059 ( .A0(n9311), .A1(n9312), .B0(n9313), .B1(n2975), .C0(n2982), 
        .C1(n9314), .Y(n9295) );
  INVX1 U11060 ( .A(n9308), .Y(n5528) );
  AOI21X1 U11061 ( .A0(n3145), .A1(n8419), .B0(n8420), .Y(n8418) );
  AOI31X1 U11062 ( .A0(n8421), .A1(n5756), .A2(n8422), .B0(n3146), .Y(n8420)
         );
  OAI222XL U11063 ( .A0(n8435), .A1(n8436), .B0(n8437), .B1(n3152), .C0(n3159), 
        .C1(n8438), .Y(n8419) );
  INVX1 U11064 ( .A(n8432), .Y(n5756) );
  AOI21X1 U11065 ( .A0(n3328), .A1(n7543), .B0(n7544), .Y(n7542) );
  AOI31X1 U11066 ( .A0(n7545), .A1(n5992), .A2(n7546), .B0(n3329), .Y(n7544)
         );
  OAI222XL U11067 ( .A0(n7559), .A1(n7560), .B0(n7561), .B1(n3335), .C0(n3342), 
        .C1(n7562), .Y(n7543) );
  INVX1 U11068 ( .A(n7556), .Y(n5992) );
  AOI21X1 U11069 ( .A0(n2543), .A1(n11339), .B0(n11340), .Y(n11338) );
  AOI31X1 U11070 ( .A0(n11341), .A1(n4898), .A2(n11342), .B0(n2544), .Y(n11340) );
  OAI222XL U11071 ( .A0(n11355), .A1(n11356), .B0(n11357), .B1(n2550), .C0(
        n2557), .C1(n11358), .Y(n11339) );
  INVX1 U11072 ( .A(n11352), .Y(n4898) );
  AOI21X1 U11073 ( .A0(n2725), .A1(n10463), .B0(n10464), .Y(n10462) );
  AOI31X1 U11074 ( .A0(n10465), .A1(n5206), .A2(n10466), .B0(n2726), .Y(n10464) );
  OAI222XL U11075 ( .A0(n10479), .A1(n10480), .B0(n10481), .B1(n2732), .C0(
        n2739), .C1(n10482), .Y(n10463) );
  INVX1 U11076 ( .A(n10476), .Y(n5206) );
  AOI21X1 U11077 ( .A0(n2907), .A1(n9587), .B0(n9588), .Y(n9586) );
  AOI31X1 U11078 ( .A0(n9589), .A1(n5452), .A2(n9590), .B0(n2908), .Y(n9588)
         );
  OAI222XL U11079 ( .A0(n9603), .A1(n9604), .B0(n9605), .B1(n2914), .C0(n2921), 
        .C1(n9606), .Y(n9587) );
  INVX1 U11080 ( .A(n9600), .Y(n5452) );
  AOI21X1 U11081 ( .A0(n3087), .A1(n8711), .B0(n8712), .Y(n8710) );
  AOI31X1 U11082 ( .A0(n8713), .A1(n5680), .A2(n8714), .B0(n3088), .Y(n8712)
         );
  OAI222XL U11083 ( .A0(n8727), .A1(n8728), .B0(n8729), .B1(n3094), .C0(n3101), 
        .C1(n8730), .Y(n8711) );
  INVX1 U11084 ( .A(n8724), .Y(n5680) );
  AOI21X1 U11085 ( .A0(n3267), .A1(n7835), .B0(n7836), .Y(n7834) );
  AOI31X1 U11086 ( .A0(n7837), .A1(n5916), .A2(n7838), .B0(n3268), .Y(n7836)
         );
  OAI222XL U11087 ( .A0(n7851), .A1(n7852), .B0(n7853), .B1(n3274), .C0(n3281), 
        .C1(n7854), .Y(n7835) );
  INVX1 U11088 ( .A(n7848), .Y(n5916) );
  AOI22X1 U11089 ( .A0(n9965), .A1(n2851), .B0(n2855), .B1(n9966), .Y(n9933)
         );
  NAND4X1 U11090 ( .A(n9885), .B(n9944), .C(n9968), .D(n9969), .Y(n9965) );
  NAND4X1 U11091 ( .A(n9958), .B(n9887), .C(n9930), .D(n9967), .Y(n9966) );
  AOI22X1 U11092 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n150), .A1(n3452), 
        .B0(n3456), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n151), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n118) );
  NAND4X1 U11093 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n67), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n129), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n154), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n155), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n150) );
  NAND4X1 U11094 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n143), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n69), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n115), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n152), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n151) );
  AOI22X1 U11095 ( .A0(n11133), .A1(n2609), .B0(n2613), .B1(n11134), .Y(n11101) );
  NAND4X1 U11096 ( .A(n11053), .B(n11112), .C(n11136), .D(n11137), .Y(n11133)
         );
  NAND4X1 U11097 ( .A(n11126), .B(n11055), .C(n11098), .D(n11135), .Y(n11134)
         );
  AOI22X1 U11098 ( .A0(n8213), .A1(n3211), .B0(n3215), .B1(n8214), .Y(n8181)
         );
  NAND4X1 U11099 ( .A(n8133), .B(n8192), .C(n8216), .D(n8217), .Y(n8213) );
  NAND4X1 U11100 ( .A(n8206), .B(n8135), .C(n8178), .D(n8215), .Y(n8214) );
  AOI22X1 U11101 ( .A0(n10841), .A1(n2670), .B0(n2674), .B1(n10842), .Y(n10809) );
  NAND4X1 U11102 ( .A(n10761), .B(n10820), .C(n10844), .D(n10845), .Y(n10841)
         );
  NAND4X1 U11103 ( .A(n10834), .B(n10763), .C(n10806), .D(n10843), .Y(n10842)
         );
  AOI22X1 U11104 ( .A0(n9089), .A1(n3031), .B0(n3035), .B1(n9090), .Y(n9057)
         );
  NAND4X1 U11105 ( .A(n9009), .B(n9068), .C(n9092), .D(n9093), .Y(n9089) );
  NAND4X1 U11106 ( .A(n9082), .B(n9011), .C(n9054), .D(n9091), .Y(n9090) );
  AOI22X1 U11107 ( .A0(n7337), .A1(n3391), .B0(n3395), .B1(n7338), .Y(n7305)
         );
  NAND4X1 U11108 ( .A(n7257), .B(n7316), .C(n7340), .D(n7341), .Y(n7337) );
  NAND4X1 U11109 ( .A(n7330), .B(n7259), .C(n7302), .D(n7339), .Y(n7338) );
  AOI22X1 U11110 ( .A0(n10257), .A1(n2791), .B0(n2795), .B1(n10258), .Y(n10225) );
  NAND4X1 U11111 ( .A(n10177), .B(n10236), .C(n10260), .D(n10261), .Y(n10257)
         );
  NAND4X1 U11112 ( .A(n10250), .B(n10179), .C(n10222), .D(n10259), .Y(n10258)
         );
  AOI22X1 U11113 ( .A0(n9381), .A1(n2973), .B0(n2977), .B1(n9382), .Y(n9349)
         );
  NAND4X1 U11114 ( .A(n9301), .B(n9360), .C(n9384), .D(n9385), .Y(n9381) );
  NAND4X1 U11115 ( .A(n9374), .B(n9303), .C(n9346), .D(n9383), .Y(n9382) );
  AOI22X1 U11116 ( .A0(n8505), .A1(n3150), .B0(n3154), .B1(n8506), .Y(n8473)
         );
  NAND4X1 U11117 ( .A(n8425), .B(n8484), .C(n8508), .D(n8509), .Y(n8505) );
  NAND4X1 U11118 ( .A(n8498), .B(n8427), .C(n8470), .D(n8507), .Y(n8506) );
  AOI22X1 U11119 ( .A0(n7629), .A1(n3333), .B0(n3337), .B1(n7630), .Y(n7597)
         );
  NAND4X1 U11120 ( .A(n7549), .B(n7608), .C(n7632), .D(n7633), .Y(n7629) );
  NAND4X1 U11121 ( .A(n7622), .B(n7551), .C(n7594), .D(n7631), .Y(n7630) );
  AOI22X1 U11122 ( .A0(n11425), .A1(n2548), .B0(n2552), .B1(n11426), .Y(n11393) );
  NAND4X1 U11123 ( .A(n11345), .B(n11404), .C(n11428), .D(n11429), .Y(n11425)
         );
  NAND4X1 U11124 ( .A(n11418), .B(n11347), .C(n11390), .D(n11427), .Y(n11426)
         );
  AOI22X1 U11125 ( .A0(n10549), .A1(n2730), .B0(n2734), .B1(n10550), .Y(n10517) );
  NAND4X1 U11126 ( .A(n10469), .B(n10528), .C(n10552), .D(n10553), .Y(n10549)
         );
  NAND4X1 U11127 ( .A(n10542), .B(n10471), .C(n10514), .D(n10551), .Y(n10550)
         );
  AOI22X1 U11128 ( .A0(n9673), .A1(n2912), .B0(n2916), .B1(n9674), .Y(n9641)
         );
  NAND4X1 U11129 ( .A(n9593), .B(n9652), .C(n9676), .D(n9677), .Y(n9673) );
  NAND4X1 U11130 ( .A(n9666), .B(n9595), .C(n9638), .D(n9675), .Y(n9674) );
  AOI22X1 U11131 ( .A0(n8797), .A1(n3092), .B0(n3096), .B1(n8798), .Y(n8765)
         );
  NAND4X1 U11132 ( .A(n8717), .B(n8776), .C(n8800), .D(n8801), .Y(n8797) );
  NAND4X1 U11133 ( .A(n8790), .B(n8719), .C(n8762), .D(n8799), .Y(n8798) );
  AOI22X1 U11134 ( .A0(n7921), .A1(n3272), .B0(n3276), .B1(n7922), .Y(n7889)
         );
  NAND4X1 U11135 ( .A(n7841), .B(n7900), .C(n7924), .D(n7925), .Y(n7921) );
  NAND4X1 U11136 ( .A(n7914), .B(n7843), .C(n7886), .D(n7923), .Y(n7922) );
  AOI22XL U11137 ( .A0(n6539), .A1(n1173), .B0(n6549), .B1(n1275), .Y(n13473)
         );
  AOI22XL U11138 ( .A0(n6834), .A1(n1213), .B0(n6844), .B1(n12652), .Y(n12843)
         );
  AOI22XL U11139 ( .A0(n6587), .A1(n1178), .B0(n6597), .B1(n13597), .Y(n13788)
         );
  AOI22XL U11140 ( .A0(n6880), .A1(n1219), .B0(n6890), .B1(n12967), .Y(n13158)
         );
  OAI21XL U11141 ( .A0(n1680), .A1(n73), .B0(n13246), .Y(n13320) );
  OAI21XL U11142 ( .A0(n1738), .A1(n74), .B0(n12616), .Y(n12690) );
  OAI21XL U11143 ( .A0(n1709), .A1(n75), .B0(n12931), .Y(n13005) );
  NAND2X1 U11144 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n131), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n254), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n298) );
  NAND2X1 U11145 ( .A(n9946), .B(n10068), .Y(n10112) );
  NAND2X1 U11146 ( .A(n8194), .B(n8316), .Y(n8360) );
  NAND2X1 U11147 ( .A(n11114), .B(n11236), .Y(n11280) );
  NAND2X1 U11148 ( .A(n10822), .B(n10944), .Y(n10988) );
  NAND2X1 U11149 ( .A(n7318), .B(n7440), .Y(n7484) );
  NAND2X1 U11150 ( .A(n9070), .B(n9192), .Y(n9236) );
  NAND2X1 U11151 ( .A(n10238), .B(n10360), .Y(n10404) );
  NAND2X1 U11152 ( .A(n9362), .B(n9484), .Y(n9528) );
  NAND2X1 U11153 ( .A(n8486), .B(n8608), .Y(n8652) );
  NAND2X1 U11154 ( .A(n7610), .B(n7732), .Y(n7776) );
  NAND2X1 U11155 ( .A(n11406), .B(n11528), .Y(n11572) );
  NAND2X1 U11156 ( .A(n10530), .B(n10652), .Y(n10696) );
  NAND2X1 U11157 ( .A(n9654), .B(n9776), .Y(n9820) );
  NAND2X1 U11158 ( .A(n8778), .B(n8900), .Y(n8944) );
  NAND2X1 U11159 ( .A(n7902), .B(n8024), .Y(n8068) );
  AOI21X1 U11160 ( .A0(n6627), .A1(n691), .B0(n6620), .Y(n12554) );
  AOI21XL U11161 ( .A0(n17065), .A1(n17126), .B0(n5391), .Y(n17286) );
  INVX1 U11162 ( .A(n17224), .Y(n5391) );
  AOI21XL U11163 ( .A0(n13915), .A1(n13976), .B0(n6173), .Y(n14136) );
  INVX1 U11164 ( .A(n14074), .Y(n6173) );
  AOI21XL U11165 ( .A0(n15175), .A1(n15236), .B0(n5863), .Y(n15396) );
  INVX1 U11166 ( .A(n15334), .Y(n5863) );
  AOI21XL U11167 ( .A0(n18325), .A1(n18386), .B0(n5037), .Y(n18546) );
  INVX1 U11168 ( .A(n18484), .Y(n5037) );
  AOI21XL U11169 ( .A0(n15490), .A1(n15551), .B0(n5779), .Y(n15711) );
  INVX1 U11170 ( .A(n15649), .Y(n5779) );
  AOI21XL U11171 ( .A0(n16750), .A1(n16811), .B0(n5475), .Y(n16971) );
  INVX1 U11172 ( .A(n16909), .Y(n5475) );
  AOI21XL U11173 ( .A0(n18640), .A1(n18701), .B0(n4921), .Y(n18861) );
  INVX1 U11174 ( .A(n18799), .Y(n4921) );
  AOI21XL U11175 ( .A0(n14860), .A1(n14921), .B0(n5939), .Y(n15081) );
  INVX1 U11176 ( .A(n15019), .Y(n5939) );
  AOI21XL U11177 ( .A0(n16435), .A1(n16496), .B0(n5551), .Y(n16656) );
  INVX1 U11178 ( .A(n16594), .Y(n5551) );
  AOI21XL U11179 ( .A0(n18010), .A1(n18071), .B0(n5121), .Y(n18231) );
  INVX1 U11180 ( .A(n18169), .Y(n5121) );
  AOI21XL U11181 ( .A0(n14545), .A1(n14606), .B0(n6015), .Y(n14766) );
  INVX1 U11182 ( .A(n14704), .Y(n6015) );
  AOI21XL U11183 ( .A0(n16120), .A1(n16181), .B0(n5627), .Y(n16341) );
  INVX1 U11184 ( .A(n16279), .Y(n5627) );
  AOI21XL U11185 ( .A0(n17695), .A1(n17756), .B0(n5229), .Y(n17916) );
  INVX1 U11186 ( .A(n17854), .Y(n5229) );
  AOI21XL U11187 ( .A0(n14230), .A1(n14291), .B0(n6091), .Y(n14451) );
  INVX1 U11188 ( .A(n14389), .Y(n6091) );
  AOI21XL U11189 ( .A0(n15805), .A1(n15866), .B0(n5703), .Y(n16026) );
  INVX1 U11190 ( .A(n15964), .Y(n5703) );
  AOI21XL U11191 ( .A0(n17380), .A1(n17441), .B0(n5307), .Y(n17601) );
  INVX1 U11192 ( .A(n17539), .Y(n5307) );
  AOI2BB2X1 U11193 ( .B0(n1139), .B1(n6119), .A0N(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n76), .A1N(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n77), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n63) );
  AOI2BB2X1 U11194 ( .B0(n996), .B1(n5333), .A0N(n9893), .A1N(n9894), .Y(n9881) );
  AOI2BB2X1 U11195 ( .B0(n940), .B1(n4979), .A0N(n11061), .A1N(n11062), .Y(
        n11049) );
  AOI2BB2X1 U11196 ( .B0(n1080), .B1(n5805), .A0N(n8141), .A1N(n8142), .Y(
        n8129) );
  AOI2BB2X1 U11197 ( .B0(n954), .B1(n5063), .A0N(n10769), .A1N(n10770), .Y(
        n10757) );
  AOI2BB2X1 U11198 ( .B0(n1038), .B1(n5569), .A0N(n9017), .A1N(n9018), .Y(
        n9005) );
  AOI2BB2X1 U11199 ( .B0(n1122), .B1(n6033), .A0N(n7265), .A1N(n7266), .Y(
        n7253) );
  AOI2BB2X1 U11200 ( .B0(n982), .B1(n5249), .A0N(n10185), .A1N(n10186), .Y(
        n10173) );
  AOI2BB2X1 U11201 ( .B0(n1024), .B1(n5493), .A0N(n9309), .A1N(n9310), .Y(
        n9297) );
  AOI2BB2X1 U11202 ( .B0(n1066), .B1(n5721), .A0N(n8433), .A1N(n8434), .Y(
        n8421) );
  AOI2BB2X1 U11203 ( .B0(n1108), .B1(n5957), .A0N(n7557), .A1N(n7558), .Y(
        n7545) );
  AOI2BB2X1 U11204 ( .B0(n926), .B1(n4863), .A0N(n11353), .A1N(n11354), .Y(
        n11341) );
  AOI2BB2X1 U11205 ( .B0(n968), .B1(n5171), .A0N(n10477), .A1N(n10478), .Y(
        n10465) );
  AOI2BB2X1 U11206 ( .B0(n1010), .B1(n5417), .A0N(n9601), .A1N(n9602), .Y(
        n9589) );
  AOI2BB2X1 U11207 ( .B0(n1052), .B1(n5645), .A0N(n8725), .A1N(n8726), .Y(
        n8713) );
  AOI2BB2X1 U11208 ( .B0(n1094), .B1(n5881), .A0N(n7849), .A1N(n7850), .Y(
        n7837) );
  INVX1 U11209 ( .A(n17205), .Y(n5385) );
  INVX1 U11210 ( .A(n14055), .Y(n6167) );
  INVX1 U11211 ( .A(n18465), .Y(n5031) );
  INVX1 U11212 ( .A(n15315), .Y(n5857) );
  INVX1 U11213 ( .A(n15630), .Y(n5773) );
  INVX1 U11214 ( .A(n16890), .Y(n5469) );
  INVX1 U11215 ( .A(n18780), .Y(n4915) );
  INVX1 U11216 ( .A(n15000), .Y(n5933) );
  INVX1 U11217 ( .A(n16575), .Y(n5545) );
  INVX1 U11218 ( .A(n18150), .Y(n5115) );
  INVX1 U11219 ( .A(n14685), .Y(n6009) );
  INVX1 U11220 ( .A(n16260), .Y(n5621) );
  INVX1 U11221 ( .A(n17835), .Y(n5223) );
  INVX1 U11222 ( .A(n14370), .Y(n6085) );
  INVX1 U11223 ( .A(n15945), .Y(n5697) );
  INVX1 U11224 ( .A(n17520), .Y(n5301) );
  CLKINVX3 U11225 ( .A(n3986), .Y(n3977) );
  CLKINVX3 U11226 ( .A(n3985), .Y(n3980) );
  CLKINVX3 U11227 ( .A(n3987), .Y(n3979) );
  CLKINVX3 U11228 ( .A(n3986), .Y(n3981) );
  CLKINVX3 U11229 ( .A(n3986), .Y(n3978) );
  CLKINVX3 U11230 ( .A(n3987), .Y(n3982) );
  CLKINVX3 U11231 ( .A(n4092), .Y(n4058) );
  NAND4X1 U11232 ( .A(n17143), .B(n5382), .C(n17144), .D(n17145), .Y(n17142)
         );
  NAND3XL U11233 ( .A(n17126), .B(n17061), .C(top_core_EC_ss_in[82]), .Y(
        n17144) );
  NAND4X1 U11234 ( .A(n13993), .B(n6153), .C(n13994), .D(n13995), .Y(n13992)
         );
  NAND3XL U11235 ( .A(n13976), .B(n13911), .C(top_core_EC_ss_in[2]), .Y(n13994) );
  NAND4X1 U11236 ( .A(n18403), .B(n5028), .C(n18404), .D(n18405), .Y(n18402)
         );
  NAND3XL U11237 ( .A(n18386), .B(n18321), .C(top_core_EC_ss_in[114]), .Y(
        n18404) );
  NAND4X1 U11238 ( .A(n15253), .B(n5854), .C(n15254), .D(n15255), .Y(n15252)
         );
  NAND3XL U11239 ( .A(n15236), .B(n15171), .C(top_core_EC_ss_in[34]), .Y(
        n15254) );
  NAND4X1 U11240 ( .A(n15568), .B(n5770), .C(n15569), .D(n15570), .Y(n15567)
         );
  NAND3XL U11241 ( .A(n15551), .B(n15486), .C(top_core_EC_ss_in[42]), .Y(
        n15569) );
  NAND4X1 U11242 ( .A(n18718), .B(n4912), .C(n18719), .D(n18720), .Y(n18717)
         );
  NAND3XL U11243 ( .A(n18701), .B(n18636), .C(top_core_EC_ss_in[122]), .Y(
        n18719) );
  NAND4X1 U11244 ( .A(n16828), .B(n5466), .C(n16829), .D(n16830), .Y(n16827)
         );
  NAND3XL U11245 ( .A(n16811), .B(n16746), .C(top_core_EC_ss_in[74]), .Y(
        n16829) );
  NAND4X1 U11246 ( .A(n14938), .B(n5930), .C(n14939), .D(n14940), .Y(n14937)
         );
  NAND3XL U11247 ( .A(n14921), .B(n14856), .C(top_core_EC_ss_in[26]), .Y(
        n14939) );
  NAND4X1 U11248 ( .A(n16513), .B(n5542), .C(n16514), .D(n16515), .Y(n16512)
         );
  NAND3XL U11249 ( .A(n16496), .B(n16431), .C(top_core_EC_ss_in[66]), .Y(
        n16514) );
  NAND4X1 U11250 ( .A(n18088), .B(n5112), .C(n18089), .D(n18090), .Y(n18087)
         );
  NAND3XL U11251 ( .A(n18071), .B(n18006), .C(top_core_EC_ss_in[106]), .Y(
        n18089) );
  NAND4X1 U11252 ( .A(n14623), .B(n6006), .C(n14624), .D(n14625), .Y(n14622)
         );
  NAND3XL U11253 ( .A(n14606), .B(n14541), .C(top_core_EC_ss_in[18]), .Y(
        n14624) );
  NAND4X1 U11254 ( .A(n16198), .B(n5618), .C(n16199), .D(n16200), .Y(n16197)
         );
  NAND3XL U11255 ( .A(n16181), .B(n16116), .C(top_core_EC_ss_in[58]), .Y(
        n16199) );
  NAND4X1 U11256 ( .A(n17773), .B(n5220), .C(n17774), .D(n17775), .Y(n17772)
         );
  NAND3XL U11257 ( .A(n17756), .B(n17691), .C(top_core_EC_ss_in[98]), .Y(
        n17774) );
  NAND4X1 U11258 ( .A(n14308), .B(n6082), .C(n14309), .D(n14310), .Y(n14307)
         );
  NAND3XL U11259 ( .A(n14291), .B(n14226), .C(top_core_EC_ss_in[10]), .Y(
        n14309) );
  NAND4X1 U11260 ( .A(n15883), .B(n5694), .C(n15884), .D(n15885), .Y(n15882)
         );
  NAND3XL U11261 ( .A(n15866), .B(n15801), .C(top_core_EC_ss_in[50]), .Y(
        n15884) );
  NAND4X1 U11262 ( .A(n17458), .B(n5298), .C(n17459), .D(n17460), .Y(n17457)
         );
  NAND3XL U11263 ( .A(n17441), .B(n17376), .C(top_core_EC_ss_in[90]), .Y(
        n17459) );
  CLKINVX3 U11264 ( .A(n4115), .Y(n4062) );
  CLKINVX3 U11265 ( .A(n4095), .Y(n4059) );
  CLKINVX3 U11266 ( .A(n4066), .Y(n4064) );
  CLKINVX3 U11267 ( .A(n4066), .Y(n4065) );
  CLKINVX3 U11268 ( .A(n4087), .Y(n4060) );
  CLKINVX3 U11269 ( .A(n4082), .Y(n4061) );
  CLKINVX3 U11270 ( .A(n4083), .Y(n4063) );
  CLKINVX3 U11271 ( .A(n4028), .Y(n4018) );
  OAI21XL U11272 ( .A0(n665), .A1(n11706), .B0(n11772), .Y(n11771) );
  OAI21XL U11273 ( .A0(n666), .A1(top_core_KE_sb1_n131), .B0(
        top_core_KE_sb1_n200), .Y(top_core_KE_sb1_n199) );
  OAI21XL U11274 ( .A0(n670), .A1(n13283), .B0(n13349), .Y(n13348) );
  OAI21XL U11275 ( .A0(n668), .A1(n12022), .B0(n12088), .Y(n12087) );
  OAI21XL U11276 ( .A0(n671), .A1(n12653), .B0(n12719), .Y(n12718) );
  OAI21XL U11277 ( .A0(n669), .A1(n13598), .B0(n13664), .Y(n13663) );
  OAI21XL U11278 ( .A0(n672), .A1(n12968), .B0(n13034), .Y(n13033) );
  AOI21XL U11279 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n76), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n70), .B0(n1145), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n114) );
  AOI21XL U11280 ( .A0(n9893), .A1(n9888), .B0(n1004), .Y(n9929) );
  AOI21XL U11281 ( .A0(n11061), .A1(n11056), .B0(n948), .Y(n11097) );
  AOI21XL U11282 ( .A0(n8141), .A1(n8136), .B0(n1088), .Y(n8177) );
  AOI21XL U11283 ( .A0(n10769), .A1(n10764), .B0(n962), .Y(n10805) );
  AOI21XL U11284 ( .A0(n9017), .A1(n9012), .B0(n1046), .Y(n9053) );
  AOI21XL U11285 ( .A0(n7265), .A1(n7260), .B0(n1130), .Y(n7301) );
  AOI21XL U11286 ( .A0(n10185), .A1(n10180), .B0(n990), .Y(n10221) );
  AOI21XL U11287 ( .A0(n9309), .A1(n9304), .B0(n1032), .Y(n9345) );
  AOI21XL U11288 ( .A0(n8433), .A1(n8428), .B0(n1074), .Y(n8469) );
  AOI21XL U11289 ( .A0(n7557), .A1(n7552), .B0(n1116), .Y(n7593) );
  AOI21XL U11290 ( .A0(n11353), .A1(n11348), .B0(n934), .Y(n11389) );
  AOI21XL U11291 ( .A0(n10477), .A1(n10472), .B0(n976), .Y(n10513) );
  AOI21XL U11292 ( .A0(n9601), .A1(n9596), .B0(n1018), .Y(n9637) );
  AOI21XL U11293 ( .A0(n8725), .A1(n8720), .B0(n1060), .Y(n8761) );
  AOI21XL U11294 ( .A0(n7849), .A1(n7844), .B0(n1102), .Y(n7885) );
  CLKINVX3 U11295 ( .A(n4086), .Y(n4056) );
  CLKINVX3 U11296 ( .A(n4073), .Y(n4053) );
  CLKINVX3 U11297 ( .A(n4074), .Y(n4051) );
  CLKINVX3 U11298 ( .A(n4090), .Y(n4055) );
  CLKINVX3 U11299 ( .A(n3974), .Y(n3970) );
  CLKINVX3 U11300 ( .A(n4114), .Y(n4057) );
  CLKINVX3 U11301 ( .A(n4075), .Y(n4052) );
  CLKINVX3 U11302 ( .A(n4072), .Y(n4050) );
  CLKINVX3 U11303 ( .A(n4092), .Y(n4054) );
  CLKINVX3 U11304 ( .A(n3975), .Y(n3968) );
  CLKINVX3 U11305 ( .A(n3973), .Y(n3965) );
  CLKINVX3 U11306 ( .A(n3974), .Y(n3967) );
  CLKINVX3 U11307 ( .A(n3973), .Y(n3969) );
  CLKINVX3 U11308 ( .A(n3973), .Y(n3966) );
  CLKINVX3 U11309 ( .A(n3974), .Y(n3971) );
  CLKINVX3 U11310 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n131), .Y(n6165) );
  CLKINVX3 U11311 ( .A(n9946), .Y(n5375) );
  CLKINVX3 U11312 ( .A(n11114), .Y(n5021) );
  CLKINVX3 U11313 ( .A(n8194), .Y(n5847) );
  CLKINVX3 U11314 ( .A(n10822), .Y(n5105) );
  CLKINVX3 U11315 ( .A(n9070), .Y(n5611) );
  CLKINVX3 U11316 ( .A(n7318), .Y(n6075) );
  CLKINVX3 U11317 ( .A(n10238), .Y(n5291) );
  CLKINVX3 U11318 ( .A(n9362), .Y(n5535) );
  CLKINVX3 U11319 ( .A(n8486), .Y(n5763) );
  CLKINVX3 U11320 ( .A(n7610), .Y(n5999) );
  CLKINVX3 U11321 ( .A(n11406), .Y(n4905) );
  CLKINVX3 U11322 ( .A(n10530), .Y(n5213) );
  CLKINVX3 U11323 ( .A(n9654), .Y(n5459) );
  CLKINVX3 U11324 ( .A(n8778), .Y(n5687) );
  CLKINVX3 U11325 ( .A(n7902), .Y(n5923) );
  CLKINVX3 U11326 ( .A(n4112), .Y(top_core_EC_n864) );
  AOI21X1 U11327 ( .A0(n5330), .A1(n17298), .B0(n17299), .Y(n17297) );
  OAI32X1 U11328 ( .A0(n2871), .A1(n17300), .A2(n2865), .B0(n1002), .B1(n17031), .Y(n17299) );
  AOI21XL U11329 ( .A0(n17126), .A1(n1311), .B0(n498), .Y(n17300) );
  AOI21X1 U11330 ( .A0(n6114), .A1(n14148), .B0(n14149), .Y(n14147) );
  OAI32X1 U11331 ( .A0(n3473), .A1(n14150), .A2(n3466), .B0(n1141), .B1(n13881), .Y(n14149) );
  AOI21XL U11332 ( .A0(n13976), .A1(n1281), .B0(n497), .Y(n14150) );
  AOI21X1 U11333 ( .A0(n5802), .A1(n15408), .B0(n15409), .Y(n15407) );
  OAI32X1 U11334 ( .A0(n3231), .A1(n15410), .A2(n3225), .B0(n1086), .B1(n15141), .Y(n15409) );
  AOI21XL U11335 ( .A0(n15236), .A1(n1293), .B0(n500), .Y(n15410) );
  AOI21X1 U11336 ( .A0(n4976), .A1(n18558), .B0(n18559), .Y(n18557) );
  OAI32X1 U11337 ( .A0(n2629), .A1(n18560), .A2(n2610), .B0(n946), .B1(n18291), 
        .Y(n18559) );
  AOI21XL U11338 ( .A0(n18386), .A1(n1323), .B0(n501), .Y(n18560) );
  AOI21X1 U11339 ( .A0(n5718), .A1(n15723), .B0(n15724), .Y(n15722) );
  OAI32X1 U11340 ( .A0(n3170), .A1(n15725), .A2(n3164), .B0(n1072), .B1(n15456), .Y(n15724) );
  AOI21XL U11341 ( .A0(n15551), .A1(n1296), .B0(n499), .Y(n15725) );
  AOI21X1 U11342 ( .A0(n5414), .A1(n16983), .B0(n16984), .Y(n16982) );
  OAI32X1 U11343 ( .A0(n2940), .A1(n16985), .A2(n2926), .B0(n1016), .B1(n16716), .Y(n16984) );
  AOI21XL U11344 ( .A0(n16811), .A1(n1308), .B0(n503), .Y(n16985) );
  AOI21X1 U11345 ( .A0(n4860), .A1(n18873), .B0(n18874), .Y(n18872) );
  OAI32X1 U11346 ( .A0(n2568), .A1(n18875), .A2(n2562), .B0(n932), .B1(n18606), 
        .Y(n18874) );
  AOI21XL U11347 ( .A0(n18701), .A1(n1326), .B0(n502), .Y(n18875) );
  AOI21X1 U11348 ( .A0(n5878), .A1(n15093), .B0(n15094), .Y(n15092) );
  OAI32X1 U11349 ( .A0(n3293), .A1(n15095), .A2(n3286), .B0(n1100), .B1(n14826), .Y(n15094) );
  AOI21XL U11350 ( .A0(n14921), .A1(n1290), .B0(n504), .Y(n15095) );
  AOI21X1 U11351 ( .A0(n5490), .A1(n16668), .B0(n16669), .Y(n16667) );
  OAI32X1 U11352 ( .A0(n3001), .A1(n16670), .A2(n2987), .B0(n1030), .B1(n16401), .Y(n16669) );
  AOI21XL U11353 ( .A0(n16496), .A1(n1305), .B0(n505), .Y(n16670) );
  AOI21X1 U11354 ( .A0(n5060), .A1(n18243), .B0(n18244), .Y(n18242) );
  OAI32X1 U11355 ( .A0(n2698), .A1(n18245), .A2(n2684), .B0(n960), .B1(n17976), 
        .Y(n18244) );
  AOI21XL U11356 ( .A0(n18071), .A1(n1320), .B0(n506), .Y(n18245) );
  AOI21X1 U11357 ( .A0(n5954), .A1(n14778), .B0(n14779), .Y(n14777) );
  OAI32X1 U11358 ( .A0(n3353), .A1(n14780), .A2(n3334), .B0(n1114), .B1(n14511), .Y(n14779) );
  AOI21XL U11359 ( .A0(n14606), .A1(n1287), .B0(n507), .Y(n14780) );
  AOI21X1 U11360 ( .A0(n5566), .A1(n16353), .B0(n16354), .Y(n16352) );
  OAI32X1 U11361 ( .A0(n3051), .A1(n16355), .A2(n3032), .B0(n1044), .B1(n16086), .Y(n16354) );
  AOI21XL U11362 ( .A0(n16181), .A1(n1302), .B0(n508), .Y(n16355) );
  AOI21X1 U11363 ( .A0(n5168), .A1(n17928), .B0(n17929), .Y(n17927) );
  OAI32X1 U11364 ( .A0(n2750), .A1(n17930), .A2(n2744), .B0(n974), .B1(n17661), 
        .Y(n17929) );
  AOI21XL U11365 ( .A0(n17756), .A1(n1317), .B0(n509), .Y(n17930) );
  AOI21X1 U11366 ( .A0(n6030), .A1(n14463), .B0(n14464), .Y(n14462) );
  OAI32X1 U11367 ( .A0(n3419), .A1(n14465), .A2(n3392), .B0(n1128), .B1(n14196), .Y(n14464) );
  AOI21XL U11368 ( .A0(n14291), .A1(n1284), .B0(n510), .Y(n14465) );
  AOI21X1 U11369 ( .A0(n5642), .A1(n16038), .B0(n16039), .Y(n16037) );
  OAI32X1 U11370 ( .A0(n3112), .A1(n16040), .A2(n3106), .B0(n1058), .B1(n15771), .Y(n16039) );
  AOI21XL U11371 ( .A0(n15866), .A1(n1299), .B0(n511), .Y(n16040) );
  AOI21X1 U11372 ( .A0(n5246), .A1(n17613), .B0(n17614), .Y(n17612) );
  OAI32X1 U11373 ( .A0(n2812), .A1(n17615), .A2(n2805), .B0(n988), .B1(n17346), 
        .Y(n17614) );
  AOI21XL U11374 ( .A0(n17441), .A1(n1314), .B0(n512), .Y(n17615) );
  OAI2BB2X1 U11375 ( .B0(n1005), .B1(n17162), .A0N(n1310), .A1N(n17167), .Y(
        n17172) );
  OAI2BB2X1 U11376 ( .B0(n1144), .B1(n14012), .A0N(n1280), .A1N(n14017), .Y(
        n14022) );
  OAI2BB2X1 U11377 ( .B0(n949), .B1(n18422), .A0N(n1322), .A1N(n18427), .Y(
        n18432) );
  OAI2BB2X1 U11378 ( .B0(n1089), .B1(n15272), .A0N(n1292), .A1N(n15277), .Y(
        n15282) );
  OAI2BB2X1 U11379 ( .B0(n1075), .B1(n15587), .A0N(n1295), .A1N(n15592), .Y(
        n15597) );
  OAI2BB2X1 U11380 ( .B0(n935), .B1(n18737), .A0N(n1325), .A1N(n18742), .Y(
        n18747) );
  OAI2BB2X1 U11381 ( .B0(n1019), .B1(n16847), .A0N(n1307), .A1N(n16852), .Y(
        n16857) );
  OAI2BB2X1 U11382 ( .B0(n1103), .B1(n14957), .A0N(n1289), .A1N(n14962), .Y(
        n14967) );
  OAI2BB2X1 U11383 ( .B0(n1033), .B1(n16532), .A0N(n1304), .A1N(n16537), .Y(
        n16542) );
  OAI2BB2X1 U11384 ( .B0(n963), .B1(n18107), .A0N(n1319), .A1N(n18112), .Y(
        n18117) );
  OAI2BB2X1 U11385 ( .B0(n1117), .B1(n14642), .A0N(n1286), .A1N(n14647), .Y(
        n14652) );
  OAI2BB2X1 U11386 ( .B0(n1047), .B1(n16217), .A0N(n1301), .A1N(n16222), .Y(
        n16227) );
  OAI2BB2X1 U11387 ( .B0(n977), .B1(n17792), .A0N(n1316), .A1N(n17797), .Y(
        n17802) );
  OAI2BB2X1 U11388 ( .B0(n1131), .B1(n14327), .A0N(n1283), .A1N(n14332), .Y(
        n14337) );
  OAI2BB2X1 U11389 ( .B0(n1061), .B1(n15902), .A0N(n1298), .A1N(n15907), .Y(
        n15912) );
  OAI2BB2X1 U11390 ( .B0(n991), .B1(n17477), .A0N(n1313), .A1N(n17482), .Y(
        n17487) );
  AOI2BB1X1 U11391 ( .A0N(n999), .A1N(n17060), .B0(n1005), .Y(n17152) );
  AOI2BB1X1 U11392 ( .A0N(n1138), .A1N(n13910), .B0(n1144), .Y(n14002) );
  AOI2BB1X1 U11393 ( .A0N(n943), .A1N(n18320), .B0(n949), .Y(n18412) );
  AOI2BB1X1 U11394 ( .A0N(n1083), .A1N(n15170), .B0(n1089), .Y(n15262) );
  AOI2BB1X1 U11395 ( .A0N(n1069), .A1N(n15485), .B0(n1075), .Y(n15577) );
  AOI2BB1X1 U11396 ( .A0N(n929), .A1N(n18635), .B0(n935), .Y(n18727) );
  AOI2BB1X1 U11397 ( .A0N(n1013), .A1N(n16745), .B0(n1019), .Y(n16837) );
  AOI2BB1X1 U11398 ( .A0N(n1097), .A1N(n14855), .B0(n1103), .Y(n14947) );
  AOI2BB1X1 U11399 ( .A0N(n1027), .A1N(n16430), .B0(n1033), .Y(n16522) );
  AOI2BB1X1 U11400 ( .A0N(n957), .A1N(n18005), .B0(n963), .Y(n18097) );
  AOI2BB1X1 U11401 ( .A0N(n1111), .A1N(n14540), .B0(n1117), .Y(n14632) );
  AOI2BB1X1 U11402 ( .A0N(n1041), .A1N(n16115), .B0(n1047), .Y(n16207) );
  AOI2BB1X1 U11403 ( .A0N(n971), .A1N(n17690), .B0(n977), .Y(n17782) );
  AOI2BB1X1 U11404 ( .A0N(n1125), .A1N(n14225), .B0(n1131), .Y(n14317) );
  AOI2BB1X1 U11405 ( .A0N(n1055), .A1N(n15800), .B0(n1061), .Y(n15892) );
  AOI2BB1X1 U11406 ( .A0N(n985), .A1N(n17375), .B0(n991), .Y(n17467) );
  NAND4X1 U11407 ( .A(n17163), .B(n17164), .C(n17165), .D(n17166), .Y(n17158)
         );
  NAND4X1 U11408 ( .A(n14013), .B(n14014), .C(n14015), .D(n14016), .Y(n14008)
         );
  NAND4X1 U11409 ( .A(n18423), .B(n18424), .C(n18425), .D(n18426), .Y(n18418)
         );
  NAND4X1 U11410 ( .A(n15273), .B(n15274), .C(n15275), .D(n15276), .Y(n15268)
         );
  NAND4X1 U11411 ( .A(n15588), .B(n15589), .C(n15590), .D(n15591), .Y(n15583)
         );
  NAND4X1 U11412 ( .A(n18738), .B(n18739), .C(n18740), .D(n18741), .Y(n18733)
         );
  NAND4X1 U11413 ( .A(n16848), .B(n16849), .C(n16850), .D(n16851), .Y(n16843)
         );
  NAND4X1 U11414 ( .A(n14958), .B(n14959), .C(n14960), .D(n14961), .Y(n14953)
         );
  NAND4X1 U11415 ( .A(n16533), .B(n16534), .C(n16535), .D(n16536), .Y(n16528)
         );
  NAND4X1 U11416 ( .A(n18108), .B(n18109), .C(n18110), .D(n18111), .Y(n18103)
         );
  NAND4X1 U11417 ( .A(n14643), .B(n14644), .C(n14645), .D(n14646), .Y(n14638)
         );
  NAND4X1 U11418 ( .A(n16218), .B(n16219), .C(n16220), .D(n16221), .Y(n16213)
         );
  NAND4X1 U11419 ( .A(n17793), .B(n17794), .C(n17795), .D(n17796), .Y(n17788)
         );
  NAND4X1 U11420 ( .A(n14328), .B(n14329), .C(n14330), .D(n14331), .Y(n14323)
         );
  NAND4X1 U11421 ( .A(n15903), .B(n15904), .C(n15905), .D(n15906), .Y(n15898)
         );
  NAND4X1 U11422 ( .A(n17478), .B(n17479), .C(n17480), .D(n17481), .Y(n17473)
         );
  NAND4BXL U11423 ( .AN(n13438), .B(n13439), .C(n13384), .D(n13363), .Y(n13437) );
  AOI21XL U11424 ( .A0(n13282), .A1(n6556), .B0(n13318), .Y(n13439) );
  CLKINVX3 U11425 ( .A(n11806), .Y(n6919) );
  CLKINVX3 U11426 ( .A(top_core_KE_sb1_n234), .Y(n6873) );
  CLKINVX3 U11427 ( .A(n13382), .Y(n6554) );
  CLKINVX3 U11428 ( .A(n12122), .Y(n6579) );
  CLKINVX3 U11429 ( .A(n12752), .Y(n6849) );
  CLKINVX3 U11430 ( .A(n13067), .Y(n6895) );
  CLKINVX3 U11431 ( .A(n13697), .Y(n6602) );
  AOI2BB2X1 U11432 ( .B0(n13860), .B1(n1138), .A0N(n13861), .A1N(n385), .Y(
        n13850) );
  AOI21X1 U11433 ( .A0(n3467), .A1(n6114), .B0(n13862), .Y(n13861) );
  AOI2BB2X1 U11434 ( .B0(n17010), .B1(n999), .A0N(n17011), .A1N(n386), .Y(
        n17000) );
  AOI21X1 U11435 ( .A0(n2866), .A1(n5330), .B0(n17012), .Y(n17011) );
  AOI2BB2X1 U11436 ( .B0(n18270), .B1(n943), .A0N(n18271), .A1N(n387), .Y(
        n18260) );
  AOI21X1 U11437 ( .A0(n2624), .A1(n4976), .B0(n18272), .Y(n18271) );
  AOI2BB2X1 U11438 ( .B0(n15120), .B1(n1083), .A0N(n15121), .A1N(n388), .Y(
        n15110) );
  AOI21X1 U11439 ( .A0(n3226), .A1(n5802), .B0(n15122), .Y(n15121) );
  AOI2BB2X1 U11440 ( .B0(n15435), .B1(n1069), .A0N(n15436), .A1N(n389), .Y(
        n15425) );
  AOI21X1 U11441 ( .A0(n3165), .A1(n5718), .B0(n15437), .Y(n15436) );
  AOI2BB2X1 U11442 ( .B0(n18585), .B1(n929), .A0N(n18586), .A1N(n390), .Y(
        n18575) );
  AOI21X1 U11443 ( .A0(n2563), .A1(n4860), .B0(n18587), .Y(n18586) );
  AOI2BB2X1 U11444 ( .B0(n16695), .B1(n1013), .A0N(n16696), .A1N(n391), .Y(
        n16685) );
  AOI21X1 U11445 ( .A0(n2927), .A1(n5414), .B0(n16697), .Y(n16696) );
  AOI2BB2X1 U11446 ( .B0(n14805), .B1(n1097), .A0N(n14806), .A1N(n392), .Y(
        n14795) );
  AOI21X1 U11447 ( .A0(n3287), .A1(n5878), .B0(n14807), .Y(n14806) );
  AOI2BB2X1 U11448 ( .B0(n16380), .B1(n1027), .A0N(n16381), .A1N(n393), .Y(
        n16370) );
  AOI21X1 U11449 ( .A0(n2988), .A1(n5490), .B0(n16382), .Y(n16381) );
  AOI2BB2X1 U11450 ( .B0(n17955), .B1(n957), .A0N(n17956), .A1N(n394), .Y(
        n17945) );
  AOI21X1 U11451 ( .A0(n2685), .A1(n5060), .B0(n17957), .Y(n17956) );
  AOI2BB2X1 U11452 ( .B0(n14490), .B1(n1111), .A0N(n14491), .A1N(n395), .Y(
        n14480) );
  AOI21X1 U11453 ( .A0(n3348), .A1(n5954), .B0(n14492), .Y(n14491) );
  AOI2BB2X1 U11454 ( .B0(n16065), .B1(n1041), .A0N(n16066), .A1N(n396), .Y(
        n16055) );
  AOI21X1 U11455 ( .A0(n3046), .A1(n5566), .B0(n16067), .Y(n16066) );
  AOI2BB2X1 U11456 ( .B0(n17640), .B1(n971), .A0N(n17641), .A1N(n397), .Y(
        n17630) );
  AOI21X1 U11457 ( .A0(n2745), .A1(n5168), .B0(n17642), .Y(n17641) );
  AOI2BB2X1 U11458 ( .B0(n14175), .B1(n1125), .A0N(n14176), .A1N(n398), .Y(
        n14165) );
  AOI21X1 U11459 ( .A0(n3406), .A1(n6030), .B0(n14177), .Y(n14176) );
  AOI2BB2X1 U11460 ( .B0(n15750), .B1(n1055), .A0N(n15751), .A1N(n399), .Y(
        n15740) );
  AOI21X1 U11461 ( .A0(n3107), .A1(n5642), .B0(n15752), .Y(n15751) );
  AOI2BB2X1 U11462 ( .B0(n17325), .B1(n985), .A0N(n17326), .A1N(n400), .Y(
        n17315) );
  AOI21X1 U11463 ( .A0(n2806), .A1(n5246), .B0(n17327), .Y(n17326) );
  NAND4BXL U11464 ( .AN(n13393), .B(n13225), .C(n13375), .D(n13384), .Y(n13391) );
  NAND4BXL U11465 ( .AN(n12763), .B(n12595), .C(n12745), .D(n12754), .Y(n12761) );
  NAND4BXL U11466 ( .AN(n13708), .B(n13540), .C(n13690), .D(n13699), .Y(n13706) );
  NAND4BXL U11467 ( .AN(n13078), .B(n12910), .C(n13060), .D(n13069), .Y(n13076) );
  NAND3XL U11468 ( .A(n1732), .B(n1269), .C(n719), .Y(n12755) );
  NAND3XL U11469 ( .A(n1703), .B(n1272), .C(n721), .Y(n13070) );
  AOI21XL U11470 ( .A0(n180), .A1(n13250), .B0(n1666), .Y(n13405) );
  AOI21XL U11471 ( .A0(n181), .A1(n12620), .B0(n1724), .Y(n12775) );
  AOI21XL U11472 ( .A0(n182), .A1(n12935), .B0(n1695), .Y(n13090) );
  CLKINVX3 U11473 ( .A(n3450), .Y(n3447) );
  CLKINVX3 U11474 ( .A(n2849), .Y(n2846) );
  CLKINVX3 U11475 ( .A(n2607), .Y(n2604) );
  CLKINVX3 U11476 ( .A(n3209), .Y(n3206) );
  CLKINVX3 U11477 ( .A(n2668), .Y(n2665) );
  CLKINVX3 U11478 ( .A(n3029), .Y(n3026) );
  CLKINVX3 U11479 ( .A(n3389), .Y(n3386) );
  CLKINVX3 U11480 ( .A(n2971), .Y(n2968) );
  CLKINVX3 U11481 ( .A(n3148), .Y(n3145) );
  CLKINVX3 U11482 ( .A(n3331), .Y(n3328) );
  CLKINVX3 U11483 ( .A(n2546), .Y(n2543) );
  CLKINVX3 U11484 ( .A(n2728), .Y(n2725) );
  CLKINVX3 U11485 ( .A(n2910), .Y(n2907) );
  CLKINVX3 U11486 ( .A(n3090), .Y(n3087) );
  CLKINVX3 U11487 ( .A(n2789), .Y(n2786) );
  CLKINVX3 U11488 ( .A(n3270), .Y(n3267) );
  CLKINVX3 U11489 ( .A(n1894), .Y(n1889) );
  CLKINVX3 U11490 ( .A(n1934), .Y(n1929) );
  CLKINVX3 U11491 ( .A(n1974), .Y(n1968) );
  CLKINVX3 U11492 ( .A(n2094), .Y(n2088) );
  CLKINVX3 U11493 ( .A(n2134), .Y(n2128) );
  CLKINVX3 U11494 ( .A(n1895), .Y(n1886) );
  CLKINVX3 U11495 ( .A(n1935), .Y(n1926) );
  CLKINVX3 U11496 ( .A(n1975), .Y(n1966) );
  CLKINVX3 U11497 ( .A(n2055), .Y(n2046) );
  CLKINVX3 U11498 ( .A(n2095), .Y(n2085) );
  CLKINVX3 U11499 ( .A(n2135), .Y(n2125) );
  CLKINVX3 U11500 ( .A(n1894), .Y(n1887) );
  CLKINVX3 U11501 ( .A(n1934), .Y(n1927) );
  CLKINVX3 U11502 ( .A(n1974), .Y(n1967) );
  CLKINVX3 U11503 ( .A(n2054), .Y(n2047) );
  CLKINVX3 U11504 ( .A(n2094), .Y(n2086) );
  CLKINVX3 U11505 ( .A(n2134), .Y(n2126) );
  CLKINVX3 U11506 ( .A(n1894), .Y(n1890) );
  CLKINVX3 U11507 ( .A(n1974), .Y(n1969) );
  CLKINVX3 U11508 ( .A(n2054), .Y(n2049) );
  CLKINVX3 U11509 ( .A(n2094), .Y(n2089) );
  CLKINVX3 U11510 ( .A(n2134), .Y(n2129) );
  CLKINVX3 U11511 ( .A(n1893), .Y(n1891) );
  CLKINVX3 U11512 ( .A(n1933), .Y(n1930) );
  CLKINVX3 U11513 ( .A(n1973), .Y(n1970) );
  CLKINVX3 U11514 ( .A(n2053), .Y(n2050) );
  CLKINVX3 U11515 ( .A(n2093), .Y(n2090) );
  CLKINVX3 U11516 ( .A(n2133), .Y(n2130) );
  CLKINVX3 U11517 ( .A(n1893), .Y(n1892) );
  CLKINVX3 U11518 ( .A(n1933), .Y(n1931) );
  CLKINVX3 U11519 ( .A(n1973), .Y(n1971) );
  CLKINVX3 U11520 ( .A(n2053), .Y(n2051) );
  CLKINVX3 U11521 ( .A(n2093), .Y(n2091) );
  CLKINVX3 U11522 ( .A(n2133), .Y(n2131) );
  CLKINVX3 U11523 ( .A(n1934), .Y(n1932) );
  CLKINVX3 U11524 ( .A(n1974), .Y(n1972) );
  CLKINVX3 U11525 ( .A(n2054), .Y(n2052) );
  CLKINVX3 U11526 ( .A(n2094), .Y(n2092) );
  CLKINVX3 U11527 ( .A(n2134), .Y(n2132) );
  CLKINVX3 U11528 ( .A(n1894), .Y(n1888) );
  CLKINVX3 U11529 ( .A(n1934), .Y(n1928) );
  CLKINVX3 U11530 ( .A(n2054), .Y(n2048) );
  CLKINVX3 U11531 ( .A(n2094), .Y(n2087) );
  CLKINVX3 U11532 ( .A(n2134), .Y(n2127) );
  CLKINVX3 U11533 ( .A(n2015), .Y(n2005) );
  CLKINVX3 U11534 ( .A(n2014), .Y(n2006) );
  CLKINVX3 U11535 ( .A(n2014), .Y(n2008) );
  CLKINVX3 U11536 ( .A(n2014), .Y(n2009) );
  CLKINVX3 U11537 ( .A(n2013), .Y(n2010) );
  CLKINVX3 U11538 ( .A(n2013), .Y(n2011) );
  CLKINVX3 U11539 ( .A(n2014), .Y(n2012) );
  CLKINVX3 U11540 ( .A(n2014), .Y(n2007) );
  CLKINVX3 U11541 ( .A(n1608), .Y(n1603) );
  CLKINVX3 U11542 ( .A(n1607), .Y(n1602) );
  CLKINVX3 U11543 ( .A(n1608), .Y(n1601) );
  CLKINVX3 U11544 ( .A(n1605), .Y(n1600) );
  CLKINVX3 U11545 ( .A(n1605), .Y(n1599) );
  CLKINVX3 U11546 ( .A(n1606), .Y(n1598) );
  CLKINVX3 U11547 ( .A(n1605), .Y(n1597) );
  CLKINVX3 U11548 ( .A(n1605), .Y(n1596) );
  CLKINVX3 U11549 ( .A(n1606), .Y(n1595) );
  CLKINVX3 U11550 ( .A(n1606), .Y(n1594) );
  CLKINVX3 U11551 ( .A(top_core_io_inter_ok), .Y(n1593) );
  CLKINVX3 U11552 ( .A(top_core_io_inter_ok), .Y(n1592) );
  CLKINVX3 U11553 ( .A(n1607), .Y(n1591) );
  CLKINVX3 U11554 ( .A(n1607), .Y(n1590) );
  CLKINVX3 U11555 ( .A(n1605), .Y(n1589) );
  CLKINVX3 U11556 ( .A(n1607), .Y(n1588) );
  CLKINVX3 U11557 ( .A(n1606), .Y(n1587) );
  CLKINVX3 U11558 ( .A(top_core_io_inter_ok), .Y(n1586) );
  CLKINVX3 U11559 ( .A(n1608), .Y(n1585) );
  CLKINVX3 U11560 ( .A(n1608), .Y(n1584) );
  CLKINVX3 U11561 ( .A(n1893), .Y(n1885) );
  CLKINVX3 U11562 ( .A(n1933), .Y(n1925) );
  CLKINVX3 U11563 ( .A(n1973), .Y(n1965) );
  CLKINVX3 U11564 ( .A(n2053), .Y(n2045) );
  CLKINVX3 U11565 ( .A(n2093), .Y(n2084) );
  CLKINVX3 U11566 ( .A(n2133), .Y(n2124) );
  CLKINVX3 U11567 ( .A(n2013), .Y(n2004) );
  CLKINVX3 U11568 ( .A(n3573), .Y(n3570) );
  CLKINVX3 U11569 ( .A(n3573), .Y(n3571) );
  CLKINVX3 U11570 ( .A(n3907), .Y(n3906) );
  CLKINVX3 U11571 ( .A(n11852), .Y(n6904) );
  CLKINVX3 U11572 ( .A(top_core_KE_sb1_n281), .Y(n6858) );
  CLKINVX3 U11573 ( .A(n13428), .Y(n6539) );
  CLKINVX3 U11574 ( .A(n12168), .Y(n6564) );
  CLKINVX3 U11575 ( .A(n12798), .Y(n6834) );
  CLKINVX3 U11576 ( .A(n13743), .Y(n6587) );
  CLKINVX3 U11577 ( .A(n13113), .Y(n6880) );
  CLKINVX3 U11578 ( .A(n1896), .Y(n1878) );
  CLKINVX3 U11579 ( .A(n1936), .Y(n1918) );
  CLKINVX3 U11580 ( .A(n1976), .Y(n1958) );
  CLKINVX3 U11581 ( .A(n2056), .Y(n2038) );
  CLKINVX3 U11582 ( .A(n2136), .Y(n2117) );
  CLKINVX3 U11583 ( .A(n1896), .Y(n1877) );
  CLKINVX3 U11584 ( .A(n1936), .Y(n1917) );
  CLKINVX3 U11585 ( .A(n1976), .Y(n1957) );
  CLKINVX3 U11586 ( .A(n2056), .Y(n2037) );
  CLKINVX3 U11587 ( .A(n2096), .Y(n2077) );
  CLKINVX3 U11588 ( .A(n1896), .Y(n1879) );
  CLKINVX3 U11589 ( .A(n1936), .Y(n1919) );
  CLKINVX3 U11590 ( .A(n1976), .Y(n1959) );
  CLKINVX3 U11591 ( .A(n2056), .Y(n2039) );
  CLKINVX3 U11592 ( .A(n2096), .Y(n2078) );
  CLKINVX3 U11593 ( .A(n2136), .Y(n2118) );
  CLKINVX3 U11594 ( .A(n1896), .Y(n1880) );
  CLKINVX3 U11595 ( .A(n1936), .Y(n1920) );
  CLKINVX3 U11596 ( .A(n1976), .Y(n1960) );
  CLKINVX3 U11597 ( .A(n2056), .Y(n2040) );
  CLKINVX3 U11598 ( .A(n2096), .Y(n2079) );
  CLKINVX3 U11599 ( .A(n2136), .Y(n2119) );
  CLKINVX3 U11600 ( .A(n1896), .Y(n1881) );
  CLKINVX3 U11601 ( .A(n1936), .Y(n1921) );
  CLKINVX3 U11602 ( .A(n1976), .Y(n1961) );
  CLKINVX3 U11603 ( .A(n2056), .Y(n2041) );
  CLKINVX3 U11604 ( .A(n2096), .Y(n2080) );
  CLKINVX3 U11605 ( .A(n2136), .Y(n2120) );
  CLKINVX3 U11606 ( .A(n1895), .Y(n1882) );
  CLKINVX3 U11607 ( .A(n1935), .Y(n1922) );
  CLKINVX3 U11608 ( .A(n1975), .Y(n1962) );
  CLKINVX3 U11609 ( .A(n2055), .Y(n2042) );
  CLKINVX3 U11610 ( .A(n2095), .Y(n2081) );
  CLKINVX3 U11611 ( .A(n2135), .Y(n2121) );
  CLKINVX3 U11612 ( .A(n1895), .Y(n1883) );
  CLKINVX3 U11613 ( .A(n1935), .Y(n1923) );
  CLKINVX3 U11614 ( .A(n1975), .Y(n1963) );
  CLKINVX3 U11615 ( .A(n2055), .Y(n2043) );
  CLKINVX3 U11616 ( .A(n2095), .Y(n2082) );
  CLKINVX3 U11617 ( .A(n2135), .Y(n2122) );
  CLKINVX3 U11618 ( .A(n1895), .Y(n1884) );
  CLKINVX3 U11619 ( .A(n1935), .Y(n1924) );
  CLKINVX3 U11620 ( .A(n1975), .Y(n1964) );
  CLKINVX3 U11621 ( .A(n2055), .Y(n2044) );
  CLKINVX3 U11622 ( .A(n2095), .Y(n2083) );
  CLKINVX3 U11623 ( .A(n2135), .Y(n2123) );
  CLKINVX3 U11624 ( .A(n2016), .Y(n1997) );
  CLKINVX3 U11625 ( .A(n2016), .Y(n1998) );
  CLKINVX3 U11626 ( .A(n2016), .Y(n1999) );
  CLKINVX3 U11627 ( .A(n2016), .Y(n2000) );
  CLKINVX3 U11628 ( .A(n2015), .Y(n2001) );
  CLKINVX3 U11629 ( .A(n2015), .Y(n2002) );
  CLKINVX3 U11630 ( .A(n2015), .Y(n2003) );
  CLKINVX3 U11631 ( .A(n741), .Y(n2312) );
  CLKINVX3 U11632 ( .A(n2316), .Y(n2313) );
  CLKINVX3 U11633 ( .A(n742), .Y(n3560) );
  CLKINVX3 U11634 ( .A(n742), .Y(n3559) );
  CLKINVX3 U11635 ( .A(n3543), .Y(n3534) );
  INVX1 U11636 ( .A(top_core_EC_n733), .Y(n3543) );
  CLKINVX3 U11637 ( .A(n2326), .Y(n2317) );
  INVX1 U11638 ( .A(n11883), .Y(n6829) );
  INVX1 U11639 ( .A(top_core_KE_sb1_n312), .Y(n6808) );
  INVX1 U11640 ( .A(n12514), .Y(n6533) );
  INVX1 U11641 ( .A(n12199), .Y(n6511) );
  INVX1 U11642 ( .A(n13459), .Y(n6476) );
  INVX1 U11643 ( .A(n12829), .Y(n6779) );
  INVX1 U11644 ( .A(n13774), .Y(n6522) );
  INVX1 U11645 ( .A(n13144), .Y(n6818) );
  NAND3XL U11646 ( .A(n2881), .B(n17126), .C(n5330), .Y(n17181) );
  NAND3XL U11647 ( .A(n3482), .B(n13976), .C(n6114), .Y(n14031) );
  NAND3XL U11648 ( .A(n2639), .B(n18386), .C(n4976), .Y(n18441) );
  NAND3XL U11649 ( .A(n3241), .B(n15236), .C(n5802), .Y(n15291) );
  NAND3XL U11650 ( .A(n3180), .B(n15551), .C(n5718), .Y(n15606) );
  NAND3XL U11651 ( .A(n2942), .B(n16811), .C(n5414), .Y(n16866) );
  NAND3XL U11652 ( .A(n2578), .B(n18701), .C(n4860), .Y(n18756) );
  NAND3XL U11653 ( .A(n3302), .B(n14921), .C(n5878), .Y(n14976) );
  NAND3XL U11654 ( .A(n3003), .B(n16496), .C(n5490), .Y(n16551) );
  NAND3XL U11655 ( .A(n2700), .B(n18071), .C(n5060), .Y(n18126) );
  NAND3XL U11656 ( .A(n3363), .B(n14606), .C(n5954), .Y(n14661) );
  NAND3XL U11657 ( .A(n3061), .B(n16181), .C(n5566), .Y(n16236) );
  NAND3XL U11658 ( .A(n2760), .B(n17756), .C(n5168), .Y(n17811) );
  NAND3XL U11659 ( .A(n3421), .B(n14291), .C(n6030), .Y(n14346) );
  NAND3XL U11660 ( .A(n3122), .B(n15866), .C(n5642), .Y(n15921) );
  NAND3XL U11661 ( .A(n2821), .B(n17441), .C(n5246), .Y(n17496) );
  NAND4X1 U11662 ( .A(n13963), .B(n13875), .C(n14112), .D(n14113), .Y(n14111)
         );
  AOI222X1 U11663 ( .A0(n1134), .A1(n1142), .B0(n6149), .B1(n497), .C0(n369), 
        .C1(n1136), .Y(n14113) );
  NAND4X1 U11664 ( .A(n17113), .B(n17025), .C(n17262), .D(n17263), .Y(n17261)
         );
  AOI222X1 U11665 ( .A0(n995), .A1(n1003), .B0(n5378), .B1(n498), .C0(n370), 
        .C1(n997), .Y(n17263) );
  NAND4X1 U11666 ( .A(n18373), .B(n18285), .C(n18522), .D(n18523), .Y(n18521)
         );
  AOI222X1 U11667 ( .A0(n939), .A1(n947), .B0(n5024), .B1(n501), .C0(n371), 
        .C1(n941), .Y(n18523) );
  NAND4X1 U11668 ( .A(n15223), .B(n15135), .C(n15372), .D(n15373), .Y(n15371)
         );
  AOI222X1 U11669 ( .A0(n1079), .A1(n1087), .B0(n5850), .B1(n500), .C0(n372), 
        .C1(n1081), .Y(n15373) );
  NAND4X1 U11670 ( .A(n15538), .B(n15450), .C(n15687), .D(n15688), .Y(n15686)
         );
  AOI222X1 U11671 ( .A0(n1065), .A1(n1073), .B0(n5766), .B1(n499), .C0(n373), 
        .C1(n1067), .Y(n15688) );
  NAND4X1 U11672 ( .A(n18688), .B(n18600), .C(n18837), .D(n18838), .Y(n18836)
         );
  AOI222X1 U11673 ( .A0(n925), .A1(n933), .B0(n4908), .B1(n502), .C0(n374), 
        .C1(n927), .Y(n18838) );
  NAND4X1 U11674 ( .A(n16798), .B(n16710), .C(n16947), .D(n16948), .Y(n16946)
         );
  AOI222X1 U11675 ( .A0(n1009), .A1(n1017), .B0(n5462), .B1(n503), .C0(n375), 
        .C1(n1011), .Y(n16948) );
  NAND4X1 U11676 ( .A(n14908), .B(n14820), .C(n15057), .D(n15058), .Y(n15056)
         );
  AOI222X1 U11677 ( .A0(n1093), .A1(n1101), .B0(n5926), .B1(n504), .C0(n376), 
        .C1(n1095), .Y(n15058) );
  NAND4X1 U11678 ( .A(n16483), .B(n16395), .C(n16632), .D(n16633), .Y(n16631)
         );
  AOI222X1 U11679 ( .A0(n1023), .A1(n1031), .B0(n5538), .B1(n505), .C0(n377), 
        .C1(n1025), .Y(n16633) );
  NAND4X1 U11680 ( .A(n18058), .B(n17970), .C(n18207), .D(n18208), .Y(n18206)
         );
  AOI222X1 U11681 ( .A0(n953), .A1(n961), .B0(n5108), .B1(n506), .C0(n378), 
        .C1(n955), .Y(n18208) );
  NAND4X1 U11682 ( .A(n14593), .B(n14505), .C(n14742), .D(n14743), .Y(n14741)
         );
  AOI222X1 U11683 ( .A0(n1107), .A1(n1115), .B0(n6002), .B1(n507), .C0(n379), 
        .C1(n1109), .Y(n14743) );
  NAND4X1 U11684 ( .A(n16168), .B(n16080), .C(n16317), .D(n16318), .Y(n16316)
         );
  AOI222X1 U11685 ( .A0(n1037), .A1(n1045), .B0(n5614), .B1(n508), .C0(n380), 
        .C1(n1039), .Y(n16318) );
  NAND4X1 U11686 ( .A(n17743), .B(n17655), .C(n17892), .D(n17893), .Y(n17891)
         );
  AOI222X1 U11687 ( .A0(n967), .A1(n975), .B0(n5216), .B1(n509), .C0(n381), 
        .C1(n969), .Y(n17893) );
  NAND4X1 U11688 ( .A(n14278), .B(n14190), .C(n14427), .D(n14428), .Y(n14426)
         );
  AOI222X1 U11689 ( .A0(n1121), .A1(n1129), .B0(n6078), .B1(n510), .C0(n382), 
        .C1(n1123), .Y(n14428) );
  NAND4X1 U11690 ( .A(n15853), .B(n15765), .C(n16002), .D(n16003), .Y(n16001)
         );
  AOI222X1 U11691 ( .A0(n1051), .A1(n1059), .B0(n5690), .B1(n511), .C0(n383), 
        .C1(n1053), .Y(n16003) );
  NAND4X1 U11692 ( .A(n17428), .B(n17340), .C(n17577), .D(n17578), .Y(n17576)
         );
  AOI222X1 U11693 ( .A0(n981), .A1(n989), .B0(n5294), .B1(n512), .C0(n384), 
        .C1(n983), .Y(n17578) );
  NAND4BXL U11694 ( .AN(n13219), .B(n13375), .C(n13484), .D(n13485), .Y(n13480) );
  AOI222X1 U11695 ( .A0(n677), .A1(n1151), .B0(n6556), .B1(n1173), .C0(n1148), 
        .C1(n670), .Y(n13485) );
  AOI2BB2X1 U11696 ( .B0(n6554), .B1(n1687), .A0N(n13443), .A1N(n677), .Y(
        n13484) );
  NAND4BXL U11697 ( .AN(n12589), .B(n12745), .C(n12854), .D(n12855), .Y(n12850) );
  AOI222X1 U11698 ( .A0(n678), .A1(n1191), .B0(n6851), .B1(n1213), .C0(n1188), 
        .C1(n688), .Y(n12855) );
  AOI2BB2X1 U11699 ( .B0(n6849), .B1(n1745), .A0N(n12813), .A1N(n678), .Y(
        n12854) );
  NAND4BXL U11700 ( .AN(n13534), .B(n13690), .C(n13799), .D(n13800), .Y(n13795) );
  AOI222X1 U11701 ( .A0(n679), .A1(n1160), .B0(n6604), .B1(n1178), .C0(n1157), 
        .C1(n685), .Y(n13800) );
  AOI2BB2X1 U11702 ( .B0(n6602), .B1(n1658), .A0N(n13758), .A1N(n679), .Y(
        n13799) );
  NAND4BXL U11703 ( .AN(n12904), .B(n13060), .C(n13169), .D(n13170), .Y(n13165) );
  AOI222X1 U11704 ( .A0(n680), .A1(n1200), .B0(n6897), .B1(n1219), .C0(n1197), 
        .C1(n687), .Y(n13170) );
  AOI2BB2X1 U11705 ( .B0(n6895), .B1(n1716), .A0N(n13128), .A1N(n680), .Y(
        n13169) );
  NAND4X1 U11706 ( .A(n14116), .B(n14117), .C(n14118), .D(n14119), .Y(n14109)
         );
  AOI2BB2X1 U11707 ( .B0(n3457), .B1(n14120), .A0N(n13881), .A1N(n497), .Y(
        n14118) );
  AOI2BB2X1 U11708 ( .B0(n6114), .B1(n14004), .A0N(n107), .A1N(n13868), .Y(
        n14116) );
  NAND4X1 U11709 ( .A(n17266), .B(n17267), .C(n17268), .D(n17269), .Y(n17259)
         );
  AOI2BB2X1 U11710 ( .B0(n2856), .B1(n17270), .A0N(n17031), .A1N(n498), .Y(
        n17268) );
  AOI2BB2X1 U11711 ( .B0(n5330), .B1(n17154), .A0N(n106), .A1N(n17018), .Y(
        n17266) );
  NAND4X1 U11712 ( .A(n18526), .B(n18527), .C(n18528), .D(n18529), .Y(n18519)
         );
  AOI2BB2X1 U11713 ( .B0(n2616), .B1(n18530), .A0N(n18291), .A1N(n501), .Y(
        n18528) );
  AOI2BB2X1 U11714 ( .B0(n4976), .B1(n18414), .A0N(n108), .A1N(n18278), .Y(
        n18526) );
  NAND4X1 U11715 ( .A(n15376), .B(n15377), .C(n15378), .D(n15379), .Y(n15369)
         );
  AOI2BB2X1 U11716 ( .B0(n3216), .B1(n15380), .A0N(n15141), .A1N(n500), .Y(
        n15378) );
  AOI2BB2X1 U11717 ( .B0(n5802), .B1(n15264), .A0N(n109), .A1N(n15128), .Y(
        n15376) );
  NAND4X1 U11718 ( .A(n15691), .B(n15692), .C(n15693), .D(n15694), .Y(n15684)
         );
  AOI2BB2X1 U11719 ( .B0(n3157), .B1(n15695), .A0N(n15456), .A1N(n499), .Y(
        n15693) );
  AOI2BB2X1 U11720 ( .B0(n5718), .B1(n15579), .A0N(n110), .A1N(n15443), .Y(
        n15691) );
  NAND4X1 U11721 ( .A(n18841), .B(n18842), .C(n18843), .D(n18844), .Y(n18834)
         );
  AOI2BB2X1 U11722 ( .B0(n2553), .B1(n18845), .A0N(n18606), .A1N(n502), .Y(
        n18843) );
  AOI2BB2X1 U11723 ( .B0(n4860), .B1(n18729), .A0N(n111), .A1N(n18593), .Y(
        n18841) );
  NAND4X1 U11724 ( .A(n16951), .B(n16952), .C(n16953), .D(n16954), .Y(n16944)
         );
  AOI2BB2X1 U11725 ( .B0(n2919), .B1(n16955), .A0N(n16716), .A1N(n503), .Y(
        n16953) );
  AOI2BB2X1 U11726 ( .B0(n5414), .B1(n16839), .A0N(n112), .A1N(n16703), .Y(
        n16951) );
  NAND4X1 U11727 ( .A(n15061), .B(n15062), .C(n15063), .D(n15064), .Y(n15054)
         );
  AOI2BB2X1 U11728 ( .B0(n3279), .B1(n15065), .A0N(n14826), .A1N(n504), .Y(
        n15063) );
  AOI2BB2X1 U11729 ( .B0(n5878), .B1(n14949), .A0N(n113), .A1N(n14813), .Y(
        n15061) );
  NAND4X1 U11730 ( .A(n16636), .B(n16637), .C(n16638), .D(n16639), .Y(n16629)
         );
  AOI2BB2X1 U11731 ( .B0(n2980), .B1(n16640), .A0N(n16401), .A1N(n505), .Y(
        n16638) );
  AOI2BB2X1 U11732 ( .B0(n5490), .B1(n16524), .A0N(n114), .A1N(n16388), .Y(
        n16636) );
  NAND4X1 U11733 ( .A(n18211), .B(n18212), .C(n18213), .D(n18214), .Y(n18204)
         );
  AOI2BB2X1 U11734 ( .B0(n2675), .B1(n18215), .A0N(n17976), .A1N(n506), .Y(
        n18213) );
  AOI2BB2X1 U11735 ( .B0(n5060), .B1(n18099), .A0N(n115), .A1N(n17963), .Y(
        n18211) );
  NAND4X1 U11736 ( .A(n14746), .B(n14747), .C(n14748), .D(n14749), .Y(n14739)
         );
  AOI2BB2X1 U11737 ( .B0(n3340), .B1(n14750), .A0N(n14511), .A1N(n507), .Y(
        n14748) );
  AOI2BB2X1 U11738 ( .B0(n5954), .B1(n14634), .A0N(n116), .A1N(n14498), .Y(
        n14746) );
  NAND4X1 U11739 ( .A(n16321), .B(n16322), .C(n16323), .D(n16324), .Y(n16314)
         );
  AOI2BB2X1 U11740 ( .B0(n3038), .B1(n16325), .A0N(n16086), .A1N(n508), .Y(
        n16323) );
  AOI2BB2X1 U11741 ( .B0(n5566), .B1(n16209), .A0N(n117), .A1N(n16073), .Y(
        n16321) );
  NAND4X1 U11742 ( .A(n17896), .B(n17897), .C(n17898), .D(n17899), .Y(n17889)
         );
  AOI2BB2X1 U11743 ( .B0(n2735), .B1(n17900), .A0N(n17661), .A1N(n509), .Y(
        n17898) );
  AOI2BB2X1 U11744 ( .B0(n5168), .B1(n17784), .A0N(n118), .A1N(n17648), .Y(
        n17896) );
  NAND4X1 U11745 ( .A(n14431), .B(n14432), .C(n14433), .D(n14434), .Y(n14424)
         );
  AOI2BB2X1 U11746 ( .B0(n3398), .B1(n14435), .A0N(n14196), .A1N(n510), .Y(
        n14433) );
  AOI2BB2X1 U11747 ( .B0(n6030), .B1(n14319), .A0N(n119), .A1N(n14183), .Y(
        n14431) );
  NAND4X1 U11748 ( .A(n16006), .B(n16007), .C(n16008), .D(n16009), .Y(n15999)
         );
  AOI2BB2X1 U11749 ( .B0(n3097), .B1(n16010), .A0N(n15771), .A1N(n511), .Y(
        n16008) );
  AOI2BB2X1 U11750 ( .B0(n5642), .B1(n15894), .A0N(n120), .A1N(n15758), .Y(
        n16006) );
  NAND4X1 U11751 ( .A(n17581), .B(n17582), .C(n17583), .D(n17584), .Y(n17574)
         );
  AOI2BB2X1 U11752 ( .B0(n2798), .B1(n17585), .A0N(n17346), .A1N(n512), .Y(
        n17583) );
  AOI2BB2X1 U11753 ( .B0(n5246), .B1(n17469), .A0N(n121), .A1N(n17333), .Y(
        n17581) );
  NAND4BXL U11754 ( .AN(n17020), .B(n17036), .C(n5382), .D(n17108), .Y(n17105)
         );
  AOI211X1 U11755 ( .A0(n5353), .A1(n370), .B0(n5389), .C0(n17109), .Y(n17108)
         );
  INVX1 U11756 ( .A(n17110), .Y(n5389) );
  AOI21XL U11757 ( .A0(n30), .A1(n17062), .B0(n17061), .Y(n17109) );
  NAND4BXL U11758 ( .AN(n13870), .B(n13886), .C(n6153), .D(n13958), .Y(n13955)
         );
  AOI211X1 U11759 ( .A0(n6121), .A1(n369), .B0(n6171), .C0(n13959), .Y(n13958)
         );
  INVX1 U11760 ( .A(n13960), .Y(n6171) );
  AOI21XL U11761 ( .A0(n31), .A1(n13912), .B0(n13911), .Y(n13959) );
  NAND4BXL U11762 ( .AN(n18280), .B(n18296), .C(n5028), .D(n18368), .Y(n18365)
         );
  AOI211X1 U11763 ( .A0(n4999), .A1(n371), .B0(n5035), .C0(n18369), .Y(n18368)
         );
  INVX1 U11764 ( .A(n18370), .Y(n5035) );
  AOI21XL U11765 ( .A0(n32), .A1(n18322), .B0(n18321), .Y(n18369) );
  NAND4BXL U11766 ( .AN(n15130), .B(n15146), .C(n5854), .D(n15218), .Y(n15215)
         );
  AOI211X1 U11767 ( .A0(n5825), .A1(n372), .B0(n5861), .C0(n15219), .Y(n15218)
         );
  INVX1 U11768 ( .A(n15220), .Y(n5861) );
  AOI21XL U11769 ( .A0(n33), .A1(n15172), .B0(n15171), .Y(n15219) );
  NAND4BXL U11770 ( .AN(n15445), .B(n15461), .C(n5770), .D(n15533), .Y(n15530)
         );
  AOI211X1 U11771 ( .A0(n5741), .A1(n373), .B0(n5777), .C0(n15534), .Y(n15533)
         );
  INVX1 U11772 ( .A(n15535), .Y(n5777) );
  AOI21XL U11773 ( .A0(n34), .A1(n15487), .B0(n15486), .Y(n15534) );
  NAND4BXL U11774 ( .AN(n18595), .B(n18611), .C(n4912), .D(n18683), .Y(n18680)
         );
  AOI211X1 U11775 ( .A0(n4883), .A1(n374), .B0(n4919), .C0(n18684), .Y(n18683)
         );
  INVX1 U11776 ( .A(n18685), .Y(n4919) );
  AOI21XL U11777 ( .A0(n35), .A1(n18637), .B0(n18636), .Y(n18684) );
  NAND4BXL U11778 ( .AN(n16705), .B(n16721), .C(n5466), .D(n16793), .Y(n16790)
         );
  AOI211X1 U11779 ( .A0(n5437), .A1(n375), .B0(n5473), .C0(n16794), .Y(n16793)
         );
  INVX1 U11780 ( .A(n16795), .Y(n5473) );
  AOI21XL U11781 ( .A0(n36), .A1(n16747), .B0(n16746), .Y(n16794) );
  NAND4BXL U11782 ( .AN(n14815), .B(n14831), .C(n5930), .D(n14903), .Y(n14900)
         );
  AOI211X1 U11783 ( .A0(n5901), .A1(n376), .B0(n5937), .C0(n14904), .Y(n14903)
         );
  INVX1 U11784 ( .A(n14905), .Y(n5937) );
  AOI21XL U11785 ( .A0(n37), .A1(n14857), .B0(n14856), .Y(n14904) );
  NAND4BXL U11786 ( .AN(n16390), .B(n16406), .C(n5542), .D(n16478), .Y(n16475)
         );
  AOI211X1 U11787 ( .A0(n5513), .A1(n377), .B0(n5549), .C0(n16479), .Y(n16478)
         );
  INVX1 U11788 ( .A(n16480), .Y(n5549) );
  AOI21XL U11789 ( .A0(n38), .A1(n16432), .B0(n16431), .Y(n16479) );
  NAND4BXL U11790 ( .AN(n17965), .B(n17981), .C(n5112), .D(n18053), .Y(n18050)
         );
  AOI211X1 U11791 ( .A0(n5083), .A1(n378), .B0(n5119), .C0(n18054), .Y(n18053)
         );
  INVX1 U11792 ( .A(n18055), .Y(n5119) );
  AOI21XL U11793 ( .A0(n39), .A1(n18007), .B0(n18006), .Y(n18054) );
  NAND4BXL U11794 ( .AN(n14500), .B(n14516), .C(n6006), .D(n14588), .Y(n14585)
         );
  AOI211X1 U11795 ( .A0(n5977), .A1(n379), .B0(n6013), .C0(n14589), .Y(n14588)
         );
  INVX1 U11796 ( .A(n14590), .Y(n6013) );
  AOI21XL U11797 ( .A0(n40), .A1(n14542), .B0(n14541), .Y(n14589) );
  NAND4BXL U11798 ( .AN(n16075), .B(n16091), .C(n5618), .D(n16163), .Y(n16160)
         );
  AOI211X1 U11799 ( .A0(n5589), .A1(n380), .B0(n5625), .C0(n16164), .Y(n16163)
         );
  INVX1 U11800 ( .A(n16165), .Y(n5625) );
  AOI21XL U11801 ( .A0(n41), .A1(n16117), .B0(n16116), .Y(n16164) );
  NAND4BXL U11802 ( .AN(n17650), .B(n17666), .C(n5220), .D(n17738), .Y(n17735)
         );
  AOI211X1 U11803 ( .A0(n5191), .A1(n381), .B0(n5227), .C0(n17739), .Y(n17738)
         );
  INVX1 U11804 ( .A(n17740), .Y(n5227) );
  AOI21XL U11805 ( .A0(n42), .A1(n17692), .B0(n17691), .Y(n17739) );
  NAND4BXL U11806 ( .AN(n14185), .B(n14201), .C(n6082), .D(n14273), .Y(n14270)
         );
  AOI211X1 U11807 ( .A0(n6053), .A1(n382), .B0(n6089), .C0(n14274), .Y(n14273)
         );
  INVX1 U11808 ( .A(n14275), .Y(n6089) );
  AOI21XL U11809 ( .A0(n43), .A1(n14227), .B0(n14226), .Y(n14274) );
  NAND4BXL U11810 ( .AN(n15760), .B(n15776), .C(n5694), .D(n15848), .Y(n15845)
         );
  AOI211X1 U11811 ( .A0(n5665), .A1(n383), .B0(n5701), .C0(n15849), .Y(n15848)
         );
  INVX1 U11812 ( .A(n15850), .Y(n5701) );
  AOI21XL U11813 ( .A0(n44), .A1(n15802), .B0(n15801), .Y(n15849) );
  NAND4BXL U11814 ( .AN(n17335), .B(n17351), .C(n5298), .D(n17423), .Y(n17420)
         );
  AOI211X1 U11815 ( .A0(n5269), .A1(n384), .B0(n5305), .C0(n17424), .Y(n17423)
         );
  INVX1 U11816 ( .A(n17425), .Y(n5305) );
  AOI21XL U11817 ( .A0(n45), .A1(n17377), .B0(n17376), .Y(n17424) );
  NAND3X1 U11818 ( .A(n17230), .B(n17231), .C(n17232), .Y(n17229) );
  NAND3XL U11819 ( .A(n1311), .B(n17135), .C(n5330), .Y(n17232) );
  NAND3X1 U11820 ( .A(n14080), .B(n14081), .C(n14082), .Y(n14079) );
  NAND3XL U11821 ( .A(n1281), .B(n13985), .C(n6114), .Y(n14082) );
  NAND3X1 U11822 ( .A(n15340), .B(n15341), .C(n15342), .Y(n15339) );
  NAND3XL U11823 ( .A(n1293), .B(n15245), .C(n5802), .Y(n15342) );
  NAND3X1 U11824 ( .A(n18490), .B(n18491), .C(n18492), .Y(n18489) );
  NAND3XL U11825 ( .A(n1323), .B(n18395), .C(n4976), .Y(n18492) );
  NAND3X1 U11826 ( .A(n15655), .B(n15656), .C(n15657), .Y(n15654) );
  NAND3XL U11827 ( .A(n1296), .B(n15560), .C(n5718), .Y(n15657) );
  NAND3X1 U11828 ( .A(n16915), .B(n16916), .C(n16917), .Y(n16914) );
  NAND3XL U11829 ( .A(n1308), .B(n16820), .C(n5414), .Y(n16917) );
  NAND3X1 U11830 ( .A(n18805), .B(n18806), .C(n18807), .Y(n18804) );
  NAND3XL U11831 ( .A(n1326), .B(n18710), .C(n4860), .Y(n18807) );
  NAND3X1 U11832 ( .A(n15025), .B(n15026), .C(n15027), .Y(n15024) );
  NAND3XL U11833 ( .A(n1290), .B(n14930), .C(n5878), .Y(n15027) );
  NAND3X1 U11834 ( .A(n16600), .B(n16601), .C(n16602), .Y(n16599) );
  NAND3XL U11835 ( .A(n1305), .B(n16505), .C(n5490), .Y(n16602) );
  NAND3X1 U11836 ( .A(n18175), .B(n18176), .C(n18177), .Y(n18174) );
  NAND3XL U11837 ( .A(n1320), .B(n18080), .C(n5060), .Y(n18177) );
  NAND3X1 U11838 ( .A(n14710), .B(n14711), .C(n14712), .Y(n14709) );
  NAND3XL U11839 ( .A(n1287), .B(n14615), .C(n5954), .Y(n14712) );
  NAND3X1 U11840 ( .A(n16285), .B(n16286), .C(n16287), .Y(n16284) );
  NAND3XL U11841 ( .A(n1302), .B(n16190), .C(n5566), .Y(n16287) );
  NAND3X1 U11842 ( .A(n17860), .B(n17861), .C(n17862), .Y(n17859) );
  NAND3XL U11843 ( .A(n1317), .B(n17765), .C(n5168), .Y(n17862) );
  NAND3X1 U11844 ( .A(n14395), .B(n14396), .C(n14397), .Y(n14394) );
  NAND3XL U11845 ( .A(n1284), .B(n14300), .C(n6030), .Y(n14397) );
  NAND3X1 U11846 ( .A(n15970), .B(n15971), .C(n15972), .Y(n15969) );
  NAND3XL U11847 ( .A(n1299), .B(n15875), .C(n5642), .Y(n15972) );
  NAND3X1 U11848 ( .A(n17545), .B(n17546), .C(n17547), .Y(n17544) );
  NAND3XL U11849 ( .A(n1314), .B(n17450), .C(n5246), .Y(n17547) );
  BUFX3 U11850 ( .A(n6541), .Y(n1148) );
  INVXL U11851 ( .A(n73), .Y(n6541) );
  BUFX3 U11852 ( .A(n6836), .Y(n1188) );
  INVXL U11853 ( .A(n74), .Y(n6836) );
  BUFX3 U11854 ( .A(n6882), .Y(n1197) );
  INVXL U11855 ( .A(n75), .Y(n6882) );
  CLKINVX3 U11856 ( .A(n765), .Y(n2146) );
  CLKINVX3 U11857 ( .A(n765), .Y(n2147) );
  CLKINVX3 U11858 ( .A(n765), .Y(n2148) );
  CLKINVX3 U11859 ( .A(n765), .Y(n2149) );
  CLKINVX3 U11860 ( .A(n765), .Y(n2150) );
  CLKINVX3 U11861 ( .A(n765), .Y(n2151) );
  CLKINVX3 U11862 ( .A(n765), .Y(n2152) );
  CLKINVX3 U11863 ( .A(n766), .Y(n3509) );
  CLKINVX3 U11864 ( .A(n766), .Y(n3510) );
  CLKINVX3 U11865 ( .A(n766), .Y(n3511) );
  CLKINVX3 U11866 ( .A(n766), .Y(n3512) );
  CLKINVX3 U11867 ( .A(n766), .Y(n3513) );
  CLKINVX3 U11868 ( .A(n766), .Y(n3514) );
  CLKINVX3 U11869 ( .A(n766), .Y(n3515) );
  CLKINVX3 U11870 ( .A(n764), .Y(n2242) );
  CLKINVX3 U11871 ( .A(n764), .Y(n2237) );
  CLKINVX3 U11872 ( .A(n764), .Y(n2243) );
  CLKINVX3 U11873 ( .A(n764), .Y(n2241) );
  CLKINVX3 U11874 ( .A(n764), .Y(n2239) );
  CLKINVX3 U11875 ( .A(n764), .Y(n2238) );
  CLKINVX3 U11876 ( .A(n764), .Y(n2240) );
  CLKINVX3 U11877 ( .A(n740), .Y(n2153) );
  CLKINVX3 U11878 ( .A(n2292), .Y(n2289) );
  CLKINVX3 U11879 ( .A(n3553), .Y(n3549) );
  CLKINVX3 U11880 ( .A(n3553), .Y(n3550) );
  CLKINVX3 U11881 ( .A(n3553), .Y(n3551) );
  CLKINVX3 U11882 ( .A(n3524), .Y(n3517) );
  CLKINVX3 U11883 ( .A(n3525), .Y(n3518) );
  CLKINVX3 U11884 ( .A(n3524), .Y(n3519) );
  CLKINVX3 U11885 ( .A(n3525), .Y(n3520) );
  CLKINVX3 U11886 ( .A(n3524), .Y(n3521) );
  CLKINVX3 U11887 ( .A(n3525), .Y(n3522) );
  CLKINVX3 U11888 ( .A(n3525), .Y(n3523) );
  XOR2X1 U11889 ( .A(top_core_EC_mc_mix_in_8[48]), .B(
        top_core_EC_mc_mix_in_4_48_), .Y(top_core_EC_mc_mix_in_8[49]) );
  XOR2X1 U11890 ( .A(top_core_EC_mc_mix_in_8[48]), .B(
        top_core_EC_mc_mix_in_4_50_), .Y(top_core_EC_mc_mix_in_8[51]) );
  XOR2X1 U11891 ( .A(top_core_EC_mc_mix_in_8[48]), .B(
        top_core_EC_mc_mix_in_4_51_), .Y(top_core_EC_mc_mix_in_8[52]) );
  XOR2X1 U11892 ( .A(top_core_EC_mc_mix_in_8[32]), .B(
        top_core_EC_mc_mix_in_4_32_), .Y(top_core_EC_mc_mix_in_8[33]) );
  XOR2X1 U11893 ( .A(top_core_EC_mc_mix_in_8[32]), .B(
        top_core_EC_mc_mix_in_4_34_), .Y(top_core_EC_mc_mix_in_8[35]) );
  XOR2X1 U11894 ( .A(top_core_EC_mc_mix_in_8[32]), .B(
        top_core_EC_mc_mix_in_4_35_), .Y(top_core_EC_mc_mix_in_8[36]) );
  XOR2X1 U11895 ( .A(top_core_EC_mc_mix_in_8[16]), .B(
        top_core_EC_mc_mix_in_4_16_), .Y(top_core_EC_mc_mix_in_8[17]) );
  NAND3BX1 U11896 ( .AN(n9906), .B(n10162), .C(n10163), .Y(n10161) );
  AOI211X1 U11897 ( .A0(n1615), .A1(n5370), .B0(n5346), .C0(n9927), .Y(n10163)
         );
  INVX1 U11898 ( .A(n9998), .Y(n5370) );
  NAND3BX1 U11899 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n89), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n348), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n349), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n347) );
  AOI211X1 U11900 ( .A0(n1625), .A1(n6160), .B0(n6142), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n112), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n349) );
  INVX1 U11901 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n184), .Y(n6160) );
  NAND3BX1 U11902 ( .AN(n8154), .B(n8410), .C(n8411), .Y(n8409) );
  AOI211X1 U11903 ( .A0(n1621), .A1(n5842), .B0(n5818), .C0(n8175), .Y(n8411)
         );
  INVX1 U11904 ( .A(n8246), .Y(n5842) );
  NAND3BX1 U11905 ( .AN(n11074), .B(n11330), .C(n11331), .Y(n11329) );
  AOI211X1 U11906 ( .A0(n1611), .A1(n5016), .B0(n4992), .C0(n11095), .Y(n11331) );
  INVX1 U11907 ( .A(n11166), .Y(n5016) );
  NAND3BX1 U11908 ( .AN(n10782), .B(n11038), .C(n11039), .Y(n11037) );
  AOI211X1 U11909 ( .A0(n1612), .A1(n5100), .B0(n5076), .C0(n10803), .Y(n11039) );
  INVX1 U11910 ( .A(n10874), .Y(n5100) );
  NAND3BX1 U11911 ( .AN(n7278), .B(n7534), .C(n7535), .Y(n7533) );
  AOI211X1 U11912 ( .A0(n1624), .A1(n6070), .B0(n6046), .C0(n7299), .Y(n7535)
         );
  INVX1 U11913 ( .A(n7370), .Y(n6070) );
  NAND3BX1 U11914 ( .AN(n9030), .B(n9286), .C(n9287), .Y(n9285) );
  AOI211X1 U11915 ( .A0(n1618), .A1(n5606), .B0(n5582), .C0(n9051), .Y(n9287)
         );
  INVX1 U11916 ( .A(n9122), .Y(n5606) );
  NAND3BX1 U11917 ( .AN(n10198), .B(n10454), .C(n10455), .Y(n10453) );
  AOI211X1 U11918 ( .A0(n1614), .A1(n5286), .B0(n5262), .C0(n10219), .Y(n10455) );
  INVX1 U11919 ( .A(n10290), .Y(n5286) );
  NAND3BX1 U11920 ( .AN(n9322), .B(n9578), .C(n9579), .Y(n9577) );
  AOI211X1 U11921 ( .A0(n1617), .A1(n5530), .B0(n5506), .C0(n9343), .Y(n9579)
         );
  INVX1 U11922 ( .A(n9414), .Y(n5530) );
  NAND3BX1 U11923 ( .AN(n8446), .B(n8702), .C(n8703), .Y(n8701) );
  AOI211X1 U11924 ( .A0(n1620), .A1(n5758), .B0(n5734), .C0(n8467), .Y(n8703)
         );
  INVX1 U11925 ( .A(n8538), .Y(n5758) );
  NAND3BX1 U11926 ( .AN(n7570), .B(n7826), .C(n7827), .Y(n7825) );
  AOI211X1 U11927 ( .A0(n1623), .A1(n5994), .B0(n5970), .C0(n7591), .Y(n7827)
         );
  INVX1 U11928 ( .A(n7662), .Y(n5994) );
  NAND3BX1 U11929 ( .AN(n11366), .B(n11622), .C(n11623), .Y(n11621) );
  AOI211X1 U11930 ( .A0(n1610), .A1(n4900), .B0(n4876), .C0(n11387), .Y(n11623) );
  INVX1 U11931 ( .A(n11458), .Y(n4900) );
  NAND3BX1 U11932 ( .AN(n10490), .B(n10746), .C(n10747), .Y(n10745) );
  AOI211X1 U11933 ( .A0(n1613), .A1(n5208), .B0(n5184), .C0(n10511), .Y(n10747) );
  INVX1 U11934 ( .A(n10582), .Y(n5208) );
  NAND3BX1 U11935 ( .AN(n9614), .B(n9870), .C(n9871), .Y(n9869) );
  AOI211X1 U11936 ( .A0(n1616), .A1(n5454), .B0(n5430), .C0(n9635), .Y(n9871)
         );
  INVX1 U11937 ( .A(n9706), .Y(n5454) );
  NAND3BX1 U11938 ( .AN(n8738), .B(n8994), .C(n8995), .Y(n8993) );
  AOI211X1 U11939 ( .A0(n1619), .A1(n5682), .B0(n5658), .C0(n8759), .Y(n8995)
         );
  INVX1 U11940 ( .A(n8830), .Y(n5682) );
  NAND3BX1 U11941 ( .AN(n7862), .B(n8118), .C(n8119), .Y(n8117) );
  AOI211X1 U11942 ( .A0(n1622), .A1(n5918), .B0(n5894), .C0(n7883), .Y(n8119)
         );
  INVX1 U11943 ( .A(n7954), .Y(n5918) );
  CLKINVX3 U11944 ( .A(n739), .Y(n2171) );
  BUFX3 U11945 ( .A(n6557), .Y(n1152) );
  INVXL U11946 ( .A(n180), .Y(n6557) );
  BUFX3 U11947 ( .A(n6898), .Y(n1201) );
  INVXL U11948 ( .A(n182), .Y(n6898) );
  BUFX3 U11949 ( .A(n6852), .Y(n1192) );
  INVXL U11950 ( .A(n181), .Y(n6852) );
  CLKINVX3 U11951 ( .A(n739), .Y(n2172) );
  INVX1 U11952 ( .A(top_core_KE_n2510), .Y(n7008) );
  CLKINVX3 U11953 ( .A(n1607), .Y(n1604) );
  XOR2X1 U11954 ( .A(top_core_EC_mc_n180), .B(top_core_EC_mc_n302), .Y(
        top_core_EC_mc_n301) );
  XOR2X1 U11955 ( .A(top_core_EC_mc_n124), .B(top_core_EC_mc_n237), .Y(
        top_core_EC_mc_n236) );
  XOR2X1 U11956 ( .A(top_core_EC_mc_n783), .B(top_core_EC_mc_n894), .Y(
        top_core_EC_mc_n893) );
  XOR2X1 U11957 ( .A(top_core_EC_mc_n43), .B(top_core_EC_mc_n832), .Y(
        top_core_EC_mc_n831) );
  XOR2X1 U11958 ( .A(top_core_EC_mc_n319), .B(top_core_EC_mc_n461), .Y(
        top_core_EC_mc_n460) );
  XOR2X1 U11959 ( .A(top_core_EC_mc_n60), .B(top_core_EC_mc_n202), .Y(
        top_core_EC_mc_n201) );
  XOR2X1 U11960 ( .A(top_core_EC_mc_n725), .B(top_core_EC_mc_n844), .Y(
        top_core_EC_mc_n843) );
  XOR2X1 U11961 ( .A(top_core_EC_mc_n132), .B(top_core_EC_mc_n245), .Y(
        top_core_EC_mc_n244) );
  XOR2X1 U11962 ( .A(top_core_EC_mc_n791), .B(top_core_EC_mc_n902), .Y(
        top_core_EC_mc_n901) );
  XOR2X1 U11963 ( .A(top_core_EC_mc_n164), .B(top_core_EC_mc_n286), .Y(
        top_core_EC_mc_n285) );
  XOR2X1 U11964 ( .A(top_core_EC_mc_n140), .B(top_core_EC_mc_n262), .Y(
        top_core_EC_mc_n261) );
  XOR2X1 U11965 ( .A(top_core_EC_mc_n799), .B(top_core_EC_mc_n910), .Y(
        top_core_EC_mc_n909) );
  XOR2X1 U11966 ( .A(top_core_EC_mc_n25), .B(top_core_EC_mc_n820), .Y(
        top_core_EC_mc_n819) );
  XOR2X1 U11967 ( .A(top_core_EC_mc_n318), .B(top_core_EC_mc_n319), .Y(
        top_core_EC_mc_n317) );
  XOR2X1 U11968 ( .A(top_core_EC_mc_n172), .B(top_core_EC_mc_n294), .Y(
        top_core_EC_mc_n293) );
  XOR2X1 U11969 ( .A(top_core_EC_mc_n156), .B(top_core_EC_mc_n278), .Y(
        top_core_EC_mc_n277) );
  XOR2X1 U11970 ( .A(top_core_EC_mc_n148), .B(top_core_EC_mc_n270), .Y(
        top_core_EC_mc_n269) );
  XOR2X1 U11971 ( .A(top_core_EC_mc_n16), .B(top_core_EC_mc_n814), .Y(
        top_core_EC_mc_n813) );
  XOR2X1 U11972 ( .A(top_core_EC_mc_n310), .B(top_core_EC_mc_n311), .Y(
        top_core_EC_mc_n309) );
  XOR2X1 U11973 ( .A(top_core_EC_mc_n376), .B(top_core_EC_mc_n491), .Y(
        top_core_EC_mc_n490) );
  XOR2X1 U11974 ( .A(top_core_EC_mc_n179), .B(top_core_EC_mc_n180), .Y(
        top_core_EC_mc_n178) );
  XOR2X1 U11975 ( .A(top_core_EC_mc_n163), .B(top_core_EC_mc_n164), .Y(
        top_core_EC_mc_n162) );
  XOR2X1 U11976 ( .A(top_core_EC_mc_n155), .B(top_core_EC_mc_n156), .Y(
        top_core_EC_mc_n154) );
  XOR2X1 U11977 ( .A(top_core_EC_mc_n147), .B(top_core_EC_mc_n148), .Y(
        top_core_EC_mc_n146) );
  XOR2X1 U11978 ( .A(top_core_EC_mc_n139), .B(top_core_EC_mc_n140), .Y(
        top_core_EC_mc_n138) );
  XOR2X1 U11979 ( .A(top_core_EC_mc_n131), .B(top_core_EC_mc_n132), .Y(
        top_core_EC_mc_n130) );
  XOR2X1 U11980 ( .A(top_core_EC_mc_n123), .B(top_core_EC_mc_n124), .Y(
        top_core_EC_mc_n122) );
  XOR2X1 U11981 ( .A(top_core_EC_mc_n116), .B(top_core_EC_mc_n117), .Y(
        top_core_EC_mc_n115) );
  XOR2X1 U11982 ( .A(top_core_EC_mc_n59), .B(top_core_EC_mc_n60), .Y(
        top_core_EC_mc_n58) );
  XOR2X1 U11983 ( .A(top_core_EC_mc_n51), .B(top_core_EC_mc_n52), .Y(
        top_core_EC_mc_n50) );
  XOR2X1 U11984 ( .A(top_core_EC_mc_n807), .B(top_core_EC_mc_n918), .Y(
        top_core_EC_mc_n917) );
  XOR2X1 U11985 ( .A(top_core_EC_mc_n117), .B(top_core_EC_mc_n232), .Y(
        top_core_EC_mc_n231) );
  XOR2X1 U11986 ( .A(top_core_EC_mc_n171), .B(top_core_EC_mc_n172), .Y(
        top_core_EC_mc_n170) );
  XOR2X1 U11987 ( .A(top_core_EC_mc_n42), .B(top_core_EC_mc_n43), .Y(
        top_core_EC_mc_n41) );
  XOR2X1 U11988 ( .A(top_core_EC_mc_n33), .B(top_core_EC_mc_n34), .Y(
        top_core_EC_mc_n32) );
  XOR2X1 U11989 ( .A(top_core_EC_mc_n24), .B(top_core_EC_mc_n25), .Y(
        top_core_EC_mc_n23) );
  XOR2X1 U11990 ( .A(top_core_EC_mc_n15), .B(top_core_EC_mc_n16), .Y(
        top_core_EC_mc_n14) );
  XOR2X1 U11991 ( .A(top_core_EC_mc_n34), .B(top_core_EC_mc_n826), .Y(
        top_core_EC_mc_n825) );
  XOR2X1 U11992 ( .A(top_core_EC_mc_n770), .B(top_core_EC_mc_n887), .Y(
        top_core_EC_mc_n886) );
  XOR2X1 U11993 ( .A(top_core_EC_mc_n806), .B(top_core_EC_mc_n807), .Y(
        top_core_EC_mc_n805) );
  XOR2X1 U11994 ( .A(top_core_EC_mc_n798), .B(top_core_EC_mc_n799), .Y(
        top_core_EC_mc_n797) );
  XOR2X1 U11995 ( .A(top_core_EC_mc_n790), .B(top_core_EC_mc_n791), .Y(
        top_core_EC_mc_n789) );
  XOR2X1 U11996 ( .A(top_core_EC_mc_n782), .B(top_core_EC_mc_n783), .Y(
        top_core_EC_mc_n781) );
  XOR2X1 U11997 ( .A(top_core_EC_mc_n769), .B(top_core_EC_mc_n770), .Y(
        top_core_EC_mc_n768) );
  XOR2X1 U11998 ( .A(top_core_EC_mc_n724), .B(top_core_EC_mc_n725), .Y(
        top_core_EC_mc_n723) );
  XOR2X1 U11999 ( .A(top_core_EC_mc_n716), .B(top_core_EC_mc_n717), .Y(
        top_core_EC_mc_n715) );
  XOR2X1 U12000 ( .A(top_core_EC_mc_n311), .B(top_core_EC_mc_n456), .Y(
        top_core_EC_mc_n455) );
  XOR2X1 U12001 ( .A(top_core_EC_mc_n52), .B(top_core_EC_mc_n197), .Y(
        top_core_EC_mc_n196) );
  XOR2X1 U12002 ( .A(top_core_EC_mc_n717), .B(top_core_EC_mc_n839), .Y(
        top_core_EC_mc_n838) );
  XOR2X1 U12003 ( .A(n1550), .B(top_core_EC_mc_mix_in_4_10_), .Y(
        top_core_EC_mc_mix_in_8[11]) );
  XOR2X1 U12004 ( .A(n1547), .B(top_core_EC_mc_mix_in_4_26_), .Y(
        top_core_EC_mc_mix_in_8[27]) );
  INVX1 U12005 ( .A(n11919), .Y(n6825) );
  INVX1 U12006 ( .A(top_core_KE_sb1_n348), .Y(n6803) );
  INVX1 U12007 ( .A(n12550), .Y(n6529) );
  INVX1 U12008 ( .A(n13495), .Y(n6471) );
  INVX1 U12009 ( .A(n12235), .Y(n6506) );
  INVX1 U12010 ( .A(n13180), .Y(n6814) );
  INVX1 U12011 ( .A(n13810), .Y(n6518) );
  INVX1 U12012 ( .A(n12865), .Y(n6774) );
  XOR2X1 U12013 ( .A(n1547), .B(n1546), .Y(top_core_EC_mc_mix_in_8[25]) );
  XOR2X1 U12014 ( .A(n1547), .B(top_core_EC_mc_mix_in_4_27_), .Y(
        top_core_EC_mc_mix_in_8[28]) );
  XOR2X1 U12015 ( .A(n1550), .B(top_core_EC_mc_mix_in_4_11_), .Y(
        top_core_EC_mc_mix_in_8[12]) );
  CLKINVX3 U12016 ( .A(n2273), .Y(n2270) );
  CLKINVX3 U12017 ( .A(n2272), .Y(n2267) );
  CLKINVX3 U12018 ( .A(n2273), .Y(n2269) );
  CLKINVX3 U12019 ( .A(n2272), .Y(n2271) );
  CLKINVX3 U12020 ( .A(n2273), .Y(n2268) );
  CLKINVX3 U12021 ( .A(n2273), .Y(n2265) );
  CLKINVX3 U12022 ( .A(n2272), .Y(n2266) );
  AND2X2 U12023 ( .A(n3467), .B(n6174), .Y(n585) );
  AND2X2 U12024 ( .A(n2866), .B(n5387), .Y(n586) );
  AND2X2 U12025 ( .A(n2624), .B(n5033), .Y(n587) );
  AND2X2 U12026 ( .A(n3226), .B(n5859), .Y(n588) );
  AND2X2 U12027 ( .A(n2685), .B(n5117), .Y(n589) );
  AND2X2 U12028 ( .A(n3046), .B(n5623), .Y(n590) );
  AND2X2 U12029 ( .A(n3406), .B(n6087), .Y(n591) );
  AND2X2 U12030 ( .A(n2806), .B(n5303), .Y(n592) );
  AND2X2 U12031 ( .A(n2988), .B(n5547), .Y(n593) );
  AND2X2 U12032 ( .A(n3165), .B(n5775), .Y(n594) );
  AND2X2 U12033 ( .A(n3348), .B(n6011), .Y(n595) );
  AND2X2 U12034 ( .A(n2563), .B(n4917), .Y(n596) );
  AND2X2 U12035 ( .A(n2745), .B(n5225), .Y(n597) );
  AND2X2 U12036 ( .A(n2927), .B(n5471), .Y(n598) );
  AND2X2 U12037 ( .A(n3107), .B(n5699), .Y(n599) );
  AND2X2 U12038 ( .A(n3287), .B(n5935), .Y(n600) );
  XOR2X1 U12039 ( .A(top_core_EC_mc_mix_in_8[0]), .B(
        top_core_EC_mc_mix_in_4_2_), .Y(top_core_EC_mc_mix_in_8[3]) );
  XOR2X1 U12040 ( .A(top_core_EC_mc_mix_in_8[0]), .B(
        top_core_EC_mc_mix_in_4_3_), .Y(top_core_EC_mc_mix_in_8[4]) );
  INVX1 U12041 ( .A(n11725), .Y(n6913) );
  INVX1 U12042 ( .A(top_core_KE_sb1_n152), .Y(n6867) );
  INVX1 U12043 ( .A(n12356), .Y(n6620) );
  INVX1 U12044 ( .A(n12041), .Y(n6573) );
  CLKINVX3 U12045 ( .A(n3553), .Y(n3552) );
  INVX1 U12046 ( .A(top_core_EC_mix_out_58_), .Y(n4947) );
  OAI22X1 U12047 ( .A0(top_core_EC_mc_n355), .A1(n2441), .B0(n2381), .B1(
        top_core_EC_mc_n356), .Y(top_core_EC_mix_out_58_) );
  XOR2X1 U12048 ( .A(top_core_EC_mc_n357), .B(top_core_EC_mc_n358), .Y(
        top_core_EC_mc_n356) );
  XNOR2X1 U12049 ( .A(top_core_EC_mc_mix_in_2_58_), .B(top_core_EC_mc_n359), 
        .Y(top_core_EC_mc_n355) );
  INVX1 U12050 ( .A(top_core_EC_mix_out_59_), .Y(n4942) );
  OAI22X1 U12051 ( .A0(top_core_EC_mc_n347), .A1(n2443), .B0(n2381), .B1(
        top_core_EC_mc_n348), .Y(top_core_EC_mix_out_59_) );
  XOR2X1 U12052 ( .A(top_core_EC_mc_n349), .B(top_core_EC_mc_n350), .Y(
        top_core_EC_mc_n348) );
  XNOR2X1 U12053 ( .A(top_core_EC_mc_mix_in_2_59_), .B(top_core_EC_mc_n351), 
        .Y(top_core_EC_mc_n347) );
  INVX1 U12054 ( .A(top_core_EC_mix_out_60_), .Y(n4952) );
  OAI22X1 U12055 ( .A0(top_core_EC_mc_n330), .A1(n2428), .B0(n2381), .B1(
        top_core_EC_mc_n331), .Y(top_core_EC_mix_out_60_) );
  XOR2X1 U12056 ( .A(top_core_EC_mc_n332), .B(top_core_EC_mc_n333), .Y(
        top_core_EC_mc_n331) );
  XNOR2X1 U12057 ( .A(top_core_EC_mc_mix_in_8[62]), .B(top_core_EC_mc_n334), 
        .Y(top_core_EC_mc_n330) );
  INVX1 U12058 ( .A(top_core_EC_mix_out_73_), .Y(n4797) );
  OAI22X1 U12059 ( .A0(top_core_EC_mc_n223), .A1(n2366), .B0(n2382), .B1(
        top_core_EC_mc_n224), .Y(top_core_EC_mix_out_73_) );
  XOR2X1 U12060 ( .A(top_core_EC_mc_n225), .B(top_core_EC_mc_n226), .Y(
        top_core_EC_mc_n224) );
  XNOR2X1 U12061 ( .A(top_core_EC_mc_mix_in_4_74_), .B(top_core_EC_mc_n227), 
        .Y(top_core_EC_mc_n223) );
  INVX1 U12062 ( .A(top_core_EC_mix_out_75_), .Y(n4794) );
  OAI22X1 U12063 ( .A0(top_core_EC_mc_n213), .A1(n2527), .B0(n2383), .B1(
        top_core_EC_mc_n214), .Y(top_core_EC_mix_out_75_) );
  XOR2X1 U12064 ( .A(top_core_EC_mc_n215), .B(top_core_EC_mc_n216), .Y(
        top_core_EC_mc_n214) );
  XNOR2X1 U12065 ( .A(top_core_EC_mc_mix_in_2_75_), .B(top_core_EC_mc_n217), 
        .Y(top_core_EC_mc_n213) );
  INVX1 U12066 ( .A(top_core_EC_mix_out_76_), .Y(n4786) );
  OAI22X1 U12067 ( .A0(top_core_EC_mc_n208), .A1(n2442), .B0(n2383), .B1(
        top_core_EC_mc_n209), .Y(top_core_EC_mix_out_76_) );
  XOR2X1 U12068 ( .A(top_core_EC_mc_n210), .B(top_core_EC_mc_n211), .Y(
        top_core_EC_mc_n209) );
  XNOR2X1 U12069 ( .A(top_core_EC_mc_mix_in_8[78]), .B(top_core_EC_mc_n212), 
        .Y(top_core_EC_mc_n208) );
  INVX1 U12070 ( .A(top_core_EC_mix_out_81_), .Y(n4792) );
  OAI22X1 U12071 ( .A0(top_core_EC_mc_n168), .A1(n2541), .B0(n2383), .B1(
        top_core_EC_mc_n169), .Y(top_core_EC_mix_out_81_) );
  XOR2X1 U12072 ( .A(top_core_EC_mc_n106), .B(top_core_EC_mc_n170), .Y(
        top_core_EC_mc_n169) );
  XNOR2X1 U12073 ( .A(top_core_EC_mc_mix_in_4_90_), .B(top_core_EC_mc_n171), 
        .Y(top_core_EC_mc_n168) );
  INVX1 U12074 ( .A(top_core_EC_mix_out_83_), .Y(n4789) );
  OAI22X1 U12075 ( .A0(top_core_EC_mc_n152), .A1(n2411), .B0(n2383), .B1(
        top_core_EC_mc_n153), .Y(top_core_EC_mix_out_83_) );
  XOR2X1 U12076 ( .A(top_core_EC_mc_n81), .B(top_core_EC_mc_n154), .Y(
        top_core_EC_mc_n153) );
  XNOR2X1 U12077 ( .A(top_core_EC_mc_mix_in_2_91_), .B(top_core_EC_mc_n155), 
        .Y(top_core_EC_mc_n152) );
  INVX1 U12078 ( .A(top_core_EC_mix_out_84_), .Y(n4779) );
  OAI22X1 U12079 ( .A0(top_core_EC_mc_n144), .A1(n2540), .B0(n2383), .B1(
        top_core_EC_mc_n145), .Y(top_core_EC_mix_out_84_) );
  XOR2X1 U12080 ( .A(top_core_EC_mc_n73), .B(top_core_EC_mc_n146), .Y(
        top_core_EC_mc_n145) );
  XNOR2X1 U12081 ( .A(top_core_EC_mc_mix_in_8[94]), .B(top_core_EC_mc_n147), 
        .Y(top_core_EC_mc_n144) );
  INVX1 U12082 ( .A(top_core_EC_mix_out_89_), .Y(n4791) );
  OAI22X1 U12083 ( .A0(top_core_EC_mc_n104), .A1(n2399), .B0(n2384), .B1(
        top_core_EC_mc_n105), .Y(top_core_EC_mix_out_89_) );
  XOR2X1 U12084 ( .A(top_core_EC_mc_n106), .B(top_core_EC_mc_n107), .Y(
        top_core_EC_mc_n105) );
  XNOR2X1 U12085 ( .A(top_core_EC_mc_mix_in_4_90_), .B(top_core_EC_mc_n108), 
        .Y(top_core_EC_mc_n104) );
  INVX1 U12086 ( .A(top_core_EC_mix_out_91_), .Y(n4790) );
  OAI22X1 U12087 ( .A0(top_core_EC_mc_n79), .A1(n2430), .B0(n2384), .B1(
        top_core_EC_mc_n80), .Y(top_core_EC_mix_out_91_) );
  XOR2X1 U12088 ( .A(top_core_EC_mc_n81), .B(top_core_EC_mc_n82), .Y(
        top_core_EC_mc_n80) );
  XNOR2X1 U12089 ( .A(top_core_EC_mc_mix_in_2_91_), .B(top_core_EC_mc_n83), 
        .Y(top_core_EC_mc_n79) );
  INVX1 U12090 ( .A(top_core_EC_mix_out_92_), .Y(n4778) );
  OAI22X1 U12091 ( .A0(top_core_EC_mc_n71), .A1(n2400), .B0(n2380), .B1(
        top_core_EC_mc_n72), .Y(top_core_EC_mix_out_92_) );
  XOR2X1 U12092 ( .A(top_core_EC_mc_n73), .B(top_core_EC_mc_n74), .Y(
        top_core_EC_mc_n72) );
  XNOR2X1 U12093 ( .A(top_core_EC_mc_mix_in_8[94]), .B(top_core_EC_mc_n75), 
        .Y(top_core_EC_mc_n71) );
  INVX1 U12094 ( .A(top_core_EC_mix_out_105_), .Y(n5152) );
  OAI22X1 U12095 ( .A0(top_core_EC_mc_n876), .A1(n2530), .B0(n2376), .B1(
        top_core_EC_mc_n877), .Y(top_core_EC_mix_out_105_) );
  XOR2X1 U12096 ( .A(top_core_EC_mc_n878), .B(top_core_EC_mc_n879), .Y(
        top_core_EC_mc_n877) );
  XNOR2X1 U12097 ( .A(top_core_EC_mc_mix_in_4_106_), .B(top_core_EC_mc_n880), 
        .Y(top_core_EC_mc_n876) );
  INVX1 U12098 ( .A(top_core_EC_mix_out_107_), .Y(n5141) );
  OAI22X1 U12099 ( .A0(top_core_EC_mc_n862), .A1(n2529), .B0(n2376), .B1(
        top_core_EC_mc_n863), .Y(top_core_EC_mix_out_107_) );
  XOR2X1 U12100 ( .A(top_core_EC_mc_n864), .B(top_core_EC_mc_n865), .Y(
        top_core_EC_mc_n863) );
  XNOR2X1 U12101 ( .A(top_core_EC_mc_mix_in_2_107_), .B(top_core_EC_mc_n866), 
        .Y(top_core_EC_mc_n862) );
  INVX1 U12102 ( .A(top_core_EC_mix_out_108_), .Y(n5151) );
  OAI22X1 U12103 ( .A0(top_core_EC_mc_n857), .A1(n2477), .B0(n2376), .B1(
        top_core_EC_mc_n858), .Y(top_core_EC_mix_out_108_) );
  XOR2X1 U12104 ( .A(top_core_EC_mc_n859), .B(top_core_EC_mc_n860), .Y(
        top_core_EC_mc_n858) );
  XNOR2X1 U12105 ( .A(top_core_EC_mc_mix_in_8[110]), .B(top_core_EC_mc_n861), 
        .Y(top_core_EC_mc_n857) );
  INVX1 U12106 ( .A(top_core_EC_mix_out_113_), .Y(n5145) );
  OAI22X1 U12107 ( .A0(top_core_EC_mc_n823), .A1(n2446), .B0(n2376), .B1(
        top_core_EC_mc_n824), .Y(top_core_EC_mix_out_113_) );
  XOR2X1 U12108 ( .A(top_core_EC_mc_n760), .B(top_core_EC_mc_n825), .Y(
        top_core_EC_mc_n824) );
  XNOR2X1 U12109 ( .A(top_core_EC_mc_mix_in_4_122_), .B(top_core_EC_mc_n826), 
        .Y(top_core_EC_mc_n823) );
  INVX1 U12110 ( .A(top_core_EC_mix_out_115_), .Y(n5142) );
  OAI22X1 U12111 ( .A0(top_core_EC_mc_n811), .A1(n2442), .B0(n2376), .B1(
        top_core_EC_mc_n812), .Y(top_core_EC_mix_out_115_) );
  XOR2X1 U12112 ( .A(top_core_EC_mc_n746), .B(top_core_EC_mc_n813), .Y(
        top_core_EC_mc_n812) );
  XNOR2X1 U12113 ( .A(top_core_EC_mc_mix_in_2_123_), .B(top_core_EC_mc_n814), 
        .Y(top_core_EC_mc_n811) );
  INVX1 U12114 ( .A(top_core_EC_mix_out_116_), .Y(n5134) );
  OAI22X1 U12115 ( .A0(top_core_EC_mc_n803), .A1(n2412), .B0(n2376), .B1(
        top_core_EC_mc_n804), .Y(top_core_EC_mix_out_116_) );
  XOR2X1 U12116 ( .A(top_core_EC_mc_n738), .B(top_core_EC_mc_n805), .Y(
        top_core_EC_mc_n804) );
  XNOR2X1 U12117 ( .A(top_core_EC_mc_mix_in_8[126]), .B(top_core_EC_mc_n806), 
        .Y(top_core_EC_mc_n803) );
  INVX1 U12118 ( .A(top_core_EC_mix_out_121_), .Y(n5139) );
  OAI22X1 U12119 ( .A0(top_core_EC_mc_n758), .A1(n2418), .B0(n2377), .B1(
        top_core_EC_mc_n759), .Y(top_core_EC_mix_out_121_) );
  XOR2X1 U12120 ( .A(top_core_EC_mc_n760), .B(top_core_EC_mc_n761), .Y(
        top_core_EC_mc_n759) );
  XNOR2X1 U12121 ( .A(top_core_EC_mc_mix_in_4_122_), .B(top_core_EC_mc_n762), 
        .Y(top_core_EC_mc_n758) );
  INVX1 U12122 ( .A(top_core_EC_mix_out_123_), .Y(n5137) );
  OAI22X1 U12123 ( .A0(top_core_EC_mc_n744), .A1(n2419), .B0(n2377), .B1(
        top_core_EC_mc_n745), .Y(top_core_EC_mix_out_123_) );
  XOR2X1 U12124 ( .A(top_core_EC_mc_n746), .B(top_core_EC_mc_n747), .Y(
        top_core_EC_mc_n745) );
  XNOR2X1 U12125 ( .A(top_core_EC_mc_mix_in_2_123_), .B(top_core_EC_mc_n748), 
        .Y(top_core_EC_mc_n744) );
  INVX1 U12126 ( .A(top_core_EC_mix_out_124_), .Y(n5127) );
  OAI22X1 U12127 ( .A0(top_core_EC_mc_n736), .A1(n2489), .B0(n2377), .B1(
        top_core_EC_mc_n737), .Y(top_core_EC_mix_out_124_) );
  XOR2X1 U12128 ( .A(top_core_EC_mc_n738), .B(top_core_EC_mc_n739), .Y(
        top_core_EC_mc_n737) );
  XNOR2X1 U12129 ( .A(top_core_EC_mc_mix_in_8[126]), .B(top_core_EC_mc_n740), 
        .Y(top_core_EC_mc_n736) );
  INVX1 U12130 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n145), .Y(n6168) );
  INVX1 U12131 ( .A(n9960), .Y(n5383) );
  INVX1 U12132 ( .A(n11128), .Y(n5029) );
  INVX1 U12133 ( .A(n8208), .Y(n5855) );
  INVX1 U12134 ( .A(n10836), .Y(n5113) );
  INVX1 U12135 ( .A(n9084), .Y(n5619) );
  INVX1 U12136 ( .A(n7332), .Y(n6083) );
  INVX1 U12137 ( .A(n10252), .Y(n5299) );
  INVX1 U12138 ( .A(n9376), .Y(n5543) );
  INVX1 U12139 ( .A(n8500), .Y(n5771) );
  INVX1 U12140 ( .A(n7624), .Y(n6007) );
  INVX1 U12141 ( .A(n11420), .Y(n4913) );
  INVX1 U12142 ( .A(n10544), .Y(n5221) );
  INVX1 U12143 ( .A(n9668), .Y(n5467) );
  INVX1 U12144 ( .A(n8792), .Y(n5695) );
  INVX1 U12145 ( .A(n7916), .Y(n5931) );
  BUFX3 U12146 ( .A(n6555), .Y(n1151) );
  INVXL U12147 ( .A(n3), .Y(n6555) );
  BUFX3 U12148 ( .A(n6850), .Y(n1191) );
  INVXL U12149 ( .A(n4), .Y(n6850) );
  BUFX3 U12150 ( .A(n6896), .Y(n1200) );
  INVXL U12151 ( .A(n5), .Y(n6896) );
  XNOR2X1 U12152 ( .A(top_core_EC_mc_mix_in_4_74_), .B(top_core_EC_mc_n173), 
        .Y(top_core_EC_mc_n225) );
  XNOR2X1 U12153 ( .A(top_core_EC_mc_mix_in_4_106_), .B(top_core_EC_mc_n35), 
        .Y(top_core_EC_mc_n878) );
  AOI221X1 U12154 ( .A0(n5026), .A1(n947), .B0(n18435), .B1(n946), .C0(n18502), 
        .Y(n18501) );
  AOI21XL U12155 ( .A0(n108), .A1(n18350), .B0(n2649), .Y(n18502) );
  AOI221X1 U12156 ( .A0(n5768), .A1(n1073), .B0(n15600), .B1(n1072), .C0(
        n15667), .Y(n15666) );
  AOI21XL U12157 ( .A0(n110), .A1(n15515), .B0(n3183), .Y(n15667) );
  AOI221X1 U12158 ( .A0(n5380), .A1(n1003), .B0(n17175), .B1(n1002), .C0(
        n17242), .Y(n17241) );
  AOI21XL U12159 ( .A0(n106), .A1(n17090), .B0(n2890), .Y(n17242) );
  AOI221X1 U12160 ( .A0(n6151), .A1(n1142), .B0(n14025), .B1(n1141), .C0(
        n14092), .Y(n14091) );
  AOI21XL U12161 ( .A0(n107), .A1(n13940), .B0(n3487), .Y(n14092) );
  AOI221X1 U12162 ( .A0(n5852), .A1(n1087), .B0(n15285), .B1(n1086), .C0(
        n15352), .Y(n15351) );
  AOI21XL U12163 ( .A0(n109), .A1(n15200), .B0(n3247), .Y(n15352) );
  AOI221X1 U12164 ( .A0(n5464), .A1(n1017), .B0(n16860), .B1(n1016), .C0(
        n16927), .Y(n16926) );
  AOI21XL U12165 ( .A0(n112), .A1(n16775), .B0(n2952), .Y(n16927) );
  AOI221X1 U12166 ( .A0(n4910), .A1(n933), .B0(n18750), .B1(n932), .C0(n18817), 
        .Y(n18816) );
  AOI21XL U12167 ( .A0(n111), .A1(n18665), .B0(n2581), .Y(n18817) );
  AOI221X1 U12168 ( .A0(n5928), .A1(n1101), .B0(n14970), .B1(n1100), .C0(
        n15037), .Y(n15036) );
  AOI21XL U12169 ( .A0(n113), .A1(n14885), .B0(n3308), .Y(n15037) );
  AOI221X1 U12170 ( .A0(n5540), .A1(n1031), .B0(n16545), .B1(n1030), .C0(
        n16612), .Y(n16611) );
  AOI21XL U12171 ( .A0(n114), .A1(n16460), .B0(n3009), .Y(n16612) );
  AOI221X1 U12172 ( .A0(n5110), .A1(n961), .B0(n18120), .B1(n960), .C0(n18187), 
        .Y(n18186) );
  AOI21XL U12173 ( .A0(n115), .A1(n18035), .B0(n2703), .Y(n18187) );
  AOI221X1 U12174 ( .A0(n6004), .A1(n1115), .B0(n14655), .B1(n1114), .C0(
        n14722), .Y(n14721) );
  AOI21XL U12175 ( .A0(n116), .A1(n14570), .B0(n3366), .Y(n14722) );
  AOI221X1 U12176 ( .A0(n5616), .A1(n1045), .B0(n16230), .B1(n1044), .C0(
        n16297), .Y(n16296) );
  AOI21XL U12177 ( .A0(n117), .A1(n16145), .B0(n3071), .Y(n16297) );
  AOI221X1 U12178 ( .A0(n5218), .A1(n975), .B0(n17805), .B1(n974), .C0(n17872), 
        .Y(n17871) );
  AOI21XL U12179 ( .A0(n118), .A1(n17720), .B0(n2763), .Y(n17872) );
  AOI221X1 U12180 ( .A0(n6080), .A1(n1129), .B0(n14340), .B1(n1128), .C0(
        n14407), .Y(n14406) );
  AOI21XL U12181 ( .A0(n119), .A1(n14255), .B0(n3431), .Y(n14407) );
  AOI221X1 U12182 ( .A0(n5692), .A1(n1059), .B0(n15915), .B1(n1058), .C0(
        n15982), .Y(n15981) );
  AOI21XL U12183 ( .A0(n120), .A1(n15830), .B0(n3125), .Y(n15982) );
  AOI221X1 U12184 ( .A0(n5296), .A1(n989), .B0(n17490), .B1(n988), .C0(n17557), 
        .Y(n17556) );
  AOI21XL U12185 ( .A0(n121), .A1(n17405), .B0(n2831), .Y(n17557) );
  XNOR2X1 U12186 ( .A(top_core_EC_mc_mix_in_8[78]), .B(top_core_EC_mc_n149), 
        .Y(top_core_EC_mc_n210) );
  XNOR2X1 U12187 ( .A(top_core_EC_mc_mix_in_8[110]), .B(top_core_EC_mc_n808), 
        .Y(top_core_EC_mc_n859) );
  XNOR2X1 U12188 ( .A(top_core_EC_mc_mix_in_2_75_), .B(top_core_EC_mc_n157), 
        .Y(top_core_EC_mc_n215) );
  XNOR2X1 U12189 ( .A(top_core_EC_mc_mix_in_2_107_), .B(top_core_EC_mc_n17), 
        .Y(top_core_EC_mc_n864) );
  NAND2X1 U12190 ( .A(n9917), .B(n10068), .Y(n10067) );
  NAND2X1 U12191 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n101), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n254), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n253) );
  NAND2X1 U12192 ( .A(n11085), .B(n11236), .Y(n11235) );
  NAND2X1 U12193 ( .A(n8165), .B(n8316), .Y(n8315) );
  NAND2X1 U12194 ( .A(n10793), .B(n10944), .Y(n10943) );
  NAND2X1 U12195 ( .A(n7289), .B(n7440), .Y(n7439) );
  NAND2X1 U12196 ( .A(n9041), .B(n9192), .Y(n9191) );
  NAND2X1 U12197 ( .A(n10209), .B(n10360), .Y(n10359) );
  NAND2X1 U12198 ( .A(n9333), .B(n9484), .Y(n9483) );
  NAND2X1 U12199 ( .A(n8457), .B(n8608), .Y(n8607) );
  NAND2X1 U12200 ( .A(n7581), .B(n7732), .Y(n7731) );
  NAND2X1 U12201 ( .A(n11377), .B(n11528), .Y(n11527) );
  NAND2X1 U12202 ( .A(n10501), .B(n10652), .Y(n10651) );
  NAND2X1 U12203 ( .A(n9625), .B(n9776), .Y(n9775) );
  NAND2X1 U12204 ( .A(n8749), .B(n8900), .Y(n8899) );
  NAND2X1 U12205 ( .A(n7873), .B(n8024), .Y(n8023) );
  XOR2X1 U12206 ( .A(n1550), .B(n1549), .Y(top_core_EC_mc_mix_in_8[9]) );
  AOI21X1 U12207 ( .A0(n17193), .A1(n17194), .B0(n2852), .Y(n17192) );
  AOI21X1 U12208 ( .A0(n14043), .A1(n14044), .B0(n3453), .Y(n14042) );
  AOI21X1 U12209 ( .A0(n18453), .A1(n18454), .B0(n2610), .Y(n18452) );
  AOI21X1 U12210 ( .A0(n15303), .A1(n15304), .B0(n3212), .Y(n15302) );
  AOI21X1 U12211 ( .A0(n15618), .A1(n15619), .B0(n3151), .Y(n15617) );
  AOI21X1 U12212 ( .A0(n16878), .A1(n16879), .B0(n2913), .Y(n16877) );
  AOI21X1 U12213 ( .A0(n18768), .A1(n18769), .B0(n2549), .Y(n18767) );
  AOI21X1 U12214 ( .A0(n14988), .A1(n14989), .B0(n3273), .Y(n14987) );
  AOI21X1 U12215 ( .A0(n16563), .A1(n16564), .B0(n2974), .Y(n16562) );
  AOI21X1 U12216 ( .A0(n18138), .A1(n18139), .B0(n2671), .Y(n18137) );
  AOI21X1 U12217 ( .A0(n14673), .A1(n14674), .B0(n3334), .Y(n14672) );
  AOI21X1 U12218 ( .A0(n16248), .A1(n16249), .B0(n3032), .Y(n16247) );
  AOI21X1 U12219 ( .A0(n17823), .A1(n17824), .B0(n2731), .Y(n17822) );
  AOI21X1 U12220 ( .A0(n14358), .A1(n14359), .B0(n3392), .Y(n14357) );
  AOI21X1 U12221 ( .A0(n15933), .A1(n15934), .B0(n3093), .Y(n15932) );
  AOI21X1 U12222 ( .A0(n17508), .A1(n17509), .B0(n2792), .Y(n17507) );
  AOI221X1 U12223 ( .A0(n2847), .A1(n17050), .B0(n17051), .B1(n17052), .C0(
        n17053), .Y(n17049) );
  AOI21X1 U12224 ( .A0(n17054), .A1(n17055), .B0(n17056), .Y(n17053) );
  NAND4X1 U12225 ( .A(n17013), .B(n17062), .C(n17063), .D(n17064), .Y(n17052)
         );
  OAI221XL U12226 ( .A0(n5354), .A1(n2852), .B0(n2859), .B1(n17066), .C0(
        n17067), .Y(n17050) );
  AOI221X1 U12227 ( .A0(n3448), .A1(n13900), .B0(n13901), .B1(n13902), .C0(
        n13903), .Y(n13899) );
  AOI21X1 U12228 ( .A0(n13904), .A1(n13905), .B0(n13906), .Y(n13903) );
  NAND4X1 U12229 ( .A(n13863), .B(n13912), .C(n13913), .D(n13914), .Y(n13902)
         );
  OAI221XL U12230 ( .A0(n6122), .A1(n3453), .B0(n3462), .B1(n13916), .C0(
        n13917), .Y(n13900) );
  AOI221X1 U12231 ( .A0(n2605), .A1(n18310), .B0(n18311), .B1(n18312), .C0(
        n18313), .Y(n18309) );
  AOI21X1 U12232 ( .A0(n18314), .A1(n18315), .B0(n18316), .Y(n18313) );
  NAND4X1 U12233 ( .A(n18273), .B(n18322), .C(n18323), .D(n18324), .Y(n18312)
         );
  OAI221XL U12234 ( .A0(n5000), .A1(n2610), .B0(n2617), .B1(n18326), .C0(
        n18327), .Y(n18310) );
  AOI221X1 U12235 ( .A0(n3207), .A1(n15160), .B0(n15161), .B1(n15162), .C0(
        n15163), .Y(n15159) );
  AOI21X1 U12236 ( .A0(n15164), .A1(n15165), .B0(n15166), .Y(n15163) );
  NAND4X1 U12237 ( .A(n15123), .B(n15172), .C(n15173), .D(n15174), .Y(n15162)
         );
  OAI221XL U12238 ( .A0(n5826), .A1(n3212), .B0(n3219), .B1(n15176), .C0(
        n15177), .Y(n15160) );
  AOI221X1 U12239 ( .A0(n3146), .A1(n15475), .B0(n15476), .B1(n15477), .C0(
        n15478), .Y(n15474) );
  AOI21X1 U12240 ( .A0(n15479), .A1(n15480), .B0(n15481), .Y(n15478) );
  NAND4X1 U12241 ( .A(n15438), .B(n15487), .C(n15488), .D(n15489), .Y(n15477)
         );
  OAI221XL U12242 ( .A0(n5742), .A1(n3151), .B0(n3158), .B1(n15491), .C0(
        n15492), .Y(n15475) );
  AOI221X1 U12243 ( .A0(n2544), .A1(n18625), .B0(n18626), .B1(n18627), .C0(
        n18628), .Y(n18624) );
  AOI21X1 U12244 ( .A0(n18629), .A1(n18630), .B0(n18631), .Y(n18628) );
  NAND4X1 U12245 ( .A(n18588), .B(n18637), .C(n18638), .D(n18639), .Y(n18627)
         );
  OAI221XL U12246 ( .A0(n4884), .A1(n2549), .B0(n2556), .B1(n18641), .C0(
        n18642), .Y(n18625) );
  AOI221X1 U12247 ( .A0(n2908), .A1(n16735), .B0(n16736), .B1(n16737), .C0(
        n16738), .Y(n16734) );
  AOI21X1 U12248 ( .A0(n16739), .A1(n16740), .B0(n16741), .Y(n16738) );
  NAND4X1 U12249 ( .A(n16698), .B(n16747), .C(n16748), .D(n16749), .Y(n16737)
         );
  OAI221XL U12250 ( .A0(n5438), .A1(n2913), .B0(n2920), .B1(n16751), .C0(
        n16752), .Y(n16735) );
  AOI221X1 U12251 ( .A0(n3268), .A1(n14845), .B0(n14846), .B1(n14847), .C0(
        n14848), .Y(n14844) );
  AOI21X1 U12252 ( .A0(n14849), .A1(n14850), .B0(n14851), .Y(n14848) );
  NAND4X1 U12253 ( .A(n14808), .B(n14857), .C(n14858), .D(n14859), .Y(n14847)
         );
  OAI221XL U12254 ( .A0(n5902), .A1(n3273), .B0(n3280), .B1(n14861), .C0(
        n14862), .Y(n14845) );
  AOI221X1 U12255 ( .A0(n2969), .A1(n16420), .B0(n16421), .B1(n16422), .C0(
        n16423), .Y(n16419) );
  AOI21X1 U12256 ( .A0(n16424), .A1(n16425), .B0(n16426), .Y(n16423) );
  NAND4X1 U12257 ( .A(n16383), .B(n16432), .C(n16433), .D(n16434), .Y(n16422)
         );
  OAI221XL U12258 ( .A0(n5514), .A1(n2974), .B0(n2981), .B1(n16436), .C0(
        n16437), .Y(n16420) );
  AOI221X1 U12259 ( .A0(n2666), .A1(n17995), .B0(n17996), .B1(n17997), .C0(
        n17998), .Y(n17994) );
  AOI21X1 U12260 ( .A0(n17999), .A1(n18000), .B0(n18001), .Y(n17998) );
  NAND4X1 U12261 ( .A(n17958), .B(n18007), .C(n18008), .D(n18009), .Y(n17997)
         );
  OAI221XL U12262 ( .A0(n5084), .A1(n2671), .B0(n2678), .B1(n18011), .C0(
        n18012), .Y(n17995) );
  AOI221X1 U12263 ( .A0(n3329), .A1(n14530), .B0(n14531), .B1(n14532), .C0(
        n14533), .Y(n14529) );
  AOI21X1 U12264 ( .A0(n14534), .A1(n14535), .B0(n14536), .Y(n14533) );
  NAND4X1 U12265 ( .A(n14493), .B(n14542), .C(n14543), .D(n14544), .Y(n14532)
         );
  OAI221XL U12266 ( .A0(n5978), .A1(n3334), .B0(n3341), .B1(n14546), .C0(
        n14547), .Y(n14530) );
  AOI221X1 U12267 ( .A0(n3027), .A1(n16105), .B0(n16106), .B1(n16107), .C0(
        n16108), .Y(n16104) );
  AOI21X1 U12268 ( .A0(n16109), .A1(n16110), .B0(n16111), .Y(n16108) );
  NAND4X1 U12269 ( .A(n16068), .B(n16117), .C(n16118), .D(n16119), .Y(n16107)
         );
  OAI221XL U12270 ( .A0(n5590), .A1(n3032), .B0(n3039), .B1(n16121), .C0(
        n16122), .Y(n16105) );
  AOI221X1 U12271 ( .A0(n2726), .A1(n17680), .B0(n17681), .B1(n17682), .C0(
        n17683), .Y(n17679) );
  AOI21X1 U12272 ( .A0(n17684), .A1(n17685), .B0(n17686), .Y(n17683) );
  NAND4X1 U12273 ( .A(n17643), .B(n17692), .C(n17693), .D(n17694), .Y(n17682)
         );
  OAI221XL U12274 ( .A0(n5192), .A1(n2731), .B0(n2738), .B1(n17696), .C0(
        n17697), .Y(n17680) );
  AOI221X1 U12275 ( .A0(n3387), .A1(n14215), .B0(n14216), .B1(n14217), .C0(
        n14218), .Y(n14214) );
  AOI21X1 U12276 ( .A0(n14219), .A1(n14220), .B0(n14221), .Y(n14218) );
  NAND4X1 U12277 ( .A(n14178), .B(n14227), .C(n14228), .D(n14229), .Y(n14217)
         );
  OAI221XL U12278 ( .A0(n6054), .A1(n3392), .B0(n3399), .B1(n14231), .C0(
        n14232), .Y(n14215) );
  AOI221X1 U12279 ( .A0(n3088), .A1(n15790), .B0(n15791), .B1(n15792), .C0(
        n15793), .Y(n15789) );
  AOI21X1 U12280 ( .A0(n15794), .A1(n15795), .B0(n15796), .Y(n15793) );
  NAND4X1 U12281 ( .A(n15753), .B(n15802), .C(n15803), .D(n15804), .Y(n15792)
         );
  OAI221XL U12282 ( .A0(n5666), .A1(n3093), .B0(n3100), .B1(n15806), .C0(
        n15807), .Y(n15790) );
  AOI221X1 U12283 ( .A0(n2787), .A1(n17365), .B0(n17366), .B1(n17367), .C0(
        n17368), .Y(n17364) );
  AOI21X1 U12284 ( .A0(n17369), .A1(n17370), .B0(n17371), .Y(n17368) );
  NAND4X1 U12285 ( .A(n17328), .B(n17377), .C(n17378), .D(n17379), .Y(n17367)
         );
  OAI221XL U12286 ( .A0(n5270), .A1(n2792), .B0(n2799), .B1(n17381), .C0(
        n17382), .Y(n17365) );
  AOI222X1 U12287 ( .A0(n2847), .A1(n10075), .B0(n9909), .B1(n10076), .C0(
        n5321), .C1(n10077), .Y(n10056) );
  NAND4BXL U12288 ( .AN(n10019), .B(n10074), .C(n10065), .D(n10078), .Y(n10077) );
  NAND4BXL U12289 ( .AN(n9995), .B(n9958), .C(n10079), .D(n10080), .Y(n10076)
         );
  OAI222XL U12290 ( .A0(n90), .A1(n9895), .B0(n10082), .B1(n2853), .C0(n2860), 
        .C1(n10083), .Y(n10075) );
  AOI222X1 U12291 ( .A0(n3448), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n261), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n93), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n262), .C0(n6105), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n263), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n242) );
  NAND4BXL U12292 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n205), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n260), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n251), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n264), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n263) );
  NAND4BXL U12293 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n181), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n143), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n265), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n266), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n262) );
  OAI222XL U12294 ( .A0(n91), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n78), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n268), .B1(n3454), .C0(n3460), 
        .C1(top_core_EC_ss_gen_tbox_0__sboxs_r_n269), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n261) );
  AOI222X1 U12295 ( .A0(n2605), .A1(n11243), .B0(n11077), .B1(n11244), .C0(
        n4967), .C1(n11245), .Y(n11224) );
  NAND4BXL U12296 ( .AN(n11187), .B(n11242), .C(n11233), .D(n11246), .Y(n11245) );
  NAND4BXL U12297 ( .AN(n11163), .B(n11126), .C(n11247), .D(n11248), .Y(n11244) );
  OAI222XL U12298 ( .A0(n92), .A1(n11063), .B0(n11250), .B1(n2611), .C0(n2618), 
        .C1(n11251), .Y(n11243) );
  AOI222X1 U12299 ( .A0(n3207), .A1(n8323), .B0(n8157), .B1(n8324), .C0(n5793), 
        .C1(n8325), .Y(n8304) );
  NAND4BXL U12300 ( .AN(n8267), .B(n8322), .C(n8313), .D(n8326), .Y(n8325) );
  NAND4BXL U12301 ( .AN(n8243), .B(n8206), .C(n8327), .D(n8328), .Y(n8324) );
  OAI222XL U12302 ( .A0(n93), .A1(n8143), .B0(n8330), .B1(n3213), .C0(n3220), 
        .C1(n8331), .Y(n8323) );
  AOI222X1 U12303 ( .A0(n2666), .A1(n10951), .B0(n10785), .B1(n10952), .C0(
        n5051), .C1(n10953), .Y(n10932) );
  NAND4BXL U12304 ( .AN(n10895), .B(n10950), .C(n10941), .D(n10954), .Y(n10953) );
  NAND4BXL U12305 ( .AN(n10871), .B(n10834), .C(n10955), .D(n10956), .Y(n10952) );
  OAI222XL U12306 ( .A0(n94), .A1(n10771), .B0(n10958), .B1(n2672), .C0(n2679), 
        .C1(n10959), .Y(n10951) );
  AOI222X1 U12307 ( .A0(n3387), .A1(n7447), .B0(n7281), .B1(n7448), .C0(n6021), 
        .C1(n7449), .Y(n7428) );
  NAND4BXL U12308 ( .AN(n7391), .B(n7446), .C(n7437), .D(n7450), .Y(n7449) );
  NAND4BXL U12309 ( .AN(n7367), .B(n7330), .C(n7451), .D(n7452), .Y(n7448) );
  OAI222XL U12310 ( .A0(n95), .A1(n7267), .B0(n7454), .B1(n3393), .C0(n3400), 
        .C1(n7455), .Y(n7447) );
  AOI222X1 U12311 ( .A0(n3027), .A1(n9199), .B0(n9033), .B1(n9200), .C0(n5557), 
        .C1(n9201), .Y(n9180) );
  NAND4BXL U12312 ( .AN(n9143), .B(n9198), .C(n9189), .D(n9202), .Y(n9201) );
  NAND4BXL U12313 ( .AN(n9119), .B(n9082), .C(n9203), .D(n9204), .Y(n9200) );
  OAI222XL U12314 ( .A0(n96), .A1(n9019), .B0(n9206), .B1(n3033), .C0(n3040), 
        .C1(n9207), .Y(n9199) );
  AOI222X1 U12315 ( .A0(n2787), .A1(n10367), .B0(n10201), .B1(n10368), .C0(
        n5237), .C1(n10369), .Y(n10348) );
  NAND4BXL U12316 ( .AN(n10311), .B(n10366), .C(n10357), .D(n10370), .Y(n10369) );
  NAND4BXL U12317 ( .AN(n10287), .B(n10250), .C(n10371), .D(n10372), .Y(n10368) );
  OAI222XL U12318 ( .A0(n97), .A1(n10187), .B0(n10374), .B1(n2793), .C0(n2800), 
        .C1(n10375), .Y(n10367) );
  AOI222X1 U12319 ( .A0(n2969), .A1(n9491), .B0(n9325), .B1(n9492), .C0(n5481), 
        .C1(n9493), .Y(n9472) );
  NAND4BXL U12320 ( .AN(n9435), .B(n9490), .C(n9481), .D(n9494), .Y(n9493) );
  NAND4BXL U12321 ( .AN(n9411), .B(n9374), .C(n9495), .D(n9496), .Y(n9492) );
  OAI222XL U12322 ( .A0(n98), .A1(n9311), .B0(n9498), .B1(n2975), .C0(n2982), 
        .C1(n9499), .Y(n9491) );
  AOI222X1 U12323 ( .A0(n3146), .A1(n8615), .B0(n8449), .B1(n8616), .C0(n5709), 
        .C1(n8617), .Y(n8596) );
  NAND4BXL U12324 ( .AN(n8559), .B(n8614), .C(n8605), .D(n8618), .Y(n8617) );
  NAND4BXL U12325 ( .AN(n8535), .B(n8498), .C(n8619), .D(n8620), .Y(n8616) );
  OAI222XL U12326 ( .A0(n99), .A1(n8435), .B0(n8622), .B1(n3152), .C0(n3159), 
        .C1(n8623), .Y(n8615) );
  AOI222X1 U12327 ( .A0(n3329), .A1(n7739), .B0(n7573), .B1(n7740), .C0(n5945), 
        .C1(n7741), .Y(n7720) );
  NAND4BXL U12328 ( .AN(n7683), .B(n7738), .C(n7729), .D(n7742), .Y(n7741) );
  NAND4BXL U12329 ( .AN(n7659), .B(n7622), .C(n7743), .D(n7744), .Y(n7740) );
  OAI222XL U12330 ( .A0(n100), .A1(n7559), .B0(n7746), .B1(n3335), .C0(n3342), 
        .C1(n7747), .Y(n7739) );
  AOI222X1 U12331 ( .A0(n2544), .A1(n11535), .B0(n11369), .B1(n11536), .C0(
        n4851), .C1(n11537), .Y(n11516) );
  NAND4BXL U12332 ( .AN(n11479), .B(n11534), .C(n11525), .D(n11538), .Y(n11537) );
  NAND4BXL U12333 ( .AN(n11455), .B(n11418), .C(n11539), .D(n11540), .Y(n11536) );
  OAI222XL U12334 ( .A0(n101), .A1(n11355), .B0(n11542), .B1(n2550), .C0(n2557), .C1(n11543), .Y(n11535) );
  AOI222X1 U12335 ( .A0(n2726), .A1(n10659), .B0(n10493), .B1(n10660), .C0(
        n5159), .C1(n10661), .Y(n10640) );
  NAND4BXL U12336 ( .AN(n10603), .B(n10658), .C(n10649), .D(n10662), .Y(n10661) );
  NAND4BXL U12337 ( .AN(n10579), .B(n10542), .C(n10663), .D(n10664), .Y(n10660) );
  OAI222XL U12338 ( .A0(n102), .A1(n10479), .B0(n10666), .B1(n2732), .C0(n2739), .C1(n10667), .Y(n10659) );
  AOI222X1 U12339 ( .A0(n2908), .A1(n9783), .B0(n9617), .B1(n9784), .C0(n5405), 
        .C1(n9785), .Y(n9764) );
  NAND4BXL U12340 ( .AN(n9727), .B(n9782), .C(n9773), .D(n9786), .Y(n9785) );
  NAND4BXL U12341 ( .AN(n9703), .B(n9666), .C(n9787), .D(n9788), .Y(n9784) );
  OAI222XL U12342 ( .A0(n103), .A1(n9603), .B0(n9790), .B1(n2914), .C0(n2921), 
        .C1(n9791), .Y(n9783) );
  AOI222X1 U12343 ( .A0(n3088), .A1(n8907), .B0(n8741), .B1(n8908), .C0(n5633), 
        .C1(n8909), .Y(n8888) );
  NAND4BXL U12344 ( .AN(n8851), .B(n8906), .C(n8897), .D(n8910), .Y(n8909) );
  NAND4BXL U12345 ( .AN(n8827), .B(n8790), .C(n8911), .D(n8912), .Y(n8908) );
  OAI222XL U12346 ( .A0(n104), .A1(n8727), .B0(n8914), .B1(n3094), .C0(n3101), 
        .C1(n8915), .Y(n8907) );
  AOI222X1 U12347 ( .A0(n3268), .A1(n8031), .B0(n7865), .B1(n8032), .C0(n5869), 
        .C1(n8033), .Y(n8012) );
  NAND4BXL U12348 ( .AN(n7975), .B(n8030), .C(n8021), .D(n8034), .Y(n8033) );
  NAND4BXL U12349 ( .AN(n7951), .B(n7914), .C(n8035), .D(n8036), .Y(n8032) );
  OAI222XL U12350 ( .A0(n105), .A1(n7851), .B0(n8038), .B1(n3274), .C0(n3281), 
        .C1(n8039), .Y(n8031) );
  AOI211X1 U12351 ( .A0(n5380), .A1(n2890), .B0(n17221), .C0(n17222), .Y(
        n17216) );
  OAI21XL U12352 ( .A0(n17223), .A1(n17047), .B0(n17224), .Y(n17222) );
  AOI211X1 U12353 ( .A0(n6151), .A1(n3488), .B0(n14071), .C0(n14072), .Y(
        n14066) );
  OAI21XL U12354 ( .A0(n14073), .A1(n13897), .B0(n14074), .Y(n14072) );
  AOI211X1 U12355 ( .A0(n5852), .A1(n3247), .B0(n15331), .C0(n15332), .Y(
        n15326) );
  OAI21XL U12356 ( .A0(n15333), .A1(n15157), .B0(n15334), .Y(n15332) );
  AOI211X1 U12357 ( .A0(n5026), .A1(n2645), .B0(n18481), .C0(n18482), .Y(
        n18476) );
  OAI21XL U12358 ( .A0(n18483), .A1(n18307), .B0(n18484), .Y(n18482) );
  AOI211X1 U12359 ( .A0(n5768), .A1(n3187), .B0(n15646), .C0(n15647), .Y(
        n15641) );
  OAI21XL U12360 ( .A0(n15648), .A1(n15472), .B0(n15649), .Y(n15647) );
  AOI211X1 U12361 ( .A0(n5464), .A1(n2948), .B0(n16906), .C0(n16907), .Y(
        n16901) );
  OAI21XL U12362 ( .A0(n16908), .A1(n16732), .B0(n16909), .Y(n16907) );
  AOI211X1 U12363 ( .A0(n4910), .A1(n2585), .B0(n18796), .C0(n18797), .Y(
        n18791) );
  OAI21XL U12364 ( .A0(n18798), .A1(n18622), .B0(n18799), .Y(n18797) );
  AOI211X1 U12365 ( .A0(n5928), .A1(n3308), .B0(n15016), .C0(n15017), .Y(
        n15011) );
  OAI21XL U12366 ( .A0(n15018), .A1(n14842), .B0(n15019), .Y(n15017) );
  AOI211X1 U12367 ( .A0(n5540), .A1(n3009), .B0(n16591), .C0(n16592), .Y(
        n16586) );
  OAI21XL U12368 ( .A0(n16593), .A1(n16417), .B0(n16594), .Y(n16592) );
  AOI211X1 U12369 ( .A0(n5110), .A1(n2707), .B0(n18166), .C0(n18167), .Y(
        n18161) );
  OAI21XL U12370 ( .A0(n18168), .A1(n17992), .B0(n18169), .Y(n18167) );
  AOI211X1 U12371 ( .A0(n6004), .A1(n3370), .B0(n14701), .C0(n14702), .Y(
        n14696) );
  OAI21XL U12372 ( .A0(n14703), .A1(n14527), .B0(n14704), .Y(n14702) );
  AOI211X1 U12373 ( .A0(n5616), .A1(n3067), .B0(n16276), .C0(n16277), .Y(
        n16271) );
  OAI21XL U12374 ( .A0(n16278), .A1(n16102), .B0(n16279), .Y(n16277) );
  AOI211X1 U12375 ( .A0(n5218), .A1(n2767), .B0(n17851), .C0(n17852), .Y(
        n17846) );
  OAI21XL U12376 ( .A0(n17853), .A1(n17677), .B0(n17854), .Y(n17852) );
  AOI211X1 U12377 ( .A0(n6080), .A1(n3427), .B0(n14386), .C0(n14387), .Y(
        n14381) );
  OAI21XL U12378 ( .A0(n14388), .A1(n14212), .B0(n14389), .Y(n14387) );
  AOI211X1 U12379 ( .A0(n5692), .A1(n3129), .B0(n15961), .C0(n15962), .Y(
        n15956) );
  OAI21XL U12380 ( .A0(n15963), .A1(n15787), .B0(n15964), .Y(n15962) );
  AOI211X1 U12381 ( .A0(n5296), .A1(n2827), .B0(n17536), .C0(n17537), .Y(
        n17531) );
  OAI21XL U12382 ( .A0(n17538), .A1(n17362), .B0(n17539), .Y(n17537) );
  AOI222X1 U12383 ( .A0(n10058), .A1(n2850), .B0(n5322), .B1(n10059), .C0(
        n5325), .C1(n10060), .Y(n10057) );
  NAND3X1 U12384 ( .A(n10061), .B(n10062), .C(n10063), .Y(n10060) );
  AOI222X1 U12385 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n244), .A1(n3451), 
        .B0(n6109), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n245), .C0(n6107), 
        .C1(top_core_EC_ss_gen_tbox_0__sboxs_r_n246), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n243) );
  NAND3X1 U12386 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n247), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n248), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n249), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n246) );
  AOI222X1 U12387 ( .A0(n11226), .A1(n2608), .B0(n4968), .B1(n11227), .C0(
        n4971), .C1(n11228), .Y(n11225) );
  NAND3X1 U12388 ( .A(n11229), .B(n11230), .C(n11231), .Y(n11228) );
  AOI222X1 U12389 ( .A0(n8306), .A1(n3210), .B0(n5794), .B1(n8307), .C0(n5797), 
        .C1(n8308), .Y(n8305) );
  NAND3X1 U12390 ( .A(n8309), .B(n8310), .C(n8311), .Y(n8308) );
  AOI222X1 U12391 ( .A0(n10934), .A1(n2669), .B0(n5052), .B1(n10935), .C0(
        n5055), .C1(n10936), .Y(n10933) );
  NAND3X1 U12392 ( .A(n10937), .B(n10938), .C(n10939), .Y(n10936) );
  AOI222X1 U12393 ( .A0(n7430), .A1(n3390), .B0(n6022), .B1(n7431), .C0(n6025), 
        .C1(n7432), .Y(n7429) );
  NAND3X1 U12394 ( .A(n7433), .B(n7434), .C(n7435), .Y(n7432) );
  AOI222X1 U12395 ( .A0(n9182), .A1(n3030), .B0(n5558), .B1(n9183), .C0(n5561), 
        .C1(n9184), .Y(n9181) );
  NAND3X1 U12396 ( .A(n9185), .B(n9186), .C(n9187), .Y(n9184) );
  AOI222X1 U12397 ( .A0(n10350), .A1(n2790), .B0(n5238), .B1(n10351), .C0(
        n5241), .C1(n10352), .Y(n10349) );
  NAND3X1 U12398 ( .A(n10353), .B(n10354), .C(n10355), .Y(n10352) );
  AOI222X1 U12399 ( .A0(n9474), .A1(n2972), .B0(n5482), .B1(n9475), .C0(n5485), 
        .C1(n9476), .Y(n9473) );
  NAND3X1 U12400 ( .A(n9477), .B(n9478), .C(n9479), .Y(n9476) );
  AOI222X1 U12401 ( .A0(n8598), .A1(n3149), .B0(n5710), .B1(n8599), .C0(n5713), 
        .C1(n8600), .Y(n8597) );
  NAND3X1 U12402 ( .A(n8601), .B(n8602), .C(n8603), .Y(n8600) );
  AOI222X1 U12403 ( .A0(n7722), .A1(n3332), .B0(n5946), .B1(n7723), .C0(n5949), 
        .C1(n7724), .Y(n7721) );
  NAND3X1 U12404 ( .A(n7725), .B(n7726), .C(n7727), .Y(n7724) );
  AOI222X1 U12405 ( .A0(n11518), .A1(n2547), .B0(n4852), .B1(n11519), .C0(
        n4855), .C1(n11520), .Y(n11517) );
  NAND3X1 U12406 ( .A(n11521), .B(n11522), .C(n11523), .Y(n11520) );
  AOI222X1 U12407 ( .A0(n10642), .A1(n2729), .B0(n5160), .B1(n10643), .C0(
        n5163), .C1(n10644), .Y(n10641) );
  NAND3X1 U12408 ( .A(n10645), .B(n10646), .C(n10647), .Y(n10644) );
  AOI222X1 U12409 ( .A0(n9766), .A1(n2911), .B0(n5406), .B1(n9767), .C0(n5409), 
        .C1(n9768), .Y(n9765) );
  NAND3X1 U12410 ( .A(n9769), .B(n9770), .C(n9771), .Y(n9768) );
  AOI222X1 U12411 ( .A0(n8890), .A1(n3091), .B0(n5634), .B1(n8891), .C0(n5637), 
        .C1(n8892), .Y(n8889) );
  NAND3X1 U12412 ( .A(n8893), .B(n8894), .C(n8895), .Y(n8892) );
  AOI222X1 U12413 ( .A0(n8014), .A1(n3271), .B0(n5870), .B1(n8015), .C0(n5873), 
        .C1(n8016), .Y(n8013) );
  NAND3X1 U12414 ( .A(n8017), .B(n8018), .C(n8019), .Y(n8016) );
  AOI211X1 U12415 ( .A0(n2867), .A1(n2902), .B0(n9997), .C0(n9964), .Y(n9989)
         );
  OAI221XL U12416 ( .A0(n2881), .A1(n9998), .B0(n1004), .B1(n9893), .C0(n9999), 
        .Y(n9997) );
  AOI211X1 U12417 ( .A0(n3468), .A1(top_core_EC_ss_in[0]), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n183), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n149), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n175) );
  OAI221XL U12418 ( .A0(n3483), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n184), 
        .B0(n1145), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n76), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n185), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n183) );
  AOI211X1 U12419 ( .A0(n2625), .A1(n2651), .B0(n11165), .C0(n11132), .Y(
        n11157) );
  OAI221XL U12420 ( .A0(n2639), .A1(n11166), .B0(n948), .B1(n11061), .C0(
        n11167), .Y(n11165) );
  AOI211X1 U12421 ( .A0(n3227), .A1(n3262), .B0(n8245), .C0(n8212), .Y(n8237)
         );
  OAI221XL U12422 ( .A0(n3241), .A1(n8246), .B0(n1088), .B1(n8141), .C0(n8247), 
        .Y(n8245) );
  AOI211X1 U12423 ( .A0(n2686), .A1(top_core_EC_ss_in[104]), .B0(n10873), .C0(
        n10840), .Y(n10865) );
  OAI221XL U12424 ( .A0(n2700), .A1(n10874), .B0(n962), .B1(n10769), .C0(
        n10875), .Y(n10873) );
  AOI211X1 U12425 ( .A0(n3047), .A1(n3073), .B0(n9121), .C0(n9088), .Y(n9113)
         );
  OAI221XL U12426 ( .A0(n3061), .A1(n9122), .B0(n1046), .B1(n9017), .C0(n9123), 
        .Y(n9121) );
  AOI211X1 U12427 ( .A0(n3407), .A1(top_core_EC_ss_in[8]), .B0(n7369), .C0(
        n7336), .Y(n7361) );
  OAI221XL U12428 ( .A0(n3421), .A1(n7370), .B0(n1130), .B1(n7265), .C0(n7371), 
        .Y(n7369) );
  AOI211X1 U12429 ( .A0(n2807), .A1(n2834), .B0(n10289), .C0(n10256), .Y(
        n10281) );
  OAI221XL U12430 ( .A0(n2821), .A1(n10290), .B0(n990), .B1(n10185), .C0(
        n10291), .Y(n10289) );
  AOI211X1 U12431 ( .A0(n2989), .A1(n3016), .B0(n9413), .C0(n9380), .Y(n9405)
         );
  OAI221XL U12432 ( .A0(n3003), .A1(n9414), .B0(n1032), .B1(n9309), .C0(n9415), 
        .Y(n9413) );
  AOI211X1 U12433 ( .A0(n3166), .A1(n3201), .B0(n8537), .C0(n8504), .Y(n8529)
         );
  OAI221XL U12434 ( .A0(n3180), .A1(n8538), .B0(n1074), .B1(n8433), .C0(n8539), 
        .Y(n8537) );
  AOI211X1 U12435 ( .A0(n3349), .A1(n3376), .B0(n7661), .C0(n7628), .Y(n7653)
         );
  OAI221XL U12436 ( .A0(n3363), .A1(n7662), .B0(n1116), .B1(n7557), .C0(n7663), 
        .Y(n7661) );
  AOI211X1 U12437 ( .A0(n2564), .A1(n2590), .B0(n11457), .C0(n11424), .Y(
        n11449) );
  OAI221XL U12438 ( .A0(n2578), .A1(n11458), .B0(n934), .B1(n11353), .C0(
        n11459), .Y(n11457) );
  AOI211X1 U12439 ( .A0(n2746), .A1(n2773), .B0(n10581), .C0(n10548), .Y(
        n10573) );
  OAI221XL U12440 ( .A0(n2760), .A1(n10582), .B0(n976), .B1(n10477), .C0(
        n10583), .Y(n10581) );
  AOI211X1 U12441 ( .A0(n2928), .A1(n2963), .B0(n9705), .C0(n9672), .Y(n9697)
         );
  OAI221XL U12442 ( .A0(n2942), .A1(n9706), .B0(n1018), .B1(n9601), .C0(n9707), 
        .Y(n9705) );
  AOI211X1 U12443 ( .A0(n3108), .A1(n3135), .B0(n8829), .C0(n8796), .Y(n8821)
         );
  OAI221XL U12444 ( .A0(n3122), .A1(n8830), .B0(n1060), .B1(n8725), .C0(n8831), 
        .Y(n8829) );
  AOI211X1 U12445 ( .A0(n3288), .A1(n3324), .B0(n7953), .C0(n7920), .Y(n7945)
         );
  OAI221XL U12446 ( .A0(n3302), .A1(n7954), .B0(n1102), .B1(n7849), .C0(n7955), 
        .Y(n7953) );
  INVX1 U12447 ( .A(n13333), .Y(n6546) );
  INVX1 U12448 ( .A(n12703), .Y(n6841) );
  INVX1 U12449 ( .A(n13648), .Y(n6594) );
  INVX1 U12450 ( .A(n13018), .Y(n6887) );
  AOI221X1 U12451 ( .A0(n17051), .A1(n17213), .B0(n5326), .B1(n17214), .C0(
        n17215), .Y(n17212) );
  NAND4BXL U12452 ( .AN(n17059), .B(n17091), .C(n17226), .D(n17227), .Y(n17213) );
  NAND4X1 U12453 ( .A(n17091), .B(n17143), .C(n17013), .D(n17225), .Y(n17214)
         );
  OAI2BB2X1 U12454 ( .B0(n17216), .B1(n17087), .A0N(n17217), .A1N(n5321), .Y(
        n17215) );
  AOI221X1 U12455 ( .A0(n13901), .A1(n14063), .B0(n6108), .B1(n14064), .C0(
        n14065), .Y(n14062) );
  NAND4BXL U12456 ( .AN(n13909), .B(n13941), .C(n14076), .D(n14077), .Y(n14063) );
  NAND4X1 U12457 ( .A(n13941), .B(n13993), .C(n13863), .D(n14075), .Y(n14064)
         );
  OAI2BB2X1 U12458 ( .B0(n14066), .B1(n13937), .A0N(n14067), .A1N(n6105), .Y(
        n14065) );
  AOI221X1 U12459 ( .A0(n15161), .A1(n15323), .B0(n5798), .B1(n15324), .C0(
        n15325), .Y(n15322) );
  NAND4BXL U12460 ( .AN(n15169), .B(n15201), .C(n15336), .D(n15337), .Y(n15323) );
  NAND4X1 U12461 ( .A(n15201), .B(n15253), .C(n15123), .D(n15335), .Y(n15324)
         );
  OAI2BB2X1 U12462 ( .B0(n15326), .B1(n15197), .A0N(n15327), .A1N(n5793), .Y(
        n15325) );
  AOI221X1 U12463 ( .A0(n18311), .A1(n18473), .B0(n4972), .B1(n18474), .C0(
        n18475), .Y(n18472) );
  NAND4BXL U12464 ( .AN(n18319), .B(n18351), .C(n18486), .D(n18487), .Y(n18473) );
  NAND4X1 U12465 ( .A(n18351), .B(n18403), .C(n18273), .D(n18485), .Y(n18474)
         );
  OAI2BB2X1 U12466 ( .B0(n18476), .B1(n18347), .A0N(n18477), .A1N(n4967), .Y(
        n18475) );
  AOI221X1 U12467 ( .A0(n15476), .A1(n15638), .B0(n5714), .B1(n15639), .C0(
        n15640), .Y(n15637) );
  NAND4BXL U12468 ( .AN(n15484), .B(n15516), .C(n15651), .D(n15652), .Y(n15638) );
  NAND4X1 U12469 ( .A(n15516), .B(n15568), .C(n15438), .D(n15650), .Y(n15639)
         );
  OAI2BB2X1 U12470 ( .B0(n15641), .B1(n15512), .A0N(n15642), .A1N(n5709), .Y(
        n15640) );
  AOI221X1 U12471 ( .A0(n16736), .A1(n16898), .B0(n5410), .B1(n16899), .C0(
        n16900), .Y(n16897) );
  NAND4BXL U12472 ( .AN(n16744), .B(n16776), .C(n16911), .D(n16912), .Y(n16898) );
  NAND4X1 U12473 ( .A(n16776), .B(n16828), .C(n16698), .D(n16910), .Y(n16899)
         );
  OAI2BB2X1 U12474 ( .B0(n16901), .B1(n16772), .A0N(n16902), .A1N(n5405), .Y(
        n16900) );
  AOI221X1 U12475 ( .A0(n18626), .A1(n18788), .B0(n4856), .B1(n18789), .C0(
        n18790), .Y(n18787) );
  NAND4BXL U12476 ( .AN(n18634), .B(n18666), .C(n18801), .D(n18802), .Y(n18788) );
  NAND4X1 U12477 ( .A(n18666), .B(n18718), .C(n18588), .D(n18800), .Y(n18789)
         );
  OAI2BB2X1 U12478 ( .B0(n18791), .B1(n18662), .A0N(n18792), .A1N(n4851), .Y(
        n18790) );
  AOI221X1 U12479 ( .A0(n14846), .A1(n15008), .B0(n5874), .B1(n15009), .C0(
        n15010), .Y(n15007) );
  NAND4BXL U12480 ( .AN(n14854), .B(n14886), .C(n15021), .D(n15022), .Y(n15008) );
  NAND4X1 U12481 ( .A(n14886), .B(n14938), .C(n14808), .D(n15020), .Y(n15009)
         );
  OAI2BB2X1 U12482 ( .B0(n15011), .B1(n14882), .A0N(n15012), .A1N(n5869), .Y(
        n15010) );
  AOI221X1 U12483 ( .A0(n16421), .A1(n16583), .B0(n5486), .B1(n16584), .C0(
        n16585), .Y(n16582) );
  NAND4BXL U12484 ( .AN(n16429), .B(n16461), .C(n16596), .D(n16597), .Y(n16583) );
  NAND4X1 U12485 ( .A(n16461), .B(n16513), .C(n16383), .D(n16595), .Y(n16584)
         );
  OAI2BB2X1 U12486 ( .B0(n16586), .B1(n16457), .A0N(n16587), .A1N(n5481), .Y(
        n16585) );
  AOI221X1 U12487 ( .A0(n17996), .A1(n18158), .B0(n5056), .B1(n18159), .C0(
        n18160), .Y(n18157) );
  NAND4BXL U12488 ( .AN(n18004), .B(n18036), .C(n18171), .D(n18172), .Y(n18158) );
  NAND4X1 U12489 ( .A(n18036), .B(n18088), .C(n17958), .D(n18170), .Y(n18159)
         );
  OAI2BB2X1 U12490 ( .B0(n18161), .B1(n18032), .A0N(n18162), .A1N(n5051), .Y(
        n18160) );
  AOI221X1 U12491 ( .A0(n14531), .A1(n14693), .B0(n5950), .B1(n14694), .C0(
        n14695), .Y(n14692) );
  NAND4BXL U12492 ( .AN(n14539), .B(n14571), .C(n14706), .D(n14707), .Y(n14693) );
  NAND4X1 U12493 ( .A(n14571), .B(n14623), .C(n14493), .D(n14705), .Y(n14694)
         );
  OAI2BB2X1 U12494 ( .B0(n14696), .B1(n14567), .A0N(n14697), .A1N(n5945), .Y(
        n14695) );
  AOI221X1 U12495 ( .A0(n16106), .A1(n16268), .B0(n5562), .B1(n16269), .C0(
        n16270), .Y(n16267) );
  NAND4BXL U12496 ( .AN(n16114), .B(n16146), .C(n16281), .D(n16282), .Y(n16268) );
  NAND4X1 U12497 ( .A(n16146), .B(n16198), .C(n16068), .D(n16280), .Y(n16269)
         );
  OAI2BB2X1 U12498 ( .B0(n16271), .B1(n16142), .A0N(n16272), .A1N(n5557), .Y(
        n16270) );
  AOI221X1 U12499 ( .A0(n17681), .A1(n17843), .B0(n5164), .B1(n17844), .C0(
        n17845), .Y(n17842) );
  NAND4BXL U12500 ( .AN(n17689), .B(n17721), .C(n17856), .D(n17857), .Y(n17843) );
  NAND4X1 U12501 ( .A(n17721), .B(n17773), .C(n17643), .D(n17855), .Y(n17844)
         );
  OAI2BB2X1 U12502 ( .B0(n17846), .B1(n17717), .A0N(n17847), .A1N(n5159), .Y(
        n17845) );
  AOI221X1 U12503 ( .A0(n14216), .A1(n14378), .B0(n6026), .B1(n14379), .C0(
        n14380), .Y(n14377) );
  NAND4BXL U12504 ( .AN(n14224), .B(n14256), .C(n14391), .D(n14392), .Y(n14378) );
  NAND4X1 U12505 ( .A(n14256), .B(n14308), .C(n14178), .D(n14390), .Y(n14379)
         );
  OAI2BB2X1 U12506 ( .B0(n14381), .B1(n14252), .A0N(n14382), .A1N(n6021), .Y(
        n14380) );
  AOI221X1 U12507 ( .A0(n15791), .A1(n15953), .B0(n5638), .B1(n15954), .C0(
        n15955), .Y(n15952) );
  NAND4BXL U12508 ( .AN(n15799), .B(n15831), .C(n15966), .D(n15967), .Y(n15953) );
  NAND4X1 U12509 ( .A(n15831), .B(n15883), .C(n15753), .D(n15965), .Y(n15954)
         );
  OAI2BB2X1 U12510 ( .B0(n15956), .B1(n15827), .A0N(n15957), .A1N(n5633), .Y(
        n15955) );
  AOI221X1 U12511 ( .A0(n17366), .A1(n17528), .B0(n5242), .B1(n17529), .C0(
        n17530), .Y(n17527) );
  NAND4BXL U12512 ( .AN(n17374), .B(n17406), .C(n17541), .D(n17542), .Y(n17528) );
  NAND4X1 U12513 ( .A(n17406), .B(n17458), .C(n17328), .D(n17540), .Y(n17529)
         );
  OAI2BB2X1 U12514 ( .B0(n17531), .B1(n17402), .A0N(n17532), .A1N(n5237), .Y(
        n17530) );
  AOI221X1 U12515 ( .A0(n722), .A1(n5333), .B0(n5348), .B1(n5392), .C0(n10016), 
        .Y(n9977) );
  OAI211X1 U12516 ( .A0(n2858), .A1(n10017), .B0(n10018), .C0(n9974), .Y(
        n10016) );
  OAI21XL U12517 ( .A0(n10019), .A1(n5369), .B0(n2860), .Y(n10018) );
  AOI221X1 U12518 ( .A0(n723), .A1(n6119), .B0(n6144), .B1(n6176), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n202), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n163) );
  OAI211X1 U12519 ( .A0(n3459), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n203), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n204), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n160), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n202) );
  OAI21XL U12520 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n205), .A1(n6159), 
        .B0(n3456), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n204) );
  AOI221X1 U12521 ( .A0(n724), .A1(n4979), .B0(n4994), .B1(n5038), .C0(n11184), 
        .Y(n11145) );
  OAI211X1 U12522 ( .A0(n2616), .A1(n11185), .B0(n11186), .C0(n11142), .Y(
        n11184) );
  OAI21XL U12523 ( .A0(n11187), .A1(n5015), .B0(n2617), .Y(n11186) );
  AOI221X1 U12524 ( .A0(n725), .A1(n5805), .B0(n5820), .B1(n5864), .C0(n8264), 
        .Y(n8225) );
  OAI211X1 U12525 ( .A0(n3218), .A1(n8265), .B0(n8266), .C0(n8222), .Y(n8264)
         );
  OAI21XL U12526 ( .A0(n8267), .A1(n5841), .B0(n3220), .Y(n8266) );
  AOI221X1 U12527 ( .A0(n731), .A1(n5063), .B0(n5078), .B1(n5122), .C0(n10892), 
        .Y(n10853) );
  OAI211X1 U12528 ( .A0(n2677), .A1(n10893), .B0(n10894), .C0(n10850), .Y(
        n10892) );
  OAI21XL U12529 ( .A0(n10895), .A1(n5099), .B0(n2679), .Y(n10894) );
  AOI221X1 U12530 ( .A0(n733), .A1(n5569), .B0(n5584), .B1(n5628), .C0(n9140), 
        .Y(n9101) );
  OAI211X1 U12531 ( .A0(n3038), .A1(n9141), .B0(n9142), .C0(n9098), .Y(n9140)
         );
  OAI21XL U12532 ( .A0(n9143), .A1(n5605), .B0(n3039), .Y(n9142) );
  AOI221X1 U12533 ( .A0(n735), .A1(n6033), .B0(n6048), .B1(n6092), .C0(n7388), 
        .Y(n7349) );
  OAI211X1 U12534 ( .A0(n3398), .A1(n7389), .B0(n7390), .C0(n7346), .Y(n7388)
         );
  OAI21XL U12535 ( .A0(n7391), .A1(n6069), .B0(n3399), .Y(n7390) );
  AOI221X1 U12536 ( .A0(n737), .A1(n5249), .B0(n5264), .B1(n5308), .C0(n10308), 
        .Y(n10269) );
  OAI211X1 U12537 ( .A0(n2798), .A1(n10309), .B0(n10310), .C0(n10266), .Y(
        n10308) );
  OAI21XL U12538 ( .A0(n10311), .A1(n5285), .B0(n2799), .Y(n10310) );
  AOI221X1 U12539 ( .A0(n730), .A1(n5493), .B0(n5508), .B1(n5552), .C0(n9432), 
        .Y(n9393) );
  OAI211X1 U12540 ( .A0(n2980), .A1(n9433), .B0(n9434), .C0(n9390), .Y(n9432)
         );
  OAI21XL U12541 ( .A0(n9435), .A1(n5529), .B0(n2981), .Y(n9434) );
  AOI221X1 U12542 ( .A0(n726), .A1(n5721), .B0(n5736), .B1(n5780), .C0(n8556), 
        .Y(n8517) );
  OAI211X1 U12543 ( .A0(n3157), .A1(n8557), .B0(n8558), .C0(n8514), .Y(n8556)
         );
  OAI21XL U12544 ( .A0(n8559), .A1(n5757), .B0(n3158), .Y(n8558) );
  AOI221X1 U12545 ( .A0(n732), .A1(n5957), .B0(n5972), .B1(n6016), .C0(n7680), 
        .Y(n7641) );
  OAI211X1 U12546 ( .A0(n3340), .A1(n7681), .B0(n7682), .C0(n7638), .Y(n7680)
         );
  OAI21XL U12547 ( .A0(n7683), .A1(n5993), .B0(n3341), .Y(n7682) );
  AOI221X1 U12548 ( .A0(n728), .A1(n4863), .B0(n4878), .B1(n4922), .C0(n11476), 
        .Y(n11437) );
  OAI211X1 U12549 ( .A0(n2555), .A1(n11477), .B0(n11478), .C0(n11434), .Y(
        n11476) );
  OAI21XL U12550 ( .A0(n11479), .A1(n4899), .B0(n2559), .Y(n11478) );
  AOI221X1 U12551 ( .A0(n734), .A1(n5171), .B0(n5186), .B1(n5230), .C0(n10600), 
        .Y(n10561) );
  OAI211X1 U12552 ( .A0(n2737), .A1(n10601), .B0(n10602), .C0(n10558), .Y(
        n10600) );
  OAI21XL U12553 ( .A0(n10603), .A1(n5207), .B0(n2739), .Y(n10602) );
  AOI221X1 U12554 ( .A0(n727), .A1(n5417), .B0(n5432), .B1(n5476), .C0(n9724), 
        .Y(n9685) );
  OAI211X1 U12555 ( .A0(n2919), .A1(n9725), .B0(n9726), .C0(n9682), .Y(n9724)
         );
  OAI21XL U12556 ( .A0(n9727), .A1(n5453), .B0(n2920), .Y(n9726) );
  AOI221X1 U12557 ( .A0(n736), .A1(n5645), .B0(n5660), .B1(n5704), .C0(n8848), 
        .Y(n8809) );
  OAI211X1 U12558 ( .A0(n3099), .A1(n8849), .B0(n8850), .C0(n8806), .Y(n8848)
         );
  OAI21XL U12559 ( .A0(n8851), .A1(n5681), .B0(n3101), .Y(n8850) );
  AOI221X1 U12560 ( .A0(n729), .A1(n5881), .B0(n5896), .B1(n5940), .C0(n7972), 
        .Y(n7933) );
  OAI211X1 U12561 ( .A0(n3279), .A1(n7973), .B0(n7974), .C0(n7930), .Y(n7972)
         );
  OAI21XL U12562 ( .A0(n7975), .A1(n5917), .B0(n3280), .Y(n7974) );
  AOI221X1 U12563 ( .A0(n9909), .A1(n10025), .B0(n5321), .B1(n10026), .C0(
        n10027), .Y(n10024) );
  NAND4BXL U12564 ( .AN(n10035), .B(n9950), .C(n10036), .D(n10037), .Y(n10026)
         );
  OAI22X1 U12565 ( .A0(n10028), .A1(n9990), .B0(n10029), .B1(n9992), .Y(n10027) );
  AOI221X1 U12566 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n93), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n211), .B0(n6105), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n212), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n213), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n210) );
  NAND4BXL U12567 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n221), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n135), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n222), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n223), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n212) );
  OAI22X1 U12568 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n214), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n176), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n215), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n178), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n213) );
  AOI221X1 U12569 ( .A0(n11077), .A1(n11193), .B0(n4967), .B1(n11194), .C0(
        n11195), .Y(n11192) );
  NAND4BXL U12570 ( .AN(n11203), .B(n11118), .C(n11204), .D(n11205), .Y(n11194) );
  OAI22X1 U12571 ( .A0(n11196), .A1(n11158), .B0(n11197), .B1(n11160), .Y(
        n11195) );
  AOI221X1 U12572 ( .A0(n8157), .A1(n8273), .B0(n5793), .B1(n8274), .C0(n8275), 
        .Y(n8272) );
  NAND4BXL U12573 ( .AN(n8283), .B(n8198), .C(n8284), .D(n8285), .Y(n8274) );
  OAI22X1 U12574 ( .A0(n8276), .A1(n8238), .B0(n8277), .B1(n8240), .Y(n8275)
         );
  AOI221X1 U12575 ( .A0(n10785), .A1(n10901), .B0(n5051), .B1(n10902), .C0(
        n10903), .Y(n10900) );
  NAND4BXL U12576 ( .AN(n10911), .B(n10826), .C(n10912), .D(n10913), .Y(n10902) );
  OAI22X1 U12577 ( .A0(n10904), .A1(n10866), .B0(n10905), .B1(n10868), .Y(
        n10903) );
  AOI221X1 U12578 ( .A0(n9033), .A1(n9149), .B0(n5557), .B1(n9150), .C0(n9151), 
        .Y(n9148) );
  NAND4BXL U12579 ( .AN(n9159), .B(n9074), .C(n9160), .D(n9161), .Y(n9150) );
  OAI22X1 U12580 ( .A0(n9152), .A1(n9114), .B0(n9153), .B1(n9116), .Y(n9151)
         );
  AOI221X1 U12581 ( .A0(n7281), .A1(n7397), .B0(n6021), .B1(n7398), .C0(n7399), 
        .Y(n7396) );
  NAND4BXL U12582 ( .AN(n7407), .B(n7322), .C(n7408), .D(n7409), .Y(n7398) );
  OAI22X1 U12583 ( .A0(n7400), .A1(n7362), .B0(n7401), .B1(n7364), .Y(n7399)
         );
  AOI221X1 U12584 ( .A0(n10201), .A1(n10317), .B0(n5237), .B1(n10318), .C0(
        n10319), .Y(n10316) );
  NAND4BXL U12585 ( .AN(n10327), .B(n10242), .C(n10328), .D(n10329), .Y(n10318) );
  OAI22X1 U12586 ( .A0(n10320), .A1(n10282), .B0(n10321), .B1(n10284), .Y(
        n10319) );
  AOI221X1 U12587 ( .A0(n9325), .A1(n9441), .B0(n5481), .B1(n9442), .C0(n9443), 
        .Y(n9440) );
  NAND4BXL U12588 ( .AN(n9451), .B(n9366), .C(n9452), .D(n9453), .Y(n9442) );
  OAI22X1 U12589 ( .A0(n9444), .A1(n9406), .B0(n9445), .B1(n9408), .Y(n9443)
         );
  AOI221X1 U12590 ( .A0(n8449), .A1(n8565), .B0(n5709), .B1(n8566), .C0(n8567), 
        .Y(n8564) );
  NAND4BXL U12591 ( .AN(n8575), .B(n8490), .C(n8576), .D(n8577), .Y(n8566) );
  OAI22X1 U12592 ( .A0(n8568), .A1(n8530), .B0(n8569), .B1(n8532), .Y(n8567)
         );
  AOI221X1 U12593 ( .A0(n7573), .A1(n7689), .B0(n5945), .B1(n7690), .C0(n7691), 
        .Y(n7688) );
  NAND4BXL U12594 ( .AN(n7699), .B(n7614), .C(n7700), .D(n7701), .Y(n7690) );
  OAI22X1 U12595 ( .A0(n7692), .A1(n7654), .B0(n7693), .B1(n7656), .Y(n7691)
         );
  AOI221X1 U12596 ( .A0(n11369), .A1(n11485), .B0(n4851), .B1(n11486), .C0(
        n11487), .Y(n11484) );
  NAND4BXL U12597 ( .AN(n11495), .B(n11410), .C(n11496), .D(n11497), .Y(n11486) );
  OAI22X1 U12598 ( .A0(n11488), .A1(n11450), .B0(n11489), .B1(n11452), .Y(
        n11487) );
  AOI221X1 U12599 ( .A0(n10493), .A1(n10609), .B0(n5159), .B1(n10610), .C0(
        n10611), .Y(n10608) );
  NAND4BXL U12600 ( .AN(n10619), .B(n10534), .C(n10620), .D(n10621), .Y(n10610) );
  OAI22X1 U12601 ( .A0(n10612), .A1(n10574), .B0(n10613), .B1(n10576), .Y(
        n10611) );
  AOI221X1 U12602 ( .A0(n9617), .A1(n9733), .B0(n5405), .B1(n9734), .C0(n9735), 
        .Y(n9732) );
  NAND4BXL U12603 ( .AN(n9743), .B(n9658), .C(n9744), .D(n9745), .Y(n9734) );
  OAI22X1 U12604 ( .A0(n9736), .A1(n9698), .B0(n9737), .B1(n9700), .Y(n9735)
         );
  AOI221X1 U12605 ( .A0(n8741), .A1(n8857), .B0(n5633), .B1(n8858), .C0(n8859), 
        .Y(n8856) );
  NAND4BXL U12606 ( .AN(n8867), .B(n8782), .C(n8868), .D(n8869), .Y(n8858) );
  OAI22X1 U12607 ( .A0(n8860), .A1(n8822), .B0(n8861), .B1(n8824), .Y(n8859)
         );
  AOI221X1 U12608 ( .A0(n7865), .A1(n7981), .B0(n5869), .B1(n7982), .C0(n7983), 
        .Y(n7980) );
  NAND4BXL U12609 ( .AN(n7991), .B(n7906), .C(n7992), .D(n7993), .Y(n7982) );
  OAI22X1 U12610 ( .A0(n7984), .A1(n7946), .B0(n7985), .B1(n7948), .Y(n7983)
         );
  AOI222X1 U12611 ( .A0(n2847), .A1(n10094), .B0(n9909), .B1(n10095), .C0(
        n5321), .C1(n10096), .Y(n10093) );
  NAND3X1 U12612 ( .A(n10099), .B(n9907), .C(n10100), .Y(n10095) );
  NAND4X1 U12613 ( .A(n10045), .B(n10051), .C(n10097), .D(n10098), .Y(n10096)
         );
  OAI221XL U12614 ( .A0(n2860), .A1(n10102), .B0(n90), .B1(n9895), .C0(n10103), 
        .Y(n10094) );
  AOI222X1 U12615 ( .A0(n3448), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n280), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n93), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n281), .C0(n6105), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n282), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n279) );
  NAND3X1 U12616 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n285), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n91), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n286), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n281) );
  NAND4X1 U12617 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n231), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n237), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n283), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n284), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n282) );
  OAI221XL U12618 ( .A0(n3461), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n288), 
        .B0(n91), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n78), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n289), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n280) );
  AOI222X1 U12619 ( .A0(n3207), .A1(n8342), .B0(n8157), .B1(n8343), .C0(n5793), 
        .C1(n8344), .Y(n8341) );
  NAND3X1 U12620 ( .A(n8347), .B(n8155), .C(n8348), .Y(n8343) );
  NAND4X1 U12621 ( .A(n8293), .B(n8299), .C(n8345), .D(n8346), .Y(n8344) );
  OAI221XL U12622 ( .A0(n3220), .A1(n8350), .B0(n93), .B1(n8143), .C0(n8351), 
        .Y(n8342) );
  AOI222X1 U12623 ( .A0(n2605), .A1(n11262), .B0(n11077), .B1(n11263), .C0(
        n4967), .C1(n11264), .Y(n11261) );
  NAND3X1 U12624 ( .A(n11267), .B(n11075), .C(n11268), .Y(n11263) );
  NAND4X1 U12625 ( .A(n11213), .B(n11219), .C(n11265), .D(n11266), .Y(n11264)
         );
  OAI221XL U12626 ( .A0(n2618), .A1(n11270), .B0(n92), .B1(n11063), .C0(n11271), .Y(n11262) );
  AOI222X1 U12627 ( .A0(n2666), .A1(n10970), .B0(n10785), .B1(n10971), .C0(
        n5051), .C1(n10972), .Y(n10969) );
  NAND3X1 U12628 ( .A(n10975), .B(n10783), .C(n10976), .Y(n10971) );
  NAND4X1 U12629 ( .A(n10921), .B(n10927), .C(n10973), .D(n10974), .Y(n10972)
         );
  OAI221XL U12630 ( .A0(n2679), .A1(n10978), .B0(n94), .B1(n10771), .C0(n10979), .Y(n10970) );
  AOI222X1 U12631 ( .A0(n3387), .A1(n7466), .B0(n7281), .B1(n7467), .C0(n6021), 
        .C1(n7468), .Y(n7465) );
  NAND3X1 U12632 ( .A(n7471), .B(n7279), .C(n7472), .Y(n7467) );
  NAND4X1 U12633 ( .A(n7417), .B(n7423), .C(n7469), .D(n7470), .Y(n7468) );
  OAI221XL U12634 ( .A0(n3400), .A1(n7474), .B0(n95), .B1(n7267), .C0(n7475), 
        .Y(n7466) );
  AOI222X1 U12635 ( .A0(n3027), .A1(n9218), .B0(n9033), .B1(n9219), .C0(n5557), 
        .C1(n9220), .Y(n9217) );
  NAND3X1 U12636 ( .A(n9223), .B(n9031), .C(n9224), .Y(n9219) );
  NAND4X1 U12637 ( .A(n9169), .B(n9175), .C(n9221), .D(n9222), .Y(n9220) );
  OAI221XL U12638 ( .A0(n3040), .A1(n9226), .B0(n96), .B1(n9019), .C0(n9227), 
        .Y(n9218) );
  AOI222X1 U12639 ( .A0(n2787), .A1(n10386), .B0(n10201), .B1(n10387), .C0(
        n5237), .C1(n10388), .Y(n10385) );
  NAND3X1 U12640 ( .A(n10391), .B(n10199), .C(n10392), .Y(n10387) );
  NAND4X1 U12641 ( .A(n10337), .B(n10343), .C(n10389), .D(n10390), .Y(n10388)
         );
  OAI221XL U12642 ( .A0(n2800), .A1(n10394), .B0(n97), .B1(n10187), .C0(n10395), .Y(n10386) );
  AOI222X1 U12643 ( .A0(n2969), .A1(n9510), .B0(n9325), .B1(n9511), .C0(n5481), 
        .C1(n9512), .Y(n9509) );
  NAND3X1 U12644 ( .A(n9515), .B(n9323), .C(n9516), .Y(n9511) );
  NAND4X1 U12645 ( .A(n9461), .B(n9467), .C(n9513), .D(n9514), .Y(n9512) );
  OAI221XL U12646 ( .A0(n2982), .A1(n9518), .B0(n98), .B1(n9311), .C0(n9519), 
        .Y(n9510) );
  AOI222X1 U12647 ( .A0(n3146), .A1(n8634), .B0(n8449), .B1(n8635), .C0(n5709), 
        .C1(n8636), .Y(n8633) );
  NAND3X1 U12648 ( .A(n8639), .B(n8447), .C(n8640), .Y(n8635) );
  NAND4X1 U12649 ( .A(n8585), .B(n8591), .C(n8637), .D(n8638), .Y(n8636) );
  OAI221XL U12650 ( .A0(n3159), .A1(n8642), .B0(n99), .B1(n8435), .C0(n8643), 
        .Y(n8634) );
  AOI222X1 U12651 ( .A0(n3329), .A1(n7758), .B0(n7573), .B1(n7759), .C0(n5945), 
        .C1(n7760), .Y(n7757) );
  NAND3X1 U12652 ( .A(n7763), .B(n7571), .C(n7764), .Y(n7759) );
  NAND4X1 U12653 ( .A(n7709), .B(n7715), .C(n7761), .D(n7762), .Y(n7760) );
  OAI221XL U12654 ( .A0(n3342), .A1(n7766), .B0(n100), .B1(n7559), .C0(n7767), 
        .Y(n7758) );
  AOI222X1 U12655 ( .A0(n2544), .A1(n11554), .B0(n11369), .B1(n11555), .C0(
        n4851), .C1(n11556), .Y(n11553) );
  NAND3X1 U12656 ( .A(n11559), .B(n11367), .C(n11560), .Y(n11555) );
  NAND4X1 U12657 ( .A(n11505), .B(n11511), .C(n11557), .D(n11558), .Y(n11556)
         );
  OAI221XL U12658 ( .A0(n2557), .A1(n11562), .B0(n101), .B1(n11355), .C0(
        n11563), .Y(n11554) );
  AOI222X1 U12659 ( .A0(n2726), .A1(n10678), .B0(n10493), .B1(n10679), .C0(
        n5159), .C1(n10680), .Y(n10677) );
  NAND3X1 U12660 ( .A(n10683), .B(n10491), .C(n10684), .Y(n10679) );
  NAND4X1 U12661 ( .A(n10629), .B(n10635), .C(n10681), .D(n10682), .Y(n10680)
         );
  OAI221XL U12662 ( .A0(n2739), .A1(n10686), .B0(n102), .B1(n10479), .C0(
        n10687), .Y(n10678) );
  AOI222X1 U12663 ( .A0(n2908), .A1(n9802), .B0(n9617), .B1(n9803), .C0(n5405), 
        .C1(n9804), .Y(n9801) );
  NAND3X1 U12664 ( .A(n9807), .B(n9615), .C(n9808), .Y(n9803) );
  NAND4X1 U12665 ( .A(n9753), .B(n9759), .C(n9805), .D(n9806), .Y(n9804) );
  OAI221XL U12666 ( .A0(n2921), .A1(n9810), .B0(n103), .B1(n9603), .C0(n9811), 
        .Y(n9802) );
  AOI222X1 U12667 ( .A0(n3088), .A1(n8926), .B0(n8741), .B1(n8927), .C0(n5633), 
        .C1(n8928), .Y(n8925) );
  NAND3X1 U12668 ( .A(n8931), .B(n8739), .C(n8932), .Y(n8927) );
  NAND4X1 U12669 ( .A(n8877), .B(n8883), .C(n8929), .D(n8930), .Y(n8928) );
  OAI221XL U12670 ( .A0(n3101), .A1(n8934), .B0(n104), .B1(n8727), .C0(n8935), 
        .Y(n8926) );
  AOI222X1 U12671 ( .A0(n3268), .A1(n8050), .B0(n7865), .B1(n8051), .C0(n5869), 
        .C1(n8052), .Y(n8049) );
  NAND3X1 U12672 ( .A(n8055), .B(n7863), .C(n8056), .Y(n8051) );
  NAND4X1 U12673 ( .A(n8001), .B(n8007), .C(n8053), .D(n8054), .Y(n8052) );
  OAI221XL U12674 ( .A0(n3281), .A1(n8058), .B0(n105), .B1(n7851), .C0(n8059), 
        .Y(n8050) );
  AOI222X1 U12675 ( .A0(n10049), .A1(n2853), .B0(n2856), .B1(n10050), .C0(
        n5333), .C1(n10040), .Y(n10022) );
  NAND4BXL U12676 ( .AN(n10038), .B(n10051), .C(n10011), .D(n10052), .Y(n10050) );
  NAND4X1 U12677 ( .A(n10011), .B(n9958), .C(n10053), .D(n10054), .Y(n10049)
         );
  AOI22X1 U12678 ( .A0(n698), .A1(n5392), .B0(n996), .B1(n433), .Y(n10052) );
  AOI222X1 U12679 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n235), .A1(n3454), 
        .B0(n3464), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n236), .C0(n6119), 
        .C1(top_core_EC_ss_gen_tbox_0__sboxs_r_n226), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n208) );
  NAND4BXL U12680 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n224), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n237), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n197), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n238), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n236) );
  NAND4X1 U12681 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n197), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n143), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n239), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n240), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n235) );
  AOI22X1 U12682 ( .A0(n699), .A1(n6176), .B0(n1139), .B1(n434), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n238) );
  AOI222X1 U12683 ( .A0(n11217), .A1(n2611), .B0(n2621), .B1(n11218), .C0(
        n4979), .C1(n11208), .Y(n11190) );
  NAND4BXL U12684 ( .AN(n11206), .B(n11219), .C(n11179), .D(n11220), .Y(n11218) );
  NAND4X1 U12685 ( .A(n11179), .B(n11126), .C(n11221), .D(n11222), .Y(n11217)
         );
  AOI22X1 U12686 ( .A0(n700), .A1(n5038), .B0(n940), .B1(n435), .Y(n11220) );
  AOI222X1 U12687 ( .A0(n8297), .A1(n3213), .B0(n3216), .B1(n8298), .C0(n5805), 
        .C1(n8288), .Y(n8270) );
  NAND4BXL U12688 ( .AN(n8286), .B(n8299), .C(n8259), .D(n8300), .Y(n8298) );
  NAND4X1 U12689 ( .A(n8259), .B(n8206), .C(n8301), .D(n8302), .Y(n8297) );
  AOI22X1 U12690 ( .A0(n701), .A1(n5864), .B0(n1080), .B1(n436), .Y(n8300) );
  AOI222X1 U12691 ( .A0(n10925), .A1(n2672), .B0(n2675), .B1(n10926), .C0(
        n5063), .C1(n10916), .Y(n10898) );
  NAND4BXL U12692 ( .AN(n10914), .B(n10927), .C(n10887), .D(n10928), .Y(n10926) );
  NAND4X1 U12693 ( .A(n10887), .B(n10834), .C(n10929), .D(n10930), .Y(n10925)
         );
  AOI22X1 U12694 ( .A0(n707), .A1(n5122), .B0(n954), .B1(n442), .Y(n10928) );
  AOI222X1 U12695 ( .A0(n9173), .A1(n3033), .B0(n3043), .B1(n9174), .C0(n5569), 
        .C1(n9164), .Y(n9146) );
  NAND4BXL U12696 ( .AN(n9162), .B(n9175), .C(n9135), .D(n9176), .Y(n9174) );
  NAND4X1 U12697 ( .A(n9135), .B(n9082), .C(n9177), .D(n9178), .Y(n9173) );
  AOI22X1 U12698 ( .A0(n709), .A1(n5628), .B0(n1038), .B1(n444), .Y(n9176) );
  AOI222X1 U12699 ( .A0(n7421), .A1(n3393), .B0(n3403), .B1(n7422), .C0(n6033), 
        .C1(n7412), .Y(n7394) );
  NAND4BXL U12700 ( .AN(n7410), .B(n7423), .C(n7383), .D(n7424), .Y(n7422) );
  NAND4X1 U12701 ( .A(n7383), .B(n7330), .C(n7425), .D(n7426), .Y(n7421) );
  AOI22X1 U12702 ( .A0(n711), .A1(n6092), .B0(n1122), .B1(n446), .Y(n7424) );
  AOI222X1 U12703 ( .A0(n10341), .A1(n2793), .B0(n2803), .B1(n10342), .C0(
        n5249), .C1(n10332), .Y(n10314) );
  NAND4BXL U12704 ( .AN(n10330), .B(n10343), .C(n10303), .D(n10344), .Y(n10342) );
  NAND4X1 U12705 ( .A(n10303), .B(n10250), .C(n10345), .D(n10346), .Y(n10341)
         );
  AOI22X1 U12706 ( .A0(n713), .A1(n5308), .B0(n982), .B1(n448), .Y(n10344) );
  AOI222X1 U12707 ( .A0(n9465), .A1(n2975), .B0(n2985), .B1(n9466), .C0(n5493), 
        .C1(n9456), .Y(n9438) );
  NAND4BXL U12708 ( .AN(n9454), .B(n9467), .C(n9427), .D(n9468), .Y(n9466) );
  NAND4X1 U12709 ( .A(n9427), .B(n9374), .C(n9469), .D(n9470), .Y(n9465) );
  AOI22X1 U12710 ( .A0(n706), .A1(n5552), .B0(n1024), .B1(n441), .Y(n9468) );
  AOI222X1 U12711 ( .A0(n8589), .A1(n3152), .B0(n3162), .B1(n8590), .C0(n5721), 
        .C1(n8580), .Y(n8562) );
  NAND4BXL U12712 ( .AN(n8578), .B(n8591), .C(n8551), .D(n8592), .Y(n8590) );
  NAND4X1 U12713 ( .A(n8551), .B(n8498), .C(n8593), .D(n8594), .Y(n8589) );
  AOI22X1 U12714 ( .A0(n702), .A1(n5780), .B0(n1066), .B1(n437), .Y(n8592) );
  AOI222X1 U12715 ( .A0(n7713), .A1(n3335), .B0(n3345), .B1(n7714), .C0(n5957), 
        .C1(n7704), .Y(n7686) );
  NAND4BXL U12716 ( .AN(n7702), .B(n7715), .C(n7675), .D(n7716), .Y(n7714) );
  NAND4X1 U12717 ( .A(n7675), .B(n7622), .C(n7717), .D(n7718), .Y(n7713) );
  AOI22X1 U12718 ( .A0(n708), .A1(n6016), .B0(n1108), .B1(n443), .Y(n7716) );
  AOI222X1 U12719 ( .A0(n11509), .A1(n2550), .B0(n2551), .B1(n11510), .C0(
        n4863), .C1(n11500), .Y(n11482) );
  NAND4BXL U12720 ( .AN(n11498), .B(n11511), .C(n11471), .D(n11512), .Y(n11510) );
  NAND4X1 U12721 ( .A(n11471), .B(n11418), .C(n11513), .D(n11514), .Y(n11509)
         );
  AOI22X1 U12722 ( .A0(n704), .A1(n4922), .B0(n926), .B1(n439), .Y(n11512) );
  AOI222X1 U12723 ( .A0(n10633), .A1(n2732), .B0(n2735), .B1(n10634), .C0(
        n5171), .C1(n10624), .Y(n10606) );
  NAND4BXL U12724 ( .AN(n10622), .B(n10635), .C(n10595), .D(n10636), .Y(n10634) );
  NAND4X1 U12725 ( .A(n10595), .B(n10542), .C(n10637), .D(n10638), .Y(n10633)
         );
  AOI22X1 U12726 ( .A0(n710), .A1(n5230), .B0(n968), .B1(n445), .Y(n10636) );
  AOI222X1 U12727 ( .A0(n9757), .A1(n2914), .B0(n2924), .B1(n9758), .C0(n5417), 
        .C1(n9748), .Y(n9730) );
  NAND4BXL U12728 ( .AN(n9746), .B(n9759), .C(n9719), .D(n9760), .Y(n9758) );
  NAND4X1 U12729 ( .A(n9719), .B(n9666), .C(n9761), .D(n9762), .Y(n9757) );
  AOI22X1 U12730 ( .A0(n703), .A1(n5476), .B0(n1010), .B1(n438), .Y(n9760) );
  AOI222X1 U12731 ( .A0(n8881), .A1(n3094), .B0(n3097), .B1(n8882), .C0(n5645), 
        .C1(n8872), .Y(n8854) );
  NAND4BXL U12732 ( .AN(n8870), .B(n8883), .C(n8843), .D(n8884), .Y(n8882) );
  NAND4X1 U12733 ( .A(n8843), .B(n8790), .C(n8885), .D(n8886), .Y(n8881) );
  AOI22X1 U12734 ( .A0(n712), .A1(n5704), .B0(n1052), .B1(n447), .Y(n8884) );
  AOI222X1 U12735 ( .A0(n8005), .A1(n3274), .B0(n3284), .B1(n8006), .C0(n5881), 
        .C1(n7996), .Y(n7978) );
  NAND4BXL U12736 ( .AN(n7994), .B(n8007), .C(n7967), .D(n8008), .Y(n8006) );
  NAND4X1 U12737 ( .A(n7967), .B(n7914), .C(n8009), .D(n8010), .Y(n8005) );
  AOI22X1 U12738 ( .A0(n705), .A1(n5940), .B0(n1094), .B1(n440), .Y(n8008) );
  NAND3BX1 U12739 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n86), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n87), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n88), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n84) );
  NAND3BX1 U12740 ( .AN(n9903), .B(n9904), .C(n9905), .Y(n9901) );
  NAND3BX1 U12741 ( .AN(n11071), .B(n11072), .C(n11073), .Y(n11069) );
  NAND3BX1 U12742 ( .AN(n8151), .B(n8152), .C(n8153), .Y(n8149) );
  NAND3BX1 U12743 ( .AN(n10779), .B(n10780), .C(n10781), .Y(n10777) );
  NAND3BX1 U12744 ( .AN(n9027), .B(n9028), .C(n9029), .Y(n9025) );
  NAND3BX1 U12745 ( .AN(n7275), .B(n7276), .C(n7277), .Y(n7273) );
  NAND3BX1 U12746 ( .AN(n10195), .B(n10196), .C(n10197), .Y(n10193) );
  NAND3BX1 U12747 ( .AN(n9319), .B(n9320), .C(n9321), .Y(n9317) );
  NAND3BX1 U12748 ( .AN(n8443), .B(n8444), .C(n8445), .Y(n8441) );
  NAND3BX1 U12749 ( .AN(n7567), .B(n7568), .C(n7569), .Y(n7565) );
  NAND3BX1 U12750 ( .AN(n11363), .B(n11364), .C(n11365), .Y(n11361) );
  NAND3BX1 U12751 ( .AN(n10487), .B(n10488), .C(n10489), .Y(n10485) );
  NAND3BX1 U12752 ( .AN(n9611), .B(n9612), .C(n9613), .Y(n9609) );
  NAND3BX1 U12753 ( .AN(n8735), .B(n8736), .C(n8737), .Y(n8733) );
  NAND3BX1 U12754 ( .AN(n7859), .B(n7860), .C(n7861), .Y(n7857) );
  AOI211X1 U12755 ( .A0(n6109), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n308), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n309), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n310), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n307) );
  NAND4BXL U12756 ( .AN(top_core_EC_ss_gen_tbox_0__sboxs_r_n287), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n133), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n140), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n319), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n308) );
  OAI2BB2X1 U12757 ( .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n313), .B1(n6110), 
        .A0N(n6105), .A1N(top_core_EC_ss_gen_tbox_0__sboxs_r_n314), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n309) );
  AOI21X1 U12758 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n311), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n312), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n176), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n310) );
  AOI211X1 U12759 ( .A0(n6107), .A1(n13841), .B0(n13842), .C0(n13843), .Y(
        n13840) );
  NAND4X1 U12760 ( .A(n13863), .B(n13864), .C(n13865), .D(n13866), .Y(n13841)
         );
  AOI31X1 U12761 ( .A0(n13844), .A1(n13845), .A2(n13846), .B0(n13847), .Y(
        n13843) );
  AOI31X1 U12762 ( .A0(n13850), .A1(n13851), .A2(n13852), .B0(n3448), .Y(
        n13842) );
  AOI211X1 U12763 ( .A0(n5322), .A1(n10122), .B0(n10123), .C0(n10124), .Y(
        n10121) );
  NAND4BXL U12764 ( .AN(n10101), .B(n9948), .C(n9955), .D(n10133), .Y(n10122)
         );
  OAI2BB2X1 U12765 ( .B0(n10127), .B1(n5323), .A0N(n5321), .A1N(n10128), .Y(
        n10123) );
  AOI21X1 U12766 ( .A0(n10125), .A1(n10126), .B0(n9990), .Y(n10124) );
  AOI211X1 U12767 ( .A0(n5325), .A1(n16991), .B0(n16992), .C0(n16993), .Y(
        n16990) );
  NAND4X1 U12768 ( .A(n17013), .B(n17014), .C(n17015), .D(n17016), .Y(n16991)
         );
  AOI31X1 U12769 ( .A0(n16994), .A1(n16995), .A2(n16996), .B0(n16997), .Y(
        n16993) );
  AOI31X1 U12770 ( .A0(n17000), .A1(n17001), .A2(n17002), .B0(n2847), .Y(
        n16992) );
  AOI211X1 U12771 ( .A0(n4968), .A1(n11290), .B0(n11291), .C0(n11292), .Y(
        n11289) );
  NAND4BXL U12772 ( .AN(n11269), .B(n11116), .C(n11123), .D(n11301), .Y(n11290) );
  OAI2BB2X1 U12773 ( .B0(n11295), .B1(n4969), .A0N(n4967), .A1N(n11296), .Y(
        n11291) );
  AOI21X1 U12774 ( .A0(n11293), .A1(n11294), .B0(n11158), .Y(n11292) );
  AOI211X1 U12775 ( .A0(n5794), .A1(n8370), .B0(n8371), .C0(n8372), .Y(n8369)
         );
  NAND4BXL U12776 ( .AN(n8349), .B(n8196), .C(n8203), .D(n8381), .Y(n8370) );
  OAI2BB2X1 U12777 ( .B0(n8375), .B1(n5795), .A0N(n5793), .A1N(n8376), .Y(
        n8371) );
  AOI21X1 U12778 ( .A0(n8373), .A1(n8374), .B0(n8238), .Y(n8372) );
  AOI211X1 U12779 ( .A0(n4971), .A1(n18251), .B0(n18252), .C0(n18253), .Y(
        n18250) );
  NAND4X1 U12780 ( .A(n18273), .B(n18274), .C(n18275), .D(n18276), .Y(n18251)
         );
  AOI31X1 U12781 ( .A0(n18254), .A1(n18255), .A2(n18256), .B0(n18257), .Y(
        n18253) );
  AOI31X1 U12782 ( .A0(n18260), .A1(n18261), .A2(n18262), .B0(n2605), .Y(
        n18252) );
  AOI211X1 U12783 ( .A0(n5797), .A1(n15101), .B0(n15102), .C0(n15103), .Y(
        n15100) );
  NAND4X1 U12784 ( .A(n15123), .B(n15124), .C(n15125), .D(n15126), .Y(n15101)
         );
  AOI31X1 U12785 ( .A0(n15104), .A1(n15105), .A2(n15106), .B0(n15107), .Y(
        n15103) );
  AOI31X1 U12786 ( .A0(n15110), .A1(n15111), .A2(n15112), .B0(n3207), .Y(
        n15102) );
  AOI211X1 U12787 ( .A0(n5713), .A1(n15416), .B0(n15417), .C0(n15418), .Y(
        n15415) );
  NAND4X1 U12788 ( .A(n15438), .B(n15439), .C(n15440), .D(n15441), .Y(n15416)
         );
  AOI31X1 U12789 ( .A0(n15419), .A1(n15420), .A2(n15421), .B0(n15422), .Y(
        n15418) );
  AOI31X1 U12790 ( .A0(n15425), .A1(n15426), .A2(n15427), .B0(n3146), .Y(
        n15417) );
  AOI211X1 U12791 ( .A0(n4855), .A1(n18566), .B0(n18567), .C0(n18568), .Y(
        n18565) );
  NAND4X1 U12792 ( .A(n18588), .B(n18589), .C(n18590), .D(n18591), .Y(n18566)
         );
  AOI31X1 U12793 ( .A0(n18569), .A1(n18570), .A2(n18571), .B0(n18572), .Y(
        n18568) );
  AOI31X1 U12794 ( .A0(n18575), .A1(n18576), .A2(n18577), .B0(n2544), .Y(
        n18567) );
  AOI211X1 U12795 ( .A0(n5409), .A1(n16676), .B0(n16677), .C0(n16678), .Y(
        n16675) );
  NAND4X1 U12796 ( .A(n16698), .B(n16699), .C(n16700), .D(n16701), .Y(n16676)
         );
  AOI31X1 U12797 ( .A0(n16679), .A1(n16680), .A2(n16681), .B0(n16682), .Y(
        n16678) );
  AOI31X1 U12798 ( .A0(n16685), .A1(n16686), .A2(n16687), .B0(n2908), .Y(
        n16677) );
  AOI211X1 U12799 ( .A0(n5052), .A1(n10998), .B0(n10999), .C0(n11000), .Y(
        n10997) );
  NAND4BXL U12800 ( .AN(n10977), .B(n10824), .C(n10831), .D(n11009), .Y(n10998) );
  OAI2BB2X1 U12801 ( .B0(n11003), .B1(n5053), .A0N(n5051), .A1N(n11004), .Y(
        n10999) );
  AOI21X1 U12802 ( .A0(n11001), .A1(n11002), .B0(n10866), .Y(n11000) );
  AOI211X1 U12803 ( .A0(n5558), .A1(n9246), .B0(n9247), .C0(n9248), .Y(n9245)
         );
  NAND4BXL U12804 ( .AN(n9225), .B(n9072), .C(n9079), .D(n9257), .Y(n9246) );
  OAI2BB2X1 U12805 ( .B0(n9251), .B1(n5559), .A0N(n5557), .A1N(n9252), .Y(
        n9247) );
  AOI21X1 U12806 ( .A0(n9249), .A1(n9250), .B0(n9114), .Y(n9248) );
  AOI211X1 U12807 ( .A0(n6022), .A1(n7494), .B0(n7495), .C0(n7496), .Y(n7493)
         );
  NAND4BXL U12808 ( .AN(n7473), .B(n7320), .C(n7327), .D(n7505), .Y(n7494) );
  OAI2BB2X1 U12809 ( .B0(n7499), .B1(n6023), .A0N(n6021), .A1N(n7500), .Y(
        n7495) );
  AOI21X1 U12810 ( .A0(n7497), .A1(n7498), .B0(n7362), .Y(n7496) );
  AOI211X1 U12811 ( .A0(n5238), .A1(n10414), .B0(n10415), .C0(n10416), .Y(
        n10413) );
  NAND4BXL U12812 ( .AN(n10393), .B(n10240), .C(n10247), .D(n10425), .Y(n10414) );
  OAI2BB2X1 U12813 ( .B0(n10419), .B1(n5239), .A0N(n5237), .A1N(n10420), .Y(
        n10415) );
  AOI21X1 U12814 ( .A0(n10417), .A1(n10418), .B0(n10282), .Y(n10416) );
  AOI211X1 U12815 ( .A0(n5873), .A1(n14786), .B0(n14787), .C0(n14788), .Y(
        n14785) );
  NAND4X1 U12816 ( .A(n14808), .B(n14809), .C(n14810), .D(n14811), .Y(n14786)
         );
  AOI31X1 U12817 ( .A0(n14789), .A1(n14790), .A2(n14791), .B0(n14792), .Y(
        n14788) );
  AOI31X1 U12818 ( .A0(n14795), .A1(n14796), .A2(n14797), .B0(n3268), .Y(
        n14787) );
  AOI211X1 U12819 ( .A0(n5482), .A1(n9538), .B0(n9539), .C0(n9540), .Y(n9537)
         );
  NAND4BXL U12820 ( .AN(n9517), .B(n9364), .C(n9371), .D(n9549), .Y(n9538) );
  OAI2BB2X1 U12821 ( .B0(n9543), .B1(n5483), .A0N(n5481), .A1N(n9544), .Y(
        n9539) );
  AOI21X1 U12822 ( .A0(n9541), .A1(n9542), .B0(n9406), .Y(n9540) );
  AOI211X1 U12823 ( .A0(n5485), .A1(n16361), .B0(n16362), .C0(n16363), .Y(
        n16360) );
  NAND4X1 U12824 ( .A(n16383), .B(n16384), .C(n16385), .D(n16386), .Y(n16361)
         );
  AOI31X1 U12825 ( .A0(n16364), .A1(n16365), .A2(n16366), .B0(n16367), .Y(
        n16363) );
  AOI31X1 U12826 ( .A0(n16370), .A1(n16371), .A2(n16372), .B0(n2969), .Y(
        n16362) );
  AOI211X1 U12827 ( .A0(n5710), .A1(n8662), .B0(n8663), .C0(n8664), .Y(n8661)
         );
  NAND4BXL U12828 ( .AN(n8641), .B(n8488), .C(n8495), .D(n8673), .Y(n8662) );
  OAI2BB2X1 U12829 ( .B0(n8667), .B1(n5711), .A0N(n5709), .A1N(n8668), .Y(
        n8663) );
  AOI21X1 U12830 ( .A0(n8665), .A1(n8666), .B0(n8530), .Y(n8664) );
  AOI211X1 U12831 ( .A0(n5055), .A1(n17936), .B0(n17937), .C0(n17938), .Y(
        n17935) );
  NAND4X1 U12832 ( .A(n17958), .B(n17959), .C(n17960), .D(n17961), .Y(n17936)
         );
  AOI31X1 U12833 ( .A0(n17939), .A1(n17940), .A2(n17941), .B0(n17942), .Y(
        n17938) );
  AOI31X1 U12834 ( .A0(n17945), .A1(n17946), .A2(n17947), .B0(n2666), .Y(
        n17937) );
  AOI211X1 U12835 ( .A0(n5946), .A1(n7786), .B0(n7787), .C0(n7788), .Y(n7785)
         );
  NAND4BXL U12836 ( .AN(n7765), .B(n7612), .C(n7619), .D(n7797), .Y(n7786) );
  OAI2BB2X1 U12837 ( .B0(n7791), .B1(n5947), .A0N(n5945), .A1N(n7792), .Y(
        n7787) );
  AOI21X1 U12838 ( .A0(n7789), .A1(n7790), .B0(n7654), .Y(n7788) );
  AOI211X1 U12839 ( .A0(n5949), .A1(n14471), .B0(n14472), .C0(n14473), .Y(
        n14470) );
  NAND4X1 U12840 ( .A(n14493), .B(n14494), .C(n14495), .D(n14496), .Y(n14471)
         );
  AOI31X1 U12841 ( .A0(n14474), .A1(n14475), .A2(n14476), .B0(n14477), .Y(
        n14473) );
  AOI31X1 U12842 ( .A0(n14480), .A1(n14481), .A2(n14482), .B0(n3329), .Y(
        n14472) );
  AOI211X1 U12843 ( .A0(n4852), .A1(n11582), .B0(n11583), .C0(n11584), .Y(
        n11581) );
  NAND4BXL U12844 ( .AN(n11561), .B(n11408), .C(n11415), .D(n11593), .Y(n11582) );
  OAI2BB2X1 U12845 ( .B0(n11587), .B1(n4853), .A0N(n4851), .A1N(n11588), .Y(
        n11583) );
  AOI21X1 U12846 ( .A0(n11585), .A1(n11586), .B0(n11450), .Y(n11584) );
  AOI211X1 U12847 ( .A0(n5561), .A1(n16046), .B0(n16047), .C0(n16048), .Y(
        n16045) );
  NAND4X1 U12848 ( .A(n16068), .B(n16069), .C(n16070), .D(n16071), .Y(n16046)
         );
  AOI31X1 U12849 ( .A0(n16049), .A1(n16050), .A2(n16051), .B0(n16052), .Y(
        n16048) );
  AOI31X1 U12850 ( .A0(n16055), .A1(n16056), .A2(n16057), .B0(n3027), .Y(
        n16047) );
  AOI211X1 U12851 ( .A0(n5160), .A1(n10706), .B0(n10707), .C0(n10708), .Y(
        n10705) );
  NAND4BXL U12852 ( .AN(n10685), .B(n10532), .C(n10539), .D(n10717), .Y(n10706) );
  OAI2BB2X1 U12853 ( .B0(n10711), .B1(n5161), .A0N(n5159), .A1N(n10712), .Y(
        n10707) );
  AOI21X1 U12854 ( .A0(n10709), .A1(n10710), .B0(n10574), .Y(n10708) );
  AOI211X1 U12855 ( .A0(n5163), .A1(n17621), .B0(n17622), .C0(n17623), .Y(
        n17620) );
  NAND4X1 U12856 ( .A(n17643), .B(n17644), .C(n17645), .D(n17646), .Y(n17621)
         );
  AOI31X1 U12857 ( .A0(n17624), .A1(n17625), .A2(n17626), .B0(n17627), .Y(
        n17623) );
  AOI31X1 U12858 ( .A0(n17630), .A1(n17631), .A2(n17632), .B0(n2726), .Y(
        n17622) );
  AOI211X1 U12859 ( .A0(n5406), .A1(n9830), .B0(n9831), .C0(n9832), .Y(n9829)
         );
  NAND4BXL U12860 ( .AN(n9809), .B(n9656), .C(n9663), .D(n9841), .Y(n9830) );
  OAI2BB2X1 U12861 ( .B0(n9835), .B1(n5407), .A0N(n5405), .A1N(n9836), .Y(
        n9831) );
  AOI21X1 U12862 ( .A0(n9833), .A1(n9834), .B0(n9698), .Y(n9832) );
  AOI211X1 U12863 ( .A0(n6025), .A1(n14156), .B0(n14157), .C0(n14158), .Y(
        n14155) );
  NAND4X1 U12864 ( .A(n14178), .B(n14179), .C(n14180), .D(n14181), .Y(n14156)
         );
  AOI31X1 U12865 ( .A0(n14159), .A1(n14160), .A2(n14161), .B0(n14162), .Y(
        n14158) );
  AOI31X1 U12866 ( .A0(n14165), .A1(n14166), .A2(n14167), .B0(n3387), .Y(
        n14157) );
  AOI211X1 U12867 ( .A0(n5634), .A1(n8954), .B0(n8955), .C0(n8956), .Y(n8953)
         );
  NAND4BXL U12868 ( .AN(n8933), .B(n8780), .C(n8787), .D(n8965), .Y(n8954) );
  OAI2BB2X1 U12869 ( .B0(n8959), .B1(n5635), .A0N(n5633), .A1N(n8960), .Y(
        n8955) );
  AOI21X1 U12870 ( .A0(n8957), .A1(n8958), .B0(n8822), .Y(n8956) );
  AOI211X1 U12871 ( .A0(n5637), .A1(n15731), .B0(n15732), .C0(n15733), .Y(
        n15730) );
  NAND4X1 U12872 ( .A(n15753), .B(n15754), .C(n15755), .D(n15756), .Y(n15731)
         );
  AOI31X1 U12873 ( .A0(n15734), .A1(n15735), .A2(n15736), .B0(n15737), .Y(
        n15733) );
  AOI31X1 U12874 ( .A0(n15740), .A1(n15741), .A2(n15742), .B0(n3088), .Y(
        n15732) );
  AOI211X1 U12875 ( .A0(n5870), .A1(n8078), .B0(n8079), .C0(n8080), .Y(n8077)
         );
  NAND4BXL U12876 ( .AN(n8057), .B(n7904), .C(n7911), .D(n8089), .Y(n8078) );
  OAI2BB2X1 U12877 ( .B0(n8083), .B1(n5871), .A0N(n5869), .A1N(n8084), .Y(
        n8079) );
  AOI21X1 U12878 ( .A0(n8081), .A1(n8082), .B0(n7946), .Y(n8080) );
  AOI211X1 U12879 ( .A0(n5241), .A1(n17306), .B0(n17307), .C0(n17308), .Y(
        n17305) );
  NAND4X1 U12880 ( .A(n17328), .B(n17329), .C(n17330), .D(n17331), .Y(n17306)
         );
  AOI31X1 U12881 ( .A0(n17309), .A1(n17310), .A2(n17311), .B0(n17312), .Y(
        n17308) );
  AOI31X1 U12882 ( .A0(n17315), .A1(n17316), .A2(n17317), .B0(n2787), .Y(
        n17307) );
  AOI211X1 U12883 ( .A0(n9909), .A1(n9980), .B0(n9981), .C0(n9982), .Y(n9979)
         );
  NAND4BXL U12884 ( .AN(n10000), .B(n9957), .C(n10001), .D(n10002), .Y(n9980)
         );
  OAI22X1 U12885 ( .A0(n9989), .A1(n9990), .B0(n9991), .B1(n9992), .Y(n9981)
         );
  AOI31X1 U12886 ( .A0(n9983), .A1(n5351), .A2(n9984), .B0(n9985), .Y(n9982)
         );
  AOI211X1 U12887 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n93), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n166), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n167), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n168), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n165) );
  NAND4BXL U12888 ( .AN(n265), .B(top_core_EC_ss_gen_tbox_0__sboxs_r_n142), 
        .C(top_core_EC_ss_gen_tbox_0__sboxs_r_n187), .D(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n188), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n166) );
  OAI22X1 U12889 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n175), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n176), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n177), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n178), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n167) );
  AOI31X1 U12890 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n169), .A1(n6147), 
        .A2(top_core_EC_ss_gen_tbox_0__sboxs_r_n170), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n171), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n168) );
  AOI211X1 U12891 ( .A0(n11077), .A1(n11148), .B0(n11149), .C0(n11150), .Y(
        n11147) );
  NAND4BXL U12892 ( .AN(n11168), .B(n11125), .C(n11169), .D(n11170), .Y(n11148) );
  OAI22X1 U12893 ( .A0(n11157), .A1(n11158), .B0(n11159), .B1(n11160), .Y(
        n11149) );
  AOI31X1 U12894 ( .A0(n11151), .A1(n4997), .A2(n11152), .B0(n11153), .Y(
        n11150) );
  AOI211X1 U12895 ( .A0(n8157), .A1(n8228), .B0(n8229), .C0(n8230), .Y(n8227)
         );
  NAND4BXL U12896 ( .AN(n264), .B(n8205), .C(n8249), .D(n8250), .Y(n8228) );
  OAI22X1 U12897 ( .A0(n8237), .A1(n8238), .B0(n8239), .B1(n8240), .Y(n8229)
         );
  AOI31X1 U12898 ( .A0(n8231), .A1(n5823), .A2(n8232), .B0(n8233), .Y(n8230)
         );
  AOI211X1 U12899 ( .A0(n10785), .A1(n10856), .B0(n10857), .C0(n10858), .Y(
        n10855) );
  NAND4BXL U12900 ( .AN(n10876), .B(n10833), .C(n10877), .D(n10878), .Y(n10856) );
  OAI22X1 U12901 ( .A0(n10865), .A1(n10866), .B0(n10867), .B1(n10868), .Y(
        n10857) );
  AOI31X1 U12902 ( .A0(n10859), .A1(n5081), .A2(n10860), .B0(n10861), .Y(
        n10858) );
  AOI211X1 U12903 ( .A0(n9033), .A1(n9104), .B0(n9105), .C0(n9106), .Y(n9103)
         );
  NAND4BXL U12904 ( .AN(n9124), .B(n9081), .C(n9125), .D(n9126), .Y(n9104) );
  OAI22X1 U12905 ( .A0(n9113), .A1(n9114), .B0(n9115), .B1(n9116), .Y(n9105)
         );
  AOI31X1 U12906 ( .A0(n9107), .A1(n5587), .A2(n9108), .B0(n9109), .Y(n9106)
         );
  AOI211X1 U12907 ( .A0(n7281), .A1(n7352), .B0(n7353), .C0(n7354), .Y(n7351)
         );
  NAND4BXL U12908 ( .AN(n7372), .B(n7329), .C(n7373), .D(n7374), .Y(n7352) );
  OAI22X1 U12909 ( .A0(n7361), .A1(n7362), .B0(n7363), .B1(n7364), .Y(n7353)
         );
  AOI31X1 U12910 ( .A0(n7355), .A1(n6051), .A2(n7356), .B0(n7357), .Y(n7354)
         );
  AOI211X1 U12911 ( .A0(n10201), .A1(n10272), .B0(n10273), .C0(n10274), .Y(
        n10271) );
  NAND4BXL U12912 ( .AN(n10292), .B(n10249), .C(n10293), .D(n10294), .Y(n10272) );
  OAI22X1 U12913 ( .A0(n10281), .A1(n10282), .B0(n10283), .B1(n10284), .Y(
        n10273) );
  AOI31X1 U12914 ( .A0(n10275), .A1(n5267), .A2(n10276), .B0(n10277), .Y(
        n10274) );
  AOI211X1 U12915 ( .A0(n9325), .A1(n9396), .B0(n9397), .C0(n9398), .Y(n9395)
         );
  NAND4BXL U12916 ( .AN(n9416), .B(n9373), .C(n9417), .D(n9418), .Y(n9396) );
  OAI22X1 U12917 ( .A0(n9405), .A1(n9406), .B0(n9407), .B1(n9408), .Y(n9397)
         );
  AOI31X1 U12918 ( .A0(n9399), .A1(n5511), .A2(n9400), .B0(n9401), .Y(n9398)
         );
  AOI211X1 U12919 ( .A0(n8449), .A1(n8520), .B0(n8521), .C0(n8522), .Y(n8519)
         );
  NAND4BXL U12920 ( .AN(n8540), .B(n8497), .C(n8541), .D(n8542), .Y(n8520) );
  OAI22X1 U12921 ( .A0(n8529), .A1(n8530), .B0(n8531), .B1(n8532), .Y(n8521)
         );
  AOI31X1 U12922 ( .A0(n8523), .A1(n5739), .A2(n8524), .B0(n8525), .Y(n8522)
         );
  AOI211X1 U12923 ( .A0(n7573), .A1(n7644), .B0(n7645), .C0(n7646), .Y(n7643)
         );
  NAND4BXL U12924 ( .AN(n7664), .B(n7621), .C(n7665), .D(n7666), .Y(n7644) );
  OAI22X1 U12925 ( .A0(n7653), .A1(n7654), .B0(n7655), .B1(n7656), .Y(n7645)
         );
  AOI31X1 U12926 ( .A0(n7647), .A1(n5975), .A2(n7648), .B0(n7649), .Y(n7646)
         );
  AOI211X1 U12927 ( .A0(n11369), .A1(n11440), .B0(n11441), .C0(n11442), .Y(
        n11439) );
  NAND4BXL U12928 ( .AN(n11460), .B(n11417), .C(n11461), .D(n11462), .Y(n11440) );
  OAI22X1 U12929 ( .A0(n11449), .A1(n11450), .B0(n11451), .B1(n11452), .Y(
        n11441) );
  AOI31X1 U12930 ( .A0(n11443), .A1(n4881), .A2(n11444), .B0(n11445), .Y(
        n11442) );
  AOI211X1 U12931 ( .A0(n10493), .A1(n10564), .B0(n10565), .C0(n10566), .Y(
        n10563) );
  NAND4BXL U12932 ( .AN(n10584), .B(n10541), .C(n10585), .D(n10586), .Y(n10564) );
  OAI22X1 U12933 ( .A0(n10573), .A1(n10574), .B0(n10575), .B1(n10576), .Y(
        n10565) );
  AOI31X1 U12934 ( .A0(n10567), .A1(n5189), .A2(n10568), .B0(n10569), .Y(
        n10566) );
  AOI211X1 U12935 ( .A0(n9617), .A1(n9688), .B0(n9689), .C0(n9690), .Y(n9687)
         );
  NAND4BXL U12936 ( .AN(n9708), .B(n9665), .C(n9709), .D(n9710), .Y(n9688) );
  OAI22X1 U12937 ( .A0(n9697), .A1(n9698), .B0(n9699), .B1(n9700), .Y(n9689)
         );
  AOI31X1 U12938 ( .A0(n9691), .A1(n5435), .A2(n9692), .B0(n9693), .Y(n9690)
         );
  AOI211X1 U12939 ( .A0(n8741), .A1(n8812), .B0(n8813), .C0(n8814), .Y(n8811)
         );
  NAND4BXL U12940 ( .AN(n8832), .B(n8789), .C(n8833), .D(n8834), .Y(n8812) );
  OAI22X1 U12941 ( .A0(n8821), .A1(n8822), .B0(n8823), .B1(n8824), .Y(n8813)
         );
  AOI31X1 U12942 ( .A0(n8815), .A1(n5663), .A2(n8816), .B0(n8817), .Y(n8814)
         );
  AOI211X1 U12943 ( .A0(n7865), .A1(n7936), .B0(n7937), .C0(n7938), .Y(n7935)
         );
  NAND4BXL U12944 ( .AN(n7956), .B(n7913), .C(n7957), .D(n7958), .Y(n7936) );
  OAI22X1 U12945 ( .A0(n7945), .A1(n7946), .B0(n7947), .B1(n7948), .Y(n7937)
         );
  AOI31X1 U12946 ( .A0(n7939), .A1(n5899), .A2(n7940), .B0(n7941), .Y(n7938)
         );
  AOI211X1 U12947 ( .A0(n13860), .A1(n1137), .B0(n13888), .C0(n13889), .Y(
        n13836) );
  OAI21XL U12948 ( .A0(n3467), .A1(n13890), .B0(n13891), .Y(n13889) );
  OAI222XL U12949 ( .A0(n13880), .A1(n13878), .B0(n3462), .B1(n13892), .C0(
        n13893), .C1(n3453), .Y(n13888) );
  AOI211X1 U12950 ( .A0(n17010), .A1(n998), .B0(n17038), .C0(n17039), .Y(
        n16986) );
  OAI21XL U12951 ( .A0(n2866), .A1(n17040), .B0(n17041), .Y(n17039) );
  OAI222XL U12952 ( .A0(n17030), .A1(n17028), .B0(n2861), .B1(n17042), .C0(
        n17043), .C1(n2852), .Y(n17038) );
  AOI211X1 U12953 ( .A0(n18270), .A1(n942), .B0(n18298), .C0(n18299), .Y(
        n18246) );
  OAI21XL U12954 ( .A0(n2624), .A1(n18300), .B0(n18301), .Y(n18299) );
  OAI222XL U12955 ( .A0(n18290), .A1(n18288), .B0(n2619), .B1(n18302), .C0(
        n18303), .C1(n2610), .Y(n18298) );
  AOI211X1 U12956 ( .A0(n15120), .A1(n1082), .B0(n15148), .C0(n15149), .Y(
        n15096) );
  OAI21XL U12957 ( .A0(n3226), .A1(n15150), .B0(n15151), .Y(n15149) );
  OAI222XL U12958 ( .A0(n15140), .A1(n15138), .B0(n3221), .B1(n15152), .C0(
        n15153), .C1(n3212), .Y(n15148) );
  AOI211X1 U12959 ( .A0(n15435), .A1(n1068), .B0(n15463), .C0(n15464), .Y(
        n15411) );
  OAI21XL U12960 ( .A0(n3165), .A1(n15465), .B0(n15466), .Y(n15464) );
  OAI222XL U12961 ( .A0(n15455), .A1(n15453), .B0(n3160), .B1(n15467), .C0(
        n15468), .C1(n3151), .Y(n15463) );
  AOI211X1 U12962 ( .A0(n18585), .A1(n928), .B0(n18613), .C0(n18614), .Y(
        n18561) );
  OAI21XL U12963 ( .A0(n2563), .A1(n18615), .B0(n18616), .Y(n18614) );
  OAI222XL U12964 ( .A0(n18605), .A1(n18603), .B0(n2552), .B1(n18617), .C0(
        n18618), .C1(n2549), .Y(n18613) );
  AOI211X1 U12965 ( .A0(n16695), .A1(n1012), .B0(n16723), .C0(n16724), .Y(
        n16671) );
  OAI21XL U12966 ( .A0(n2927), .A1(n16725), .B0(n16726), .Y(n16724) );
  OAI222XL U12967 ( .A0(n16715), .A1(n16713), .B0(n2922), .B1(n16727), .C0(
        n16728), .C1(n2913), .Y(n16723) );
  AOI211X1 U12968 ( .A0(n14805), .A1(n1096), .B0(n14833), .C0(n14834), .Y(
        n14781) );
  OAI21XL U12969 ( .A0(n3287), .A1(n14835), .B0(n14836), .Y(n14834) );
  OAI222XL U12970 ( .A0(n14825), .A1(n14823), .B0(n3282), .B1(n14837), .C0(
        n14838), .C1(n3273), .Y(n14833) );
  AOI211X1 U12971 ( .A0(n16380), .A1(n1026), .B0(n16408), .C0(n16409), .Y(
        n16356) );
  OAI21XL U12972 ( .A0(n2988), .A1(n16410), .B0(n16411), .Y(n16409) );
  OAI222XL U12973 ( .A0(n16400), .A1(n16398), .B0(n2983), .B1(n16412), .C0(
        n16413), .C1(n2974), .Y(n16408) );
  AOI211X1 U12974 ( .A0(n17955), .A1(n956), .B0(n17983), .C0(n17984), .Y(
        n17931) );
  OAI21XL U12975 ( .A0(n2685), .A1(n17985), .B0(n17986), .Y(n17984) );
  OAI222XL U12976 ( .A0(n17975), .A1(n17973), .B0(n2680), .B1(n17987), .C0(
        n17988), .C1(n2671), .Y(n17983) );
  AOI211X1 U12977 ( .A0(n14490), .A1(n1110), .B0(n14518), .C0(n14519), .Y(
        n14466) );
  OAI21XL U12978 ( .A0(n3348), .A1(n14520), .B0(n14521), .Y(n14519) );
  OAI222XL U12979 ( .A0(n14510), .A1(n14508), .B0(n3343), .B1(n14522), .C0(
        n14523), .C1(n3334), .Y(n14518) );
  AOI211X1 U12980 ( .A0(n16065), .A1(n1040), .B0(n16093), .C0(n16094), .Y(
        n16041) );
  OAI21XL U12981 ( .A0(n3046), .A1(n16095), .B0(n16096), .Y(n16094) );
  OAI222XL U12982 ( .A0(n16085), .A1(n16083), .B0(n3041), .B1(n16097), .C0(
        n16098), .C1(n3032), .Y(n16093) );
  AOI211X1 U12983 ( .A0(n17640), .A1(n970), .B0(n17668), .C0(n17669), .Y(
        n17616) );
  OAI21XL U12984 ( .A0(n2745), .A1(n17670), .B0(n17671), .Y(n17669) );
  OAI222XL U12985 ( .A0(n17660), .A1(n17658), .B0(n2740), .B1(n17672), .C0(
        n17673), .C1(n2731), .Y(n17668) );
  AOI211X1 U12986 ( .A0(n14175), .A1(n1124), .B0(n14203), .C0(n14204), .Y(
        n14151) );
  OAI21XL U12987 ( .A0(n3406), .A1(n14205), .B0(n14206), .Y(n14204) );
  OAI222XL U12988 ( .A0(n14195), .A1(n14193), .B0(n3401), .B1(n14207), .C0(
        n14208), .C1(n3392), .Y(n14203) );
  AOI211X1 U12989 ( .A0(n15750), .A1(n1054), .B0(n15778), .C0(n15779), .Y(
        n15726) );
  OAI21XL U12990 ( .A0(n3107), .A1(n15780), .B0(n15781), .Y(n15779) );
  OAI222XL U12991 ( .A0(n15770), .A1(n15768), .B0(n3102), .B1(n15782), .C0(
        n15783), .C1(n3093), .Y(n15778) );
  AOI211X1 U12992 ( .A0(n17325), .A1(n984), .B0(n17353), .C0(n17354), .Y(
        n17301) );
  OAI21XL U12993 ( .A0(n2806), .A1(n17355), .B0(n17356), .Y(n17354) );
  OAI222XL U12994 ( .A0(n17345), .A1(n17343), .B0(n2801), .B1(n17357), .C0(
        n17358), .C1(n2792), .Y(n17353) );
  NAND3X1 U12995 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n237), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n67), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n329), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n325) );
  OAI22X1 U12996 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n78), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n98), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n327), .B1(n3452), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n326) );
  AOI2BB2X1 U12997 ( .B0(n1143), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n82), 
        .A0N(top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .A1N(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n162), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n329) );
  NAND3X1 U12998 ( .A(n10051), .B(n9885), .C(n10143), .Y(n10139) );
  OAI22X1 U12999 ( .A0(n9895), .A1(n9914), .B0(n10141), .B1(n2851), .Y(n10140)
         );
  AOI2BB2X1 U13000 ( .B0(n1001), .B1(n9899), .A0N(n9913), .A1N(n9976), .Y(
        n10143) );
  NAND3X1 U13001 ( .A(n11219), .B(n11053), .C(n11311), .Y(n11307) );
  OAI22X1 U13002 ( .A0(n11063), .A1(n11082), .B0(n11309), .B1(n2609), .Y(
        n11308) );
  AOI2BB2X1 U13003 ( .B0(n945), .B1(n11067), .A0N(n11081), .A1N(n11144), .Y(
        n11311) );
  NAND3X1 U13004 ( .A(n8299), .B(n8133), .C(n8391), .Y(n8387) );
  OAI22X1 U13005 ( .A0(n8143), .A1(n8162), .B0(n8389), .B1(n3211), .Y(n8388)
         );
  AOI2BB2X1 U13006 ( .B0(n1085), .B1(n8147), .A0N(n8161), .A1N(n8224), .Y(
        n8391) );
  NAND3X1 U13007 ( .A(n10927), .B(n10761), .C(n11019), .Y(n11015) );
  OAI22X1 U13008 ( .A0(n10771), .A1(n10790), .B0(n11017), .B1(n2670), .Y(
        n11016) );
  AOI2BB2X1 U13009 ( .B0(n959), .B1(n10775), .A0N(n10789), .A1N(n10852), .Y(
        n11019) );
  NAND3X1 U13010 ( .A(n9175), .B(n9009), .C(n9267), .Y(n9263) );
  OAI22X1 U13011 ( .A0(n9019), .A1(n9038), .B0(n9265), .B1(n3031), .Y(n9264)
         );
  AOI2BB2X1 U13012 ( .B0(n1043), .B1(n9023), .A0N(n9037), .A1N(n9100), .Y(
        n9267) );
  NAND3X1 U13013 ( .A(n7423), .B(n7257), .C(n7515), .Y(n7511) );
  OAI22X1 U13014 ( .A0(n7267), .A1(n7286), .B0(n7513), .B1(n3391), .Y(n7512)
         );
  AOI2BB2X1 U13015 ( .B0(n1127), .B1(n7271), .A0N(n7285), .A1N(n7348), .Y(
        n7515) );
  NAND3X1 U13016 ( .A(n10343), .B(n10177), .C(n10435), .Y(n10431) );
  OAI22X1 U13017 ( .A0(n10187), .A1(n10206), .B0(n10433), .B1(n2791), .Y(
        n10432) );
  AOI2BB2X1 U13018 ( .B0(n987), .B1(n10191), .A0N(n10205), .A1N(n10268), .Y(
        n10435) );
  NAND3X1 U13019 ( .A(n9467), .B(n9301), .C(n9559), .Y(n9555) );
  OAI22X1 U13020 ( .A0(n9311), .A1(n9330), .B0(n9557), .B1(n2973), .Y(n9556)
         );
  AOI2BB2X1 U13021 ( .B0(n1029), .B1(n9315), .A0N(n9329), .A1N(n9392), .Y(
        n9559) );
  NAND3X1 U13022 ( .A(n8591), .B(n8425), .C(n8683), .Y(n8679) );
  OAI22X1 U13023 ( .A0(n8435), .A1(n8454), .B0(n8681), .B1(n3150), .Y(n8680)
         );
  AOI2BB2X1 U13024 ( .B0(n1071), .B1(n8439), .A0N(n8453), .A1N(n8516), .Y(
        n8683) );
  NAND3X1 U13025 ( .A(n7715), .B(n7549), .C(n7807), .Y(n7803) );
  OAI22X1 U13026 ( .A0(n7559), .A1(n7578), .B0(n7805), .B1(n3333), .Y(n7804)
         );
  AOI2BB2X1 U13027 ( .B0(n1113), .B1(n7563), .A0N(n7577), .A1N(n7640), .Y(
        n7807) );
  NAND3X1 U13028 ( .A(n11511), .B(n11345), .C(n11603), .Y(n11599) );
  OAI22X1 U13029 ( .A0(n11355), .A1(n11374), .B0(n11601), .B1(n2548), .Y(
        n11600) );
  AOI2BB2X1 U13030 ( .B0(n931), .B1(n11359), .A0N(n11373), .A1N(n11436), .Y(
        n11603) );
  NAND3X1 U13031 ( .A(n10635), .B(n10469), .C(n10727), .Y(n10723) );
  OAI22X1 U13032 ( .A0(n10479), .A1(n10498), .B0(n10725), .B1(n2730), .Y(
        n10724) );
  AOI2BB2X1 U13033 ( .B0(n973), .B1(n10483), .A0N(n10497), .A1N(n10560), .Y(
        n10727) );
  NAND3X1 U13034 ( .A(n9759), .B(n9593), .C(n9851), .Y(n9847) );
  OAI22X1 U13035 ( .A0(n9603), .A1(n9622), .B0(n9849), .B1(n2912), .Y(n9848)
         );
  AOI2BB2X1 U13036 ( .B0(n1015), .B1(n9607), .A0N(n9621), .A1N(n9684), .Y(
        n9851) );
  NAND3X1 U13037 ( .A(n8883), .B(n8717), .C(n8975), .Y(n8971) );
  OAI22X1 U13038 ( .A0(n8727), .A1(n8746), .B0(n8973), .B1(n3092), .Y(n8972)
         );
  AOI2BB2X1 U13039 ( .B0(n1057), .B1(n8731), .A0N(n8745), .A1N(n8808), .Y(
        n8975) );
  NAND3X1 U13040 ( .A(n8007), .B(n7841), .C(n8099), .Y(n8095) );
  OAI22X1 U13041 ( .A0(n7851), .A1(n7870), .B0(n8097), .B1(n3272), .Y(n8096)
         );
  AOI2BB2X1 U13042 ( .B0(n1099), .B1(n7855), .A0N(n7869), .A1N(n7932), .Y(
        n8099) );
  INVX1 U13043 ( .A(n13375), .Y(n6547) );
  INVX1 U13044 ( .A(n12745), .Y(n6842) );
  INVX1 U13045 ( .A(n13690), .Y(n6595) );
  INVX1 U13046 ( .A(n13060), .Y(n6888) );
  AOI211X1 U13047 ( .A0(n5357), .A1(n2882), .B0(n17127), .C0(n17128), .Y(
        n17124) );
  NAND4X1 U13048 ( .A(n17110), .B(n17130), .C(n17026), .D(n17114), .Y(n17127)
         );
  OAI21XL U13049 ( .A0(n450), .A1(n17062), .B0(n17129), .Y(n17128) );
  AOI211X1 U13050 ( .A0(n6125), .A1(n3483), .B0(n13977), .C0(n13978), .Y(
        n13974) );
  NAND4X1 U13051 ( .A(n13960), .B(n13980), .C(n13876), .D(n13964), .Y(n13977)
         );
  OAI21XL U13052 ( .A0(n449), .A1(n13912), .B0(n13979), .Y(n13978) );
  AOI211X1 U13053 ( .A0(n5003), .A1(n2640), .B0(n18387), .C0(n18388), .Y(
        n18384) );
  NAND4X1 U13054 ( .A(n18370), .B(n18390), .C(n18286), .D(n18374), .Y(n18387)
         );
  OAI21XL U13055 ( .A0(n451), .A1(n18322), .B0(n18389), .Y(n18388) );
  AOI211X1 U13056 ( .A0(n5829), .A1(n3242), .B0(n15237), .C0(n15238), .Y(
        n15234) );
  NAND4X1 U13057 ( .A(n15220), .B(n15240), .C(n15136), .D(n15224), .Y(n15237)
         );
  OAI21XL U13058 ( .A0(n452), .A1(n15172), .B0(n15239), .Y(n15238) );
  AOI211X1 U13059 ( .A0(n5745), .A1(n3181), .B0(n15552), .C0(n15553), .Y(
        n15549) );
  NAND4X1 U13060 ( .A(n15535), .B(n15555), .C(n15451), .D(n15539), .Y(n15552)
         );
  OAI21XL U13061 ( .A0(n453), .A1(n15487), .B0(n15554), .Y(n15553) );
  AOI211X1 U13062 ( .A0(n4887), .A1(n2579), .B0(n18702), .C0(n18703), .Y(
        n18699) );
  NAND4X1 U13063 ( .A(n18685), .B(n18705), .C(n18601), .D(n18689), .Y(n18702)
         );
  OAI21XL U13064 ( .A0(n454), .A1(n18637), .B0(n18704), .Y(n18703) );
  AOI211X1 U13065 ( .A0(n5441), .A1(n2943), .B0(n16812), .C0(n16813), .Y(
        n16809) );
  NAND4X1 U13066 ( .A(n16795), .B(n16815), .C(n16711), .D(n16799), .Y(n16812)
         );
  OAI21XL U13067 ( .A0(n455), .A1(n16747), .B0(n16814), .Y(n16813) );
  AOI211X1 U13068 ( .A0(n5905), .A1(n3303), .B0(n14922), .C0(n14923), .Y(
        n14919) );
  NAND4X1 U13069 ( .A(n14905), .B(n14925), .C(n14821), .D(n14909), .Y(n14922)
         );
  OAI21XL U13070 ( .A0(n456), .A1(n14857), .B0(n14924), .Y(n14923) );
  AOI211X1 U13071 ( .A0(n5517), .A1(n3004), .B0(n16497), .C0(n16498), .Y(
        n16494) );
  NAND4X1 U13072 ( .A(n16480), .B(n16500), .C(n16396), .D(n16484), .Y(n16497)
         );
  OAI21XL U13073 ( .A0(n457), .A1(n16432), .B0(n16499), .Y(n16498) );
  AOI211X1 U13074 ( .A0(n5087), .A1(n2701), .B0(n18072), .C0(n18073), .Y(
        n18069) );
  NAND4X1 U13075 ( .A(n18055), .B(n18075), .C(n17971), .D(n18059), .Y(n18072)
         );
  OAI21XL U13076 ( .A0(n458), .A1(n18007), .B0(n18074), .Y(n18073) );
  AOI211X1 U13077 ( .A0(n5981), .A1(n3364), .B0(n14607), .C0(n14608), .Y(
        n14604) );
  NAND4X1 U13078 ( .A(n14590), .B(n14610), .C(n14506), .D(n14594), .Y(n14607)
         );
  OAI21XL U13079 ( .A0(n459), .A1(n14542), .B0(n14609), .Y(n14608) );
  AOI211X1 U13080 ( .A0(n5593), .A1(n3062), .B0(n16182), .C0(n16183), .Y(
        n16179) );
  NAND4X1 U13081 ( .A(n16165), .B(n16185), .C(n16081), .D(n16169), .Y(n16182)
         );
  OAI21XL U13082 ( .A0(n460), .A1(n16117), .B0(n16184), .Y(n16183) );
  AOI211X1 U13083 ( .A0(n5195), .A1(n2761), .B0(n17757), .C0(n17758), .Y(
        n17754) );
  NAND4X1 U13084 ( .A(n17740), .B(n17760), .C(n17656), .D(n17744), .Y(n17757)
         );
  OAI21XL U13085 ( .A0(n461), .A1(n17692), .B0(n17759), .Y(n17758) );
  AOI211X1 U13086 ( .A0(n6057), .A1(n3422), .B0(n14292), .C0(n14293), .Y(
        n14289) );
  NAND4X1 U13087 ( .A(n14275), .B(n14295), .C(n14191), .D(n14279), .Y(n14292)
         );
  OAI21XL U13088 ( .A0(n462), .A1(n14227), .B0(n14294), .Y(n14293) );
  AOI211X1 U13089 ( .A0(n5669), .A1(n3123), .B0(n15867), .C0(n15868), .Y(
        n15864) );
  NAND4X1 U13090 ( .A(n15850), .B(n15870), .C(n15766), .D(n15854), .Y(n15867)
         );
  OAI21XL U13091 ( .A0(n463), .A1(n15802), .B0(n15869), .Y(n15868) );
  AOI211X1 U13092 ( .A0(n5273), .A1(n2822), .B0(n17442), .C0(n17443), .Y(
        n17439) );
  NAND4X1 U13093 ( .A(n17425), .B(n17445), .C(n17341), .D(n17429), .Y(n17442)
         );
  OAI21XL U13094 ( .A0(n464), .A1(n17377), .B0(n17444), .Y(n17443) );
  AOI211X1 U13095 ( .A0(n17183), .A1(n1003), .B0(n17184), .C0(n17185), .Y(
        n17182) );
  AOI21X1 U13096 ( .A0(n17186), .A1(n17187), .B0(n2852), .Y(n17184) );
  AOI211X1 U13097 ( .A0(n5357), .A1(n2882), .B0(n17098), .C0(n17188), .Y(
        n17187) );
  AOI211X1 U13098 ( .A0(n14033), .A1(n1142), .B0(n14034), .C0(n14035), .Y(
        n14032) );
  AOI21X1 U13099 ( .A0(n14036), .A1(n14037), .B0(n3453), .Y(n14034) );
  AOI211X1 U13100 ( .A0(n6125), .A1(n3483), .B0(n13948), .C0(n14038), .Y(
        n14037) );
  AOI211X1 U13101 ( .A0(n18443), .A1(n947), .B0(n18444), .C0(n18445), .Y(
        n18442) );
  AOI21X1 U13102 ( .A0(n18446), .A1(n18447), .B0(n2610), .Y(n18444) );
  AOI211X1 U13103 ( .A0(n5003), .A1(n2640), .B0(n18358), .C0(n18448), .Y(
        n18447) );
  AOI211X1 U13104 ( .A0(n15293), .A1(n1087), .B0(n15294), .C0(n15295), .Y(
        n15292) );
  AOI21X1 U13105 ( .A0(n15296), .A1(n15297), .B0(n3212), .Y(n15294) );
  AOI211X1 U13106 ( .A0(n5829), .A1(n3242), .B0(n15208), .C0(n15298), .Y(
        n15297) );
  AOI211X1 U13107 ( .A0(n15608), .A1(n1073), .B0(n15609), .C0(n15610), .Y(
        n15607) );
  AOI21X1 U13108 ( .A0(n15611), .A1(n15612), .B0(n3151), .Y(n15609) );
  AOI211X1 U13109 ( .A0(n5745), .A1(n3181), .B0(n15523), .C0(n15613), .Y(
        n15612) );
  AOI211X1 U13110 ( .A0(n16868), .A1(n1017), .B0(n16869), .C0(n16870), .Y(
        n16867) );
  AOI21X1 U13111 ( .A0(n16871), .A1(n16872), .B0(n2913), .Y(n16869) );
  AOI211X1 U13112 ( .A0(n5441), .A1(n2943), .B0(n16783), .C0(n16873), .Y(
        n16872) );
  AOI211X1 U13113 ( .A0(n18758), .A1(n933), .B0(n18759), .C0(n18760), .Y(
        n18757) );
  AOI21X1 U13114 ( .A0(n18761), .A1(n18762), .B0(n2549), .Y(n18759) );
  AOI211X1 U13115 ( .A0(n4887), .A1(n2579), .B0(n18673), .C0(n18763), .Y(
        n18762) );
  AOI211X1 U13116 ( .A0(n14978), .A1(n1101), .B0(n14979), .C0(n14980), .Y(
        n14977) );
  AOI21X1 U13117 ( .A0(n14981), .A1(n14982), .B0(n3273), .Y(n14979) );
  AOI211X1 U13118 ( .A0(n5905), .A1(n3303), .B0(n14893), .C0(n14983), .Y(
        n14982) );
  AOI211X1 U13119 ( .A0(n16553), .A1(n1031), .B0(n16554), .C0(n16555), .Y(
        n16552) );
  AOI21X1 U13120 ( .A0(n16556), .A1(n16557), .B0(n2974), .Y(n16554) );
  AOI211X1 U13121 ( .A0(n5517), .A1(n3004), .B0(n16468), .C0(n16558), .Y(
        n16557) );
  AOI211X1 U13122 ( .A0(n18128), .A1(n961), .B0(n18129), .C0(n18130), .Y(
        n18127) );
  AOI21X1 U13123 ( .A0(n18131), .A1(n18132), .B0(n2671), .Y(n18129) );
  AOI211X1 U13124 ( .A0(n5087), .A1(n2701), .B0(n18043), .C0(n18133), .Y(
        n18132) );
  AOI211X1 U13125 ( .A0(n14663), .A1(n1115), .B0(n14664), .C0(n14665), .Y(
        n14662) );
  AOI21X1 U13126 ( .A0(n14666), .A1(n14667), .B0(n3334), .Y(n14664) );
  AOI211X1 U13127 ( .A0(n5981), .A1(n3364), .B0(n14578), .C0(n14668), .Y(
        n14667) );
  AOI211X1 U13128 ( .A0(n16238), .A1(n1045), .B0(n16239), .C0(n16240), .Y(
        n16237) );
  AOI21X1 U13129 ( .A0(n16241), .A1(n16242), .B0(n3032), .Y(n16239) );
  AOI211X1 U13130 ( .A0(n5593), .A1(n3062), .B0(n16153), .C0(n16243), .Y(
        n16242) );
  AOI211X1 U13131 ( .A0(n17813), .A1(n975), .B0(n17814), .C0(n17815), .Y(
        n17812) );
  AOI21X1 U13132 ( .A0(n17816), .A1(n17817), .B0(n2731), .Y(n17814) );
  AOI211X1 U13133 ( .A0(n5195), .A1(n2761), .B0(n17728), .C0(n17818), .Y(
        n17817) );
  AOI211X1 U13134 ( .A0(n14348), .A1(n1129), .B0(n14349), .C0(n14350), .Y(
        n14347) );
  AOI21X1 U13135 ( .A0(n14351), .A1(n14352), .B0(n3392), .Y(n14349) );
  AOI211X1 U13136 ( .A0(n6057), .A1(n3422), .B0(n14263), .C0(n14353), .Y(
        n14352) );
  AOI211X1 U13137 ( .A0(n15923), .A1(n1059), .B0(n15924), .C0(n15925), .Y(
        n15922) );
  AOI21X1 U13138 ( .A0(n15926), .A1(n15927), .B0(n3093), .Y(n15924) );
  AOI211X1 U13139 ( .A0(n5669), .A1(n3123), .B0(n15838), .C0(n15928), .Y(
        n15927) );
  AOI211X1 U13140 ( .A0(n17498), .A1(n989), .B0(n17499), .C0(n17500), .Y(
        n17497) );
  AOI21X1 U13141 ( .A0(n17501), .A1(n17502), .B0(n2792), .Y(n17499) );
  AOI211X1 U13142 ( .A0(n5273), .A1(n2822), .B0(n17413), .C0(n17503), .Y(
        n17502) );
  AOI211X1 U13143 ( .A0(n5333), .A1(n5341), .B0(n10155), .C0(n10156), .Y(
        n10154) );
  AOI211X1 U13144 ( .A0(n6119), .A1(n6137), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n341), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n342), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n340) );
  AOI211X1 U13145 ( .A0(n5805), .A1(n5813), .B0(n8403), .C0(n8404), .Y(n8402)
         );
  AOI211X1 U13146 ( .A0(n4979), .A1(n4987), .B0(n11323), .C0(n11324), .Y(
        n11322) );
  AOI211X1 U13147 ( .A0(n5063), .A1(n5071), .B0(n11031), .C0(n11032), .Y(
        n11030) );
  AOI211X1 U13148 ( .A0(n6033), .A1(n6041), .B0(n7527), .C0(n7528), .Y(n7526)
         );
  AOI211X1 U13149 ( .A0(n5569), .A1(n5577), .B0(n9279), .C0(n9280), .Y(n9278)
         );
  AOI211X1 U13150 ( .A0(n5249), .A1(n5257), .B0(n10447), .C0(n10448), .Y(
        n10446) );
  AOI211X1 U13151 ( .A0(n5493), .A1(n5501), .B0(n9571), .C0(n9572), .Y(n9570)
         );
  AOI211X1 U13152 ( .A0(n5721), .A1(n5729), .B0(n8695), .C0(n8696), .Y(n8694)
         );
  AOI211X1 U13153 ( .A0(n5957), .A1(n5965), .B0(n7819), .C0(n7820), .Y(n7818)
         );
  AOI211X1 U13154 ( .A0(n4863), .A1(n4871), .B0(n11615), .C0(n11616), .Y(
        n11614) );
  AOI211X1 U13155 ( .A0(n5171), .A1(n5179), .B0(n10739), .C0(n10740), .Y(
        n10738) );
  AOI211X1 U13156 ( .A0(n5417), .A1(n5425), .B0(n9863), .C0(n9864), .Y(n9862)
         );
  AOI211X1 U13157 ( .A0(n5645), .A1(n5653), .B0(n8987), .C0(n8988), .Y(n8986)
         );
  AOI211X1 U13158 ( .A0(n5881), .A1(n5889), .B0(n8111), .C0(n8112), .Y(n8110)
         );
  AOI211X1 U13159 ( .A0(n17060), .A1(n2882), .B0(n994), .C0(n17020), .Y(n17156) );
  AOI211X1 U13160 ( .A0(n13910), .A1(n3483), .B0(n1133), .C0(n13870), .Y(
        n14006) );
  AOI211X1 U13161 ( .A0(n18320), .A1(n2640), .B0(n938), .C0(n18280), .Y(n18416) );
  AOI211X1 U13162 ( .A0(n15170), .A1(n3242), .B0(n1078), .C0(n15130), .Y(
        n15266) );
  AOI211X1 U13163 ( .A0(n15485), .A1(n3181), .B0(n1064), .C0(n15445), .Y(
        n15581) );
  AOI211X1 U13164 ( .A0(n18635), .A1(n2579), .B0(n924), .C0(n18595), .Y(n18731) );
  AOI211X1 U13165 ( .A0(n16745), .A1(n2943), .B0(n1008), .C0(n16705), .Y(
        n16841) );
  AOI211X1 U13166 ( .A0(n14855), .A1(n3303), .B0(n1092), .C0(n14815), .Y(
        n14951) );
  AOI211X1 U13167 ( .A0(n16430), .A1(n3004), .B0(n1022), .C0(n16390), .Y(
        n16526) );
  AOI211X1 U13168 ( .A0(n18005), .A1(n2701), .B0(n952), .C0(n17965), .Y(n18101) );
  AOI211X1 U13169 ( .A0(n14540), .A1(n3364), .B0(n1106), .C0(n14500), .Y(
        n14636) );
  AOI211X1 U13170 ( .A0(n16115), .A1(n3062), .B0(n1036), .C0(n16075), .Y(
        n16211) );
  AOI211X1 U13171 ( .A0(n17690), .A1(n2761), .B0(n966), .C0(n17650), .Y(n17786) );
  AOI211X1 U13172 ( .A0(n14225), .A1(n3422), .B0(n1120), .C0(n14185), .Y(
        n14321) );
  AOI211X1 U13173 ( .A0(n15800), .A1(n3123), .B0(n1050), .C0(n15760), .Y(
        n15896) );
  AOI211X1 U13174 ( .A0(n17375), .A1(n2822), .B0(n980), .C0(n17335), .Y(n17471) );
  INVX1 U13175 ( .A(n17076), .Y(n5354) );
  OAI211XL U13176 ( .A0(n106), .A1(n2882), .B0(n17077), .C0(n17026), .Y(n17076) );
  INVX1 U13177 ( .A(n13926), .Y(n6122) );
  OAI211XL U13178 ( .A0(n107), .A1(n3483), .B0(n13927), .C0(n13876), .Y(n13926) );
  INVX1 U13179 ( .A(n18336), .Y(n5000) );
  OAI211XL U13180 ( .A0(n108), .A1(n2640), .B0(n18337), .C0(n18286), .Y(n18336) );
  INVX1 U13181 ( .A(n15186), .Y(n5826) );
  OAI211XL U13182 ( .A0(n109), .A1(n3242), .B0(n15187), .C0(n15136), .Y(n15186) );
  INVX1 U13183 ( .A(n15501), .Y(n5742) );
  OAI211XL U13184 ( .A0(n110), .A1(n3181), .B0(n15502), .C0(n15451), .Y(n15501) );
  INVX1 U13185 ( .A(n18651), .Y(n4884) );
  OAI211XL U13186 ( .A0(n111), .A1(n2579), .B0(n18652), .C0(n18601), .Y(n18651) );
  INVX1 U13187 ( .A(n16761), .Y(n5438) );
  OAI211XL U13188 ( .A0(n112), .A1(n2943), .B0(n16762), .C0(n16711), .Y(n16761) );
  INVX1 U13189 ( .A(n14871), .Y(n5902) );
  OAI211XL U13190 ( .A0(n113), .A1(n3303), .B0(n14872), .C0(n14821), .Y(n14871) );
  INVX1 U13191 ( .A(n16446), .Y(n5514) );
  OAI211XL U13192 ( .A0(n114), .A1(n3004), .B0(n16447), .C0(n16396), .Y(n16446) );
  INVX1 U13193 ( .A(n18021), .Y(n5084) );
  OAI211XL U13194 ( .A0(n115), .A1(n2701), .B0(n18022), .C0(n17971), .Y(n18021) );
  INVX1 U13195 ( .A(n14556), .Y(n5978) );
  OAI211XL U13196 ( .A0(n116), .A1(n3364), .B0(n14557), .C0(n14506), .Y(n14556) );
  INVX1 U13197 ( .A(n16131), .Y(n5590) );
  OAI211XL U13198 ( .A0(n117), .A1(n3062), .B0(n16132), .C0(n16081), .Y(n16131) );
  INVX1 U13199 ( .A(n17706), .Y(n5192) );
  OAI211XL U13200 ( .A0(n118), .A1(n2761), .B0(n17707), .C0(n17656), .Y(n17706) );
  INVX1 U13201 ( .A(n14241), .Y(n6054) );
  OAI211XL U13202 ( .A0(n119), .A1(n3422), .B0(n14242), .C0(n14191), .Y(n14241) );
  INVX1 U13203 ( .A(n15816), .Y(n5666) );
  OAI211XL U13204 ( .A0(n120), .A1(n3123), .B0(n15817), .C0(n15766), .Y(n15816) );
  INVX1 U13205 ( .A(n17391), .Y(n5270) );
  OAI211XL U13206 ( .A0(n121), .A1(n2822), .B0(n17392), .C0(n17341), .Y(n17391) );
  AND2X2 U13207 ( .A(n1767), .B(n1760), .Y(n601) );
  INVX1 U13208 ( .A(n11672), .Y(n6903) );
  INVX1 U13209 ( .A(top_core_KE_sb1_n97), .Y(n6857) );
  INVX1 U13210 ( .A(n12303), .Y(n6610) );
  INVX1 U13211 ( .A(n13249), .Y(n6538) );
  INVX1 U13212 ( .A(n11988), .Y(n6563) );
  INVX1 U13213 ( .A(n12619), .Y(n6833) );
  INVX1 U13214 ( .A(n13564), .Y(n6586) );
  INVX1 U13215 ( .A(n12934), .Y(n6879) );
  AND2X2 U13216 ( .A(n1687), .B(n1681), .Y(n602) );
  AND2X2 U13217 ( .A(n1745), .B(n1739), .Y(n603) );
  AND2X2 U13218 ( .A(n1716), .B(n1710), .Y(n604) );
  AND2X2 U13219 ( .A(n1809), .B(n1802), .Y(n605) );
  AND2X2 U13220 ( .A(n1830), .B(n1823), .Y(n606) );
  AND2X2 U13221 ( .A(n1767), .B(n1760), .Y(n607) );
  AND2X2 U13222 ( .A(n1788), .B(n1781), .Y(n608) );
  AND2X2 U13223 ( .A(n1658), .B(n1651), .Y(n609) );
  AND2X2 U13224 ( .A(n1687), .B(n1681), .Y(n610) );
  AND2X2 U13225 ( .A(n1745), .B(n1739), .Y(n611) );
  AND2X2 U13226 ( .A(n1716), .B(n1710), .Y(n612) );
  AND2X2 U13227 ( .A(n1809), .B(n1802), .Y(n613) );
  AND2X2 U13228 ( .A(n1830), .B(n1823), .Y(n614) );
  AND2X2 U13229 ( .A(n1788), .B(n1781), .Y(n615) );
  AND2X2 U13230 ( .A(n1658), .B(n1651), .Y(n616) );
  CLKINVX3 U13231 ( .A(n3987), .Y(n3984) );
  INVX1 U13232 ( .A(n11728), .Y(n6827) );
  INVX1 U13233 ( .A(top_core_KE_sb1_n155), .Y(n6805) );
  INVX1 U13234 ( .A(n12359), .Y(n6531) );
  INVX1 U13235 ( .A(n13305), .Y(n6473) );
  INVX1 U13236 ( .A(n12044), .Y(n6508) );
  INVX1 U13237 ( .A(n12675), .Y(n6776) );
  INVX1 U13238 ( .A(n13620), .Y(n6520) );
  INVX1 U13239 ( .A(n12990), .Y(n6816) );
  INVX1 U13240 ( .A(n11875), .Y(n6828) );
  INVX1 U13241 ( .A(top_core_KE_sb1_n304), .Y(n6806) );
  INVX1 U13242 ( .A(n12506), .Y(n6532) );
  INVX1 U13243 ( .A(n12191), .Y(n6509) );
  INVX1 U13244 ( .A(n13766), .Y(n6521) );
  INVX1 U13245 ( .A(n13451), .Y(n6474) );
  INVX1 U13246 ( .A(n12821), .Y(n6777) );
  INVX1 U13247 ( .A(n13136), .Y(n6817) );
  INVX1 U13248 ( .A(n3955), .Y(n3920) );
  INVX1 U13249 ( .A(n3956), .Y(n3919) );
  INVX1 U13250 ( .A(n3956), .Y(n3917) );
  INVX1 U13251 ( .A(n3956), .Y(n3918) );
  INVX1 U13252 ( .A(n3954), .Y(n3925) );
  INVX1 U13253 ( .A(n3953), .Y(n3927) );
  INVX1 U13254 ( .A(n3953), .Y(n3926) );
  INVX1 U13255 ( .A(n3955), .Y(n3922) );
  INVX1 U13256 ( .A(n3954), .Y(n3924) );
  INVX1 U13257 ( .A(n3954), .Y(n3923) );
  INVX1 U13258 ( .A(n3955), .Y(n3921) );
  INVX1 U13259 ( .A(top_core_clk_slow), .Y(n3910) );
  INVX1 U13260 ( .A(n3959), .Y(n3912) );
  INVX1 U13261 ( .A(n3959), .Y(n3911) );
  INVX1 U13262 ( .A(n3949), .Y(n3908) );
  INVX1 U13263 ( .A(top_core_clk_slow), .Y(n3909) );
  INVX1 U13264 ( .A(n3958), .Y(n3914) );
  INVX1 U13265 ( .A(n3958), .Y(n3916) );
  INVX1 U13266 ( .A(n3958), .Y(n3915) );
  INVX1 U13267 ( .A(n3959), .Y(n3913) );
  INVX1 U13268 ( .A(n3957), .Y(n3942) );
  INVX1 U13269 ( .A(n3952), .Y(n3943) );
  INVX1 U13270 ( .A(n3957), .Y(n3941) );
  INVX1 U13271 ( .A(n3948), .Y(n3946) );
  INVX1 U13272 ( .A(n3948), .Y(n3944) );
  INVX1 U13273 ( .A(n3948), .Y(n3945) );
  INVX1 U13274 ( .A(n3951), .Y(n3932) );
  INVX1 U13275 ( .A(n3953), .Y(n3929) );
  INVX1 U13276 ( .A(n3956), .Y(n3931) );
  INVX1 U13277 ( .A(n3955), .Y(n3930) );
  INVX1 U13278 ( .A(n3949), .Y(n3938) );
  INVX1 U13279 ( .A(n3949), .Y(n3940) );
  INVX1 U13280 ( .A(n3949), .Y(n3939) );
  INVX1 U13281 ( .A(n3951), .Y(n3934) );
  INVX1 U13282 ( .A(n3950), .Y(n3936) );
  INVX1 U13283 ( .A(n3950), .Y(n3937) );
  INVX1 U13284 ( .A(n3950), .Y(n3935) );
  INVX1 U13285 ( .A(n3951), .Y(n3933) );
  INVX1 U13286 ( .A(n3953), .Y(n3928) );
  INVX1 U13287 ( .A(n2539), .Y(n2395) );
  INVX1 U13288 ( .A(n2521), .Y(n2397) );
  INVX1 U13289 ( .A(n2521), .Y(n2399) );
  INVX1 U13290 ( .A(n2521), .Y(n2398) );
  INVX1 U13291 ( .A(n2538), .Y(n2396) );
  INVX1 U13292 ( .A(n2852), .Y(n2854) );
  INVX1 U13293 ( .A(n3453), .Y(n3455) );
  INVX1 U13294 ( .A(n2622), .Y(n2612) );
  INVX1 U13295 ( .A(n3212), .Y(n3214) );
  INVX1 U13296 ( .A(n3151), .Y(n3153) );
  INVX1 U13297 ( .A(n2549), .Y(n2551) );
  INVX1 U13298 ( .A(n2913), .Y(n2915) );
  INVX1 U13299 ( .A(n3273), .Y(n3275) );
  INVX1 U13300 ( .A(n2974), .Y(n2976) );
  INVX1 U13301 ( .A(n3346), .Y(n3336) );
  INVX1 U13302 ( .A(n2731), .Y(n2733) );
  INVX1 U13303 ( .A(n3093), .Y(n3095) );
  INVX1 U13304 ( .A(n2792), .Y(n2794) );
  INVX1 U13305 ( .A(n2671), .Y(n2673) );
  INVX1 U13306 ( .A(n3044), .Y(n3034) );
  INVX1 U13307 ( .A(n3404), .Y(n3394) );
  INVX1 U13308 ( .A(n2285), .Y(n2297) );
  INVX1 U13309 ( .A(n2305), .Y(n2300) );
  INVX1 U13310 ( .A(n2285), .Y(n2295) );
  INVX1 U13311 ( .A(n2285), .Y(n2299) );
  INVX1 U13312 ( .A(n2289), .Y(n2294) );
  INVX1 U13313 ( .A(n2305), .Y(n2301) );
  INVX1 U13314 ( .A(n2285), .Y(n2298) );
  INVX1 U13315 ( .A(n2285), .Y(n2296) );
  INVX1 U13316 ( .A(n2289), .Y(n2293) );
  INVX1 U13317 ( .A(n2204), .Y(n2212) );
  INVX1 U13318 ( .A(n2204), .Y(n2213) );
  INVX1 U13319 ( .A(n2204), .Y(n2214) );
  INVX1 U13320 ( .A(top_core_KE_n915), .Y(n2215) );
  INVX1 U13321 ( .A(n2210), .Y(n2216) );
  INVX1 U13322 ( .A(top_core_KE_n915), .Y(n2217) );
  INVX1 U13323 ( .A(n2204), .Y(n2218) );
  INVX1 U13324 ( .A(top_core_KE_n914), .Y(n2197) );
  INVX1 U13325 ( .A(n2190), .Y(n2198) );
  INVX1 U13326 ( .A(top_core_KE_n914), .Y(n2199) );
  INVX1 U13327 ( .A(top_core_KE_n914), .Y(n2200) );
  INVX1 U13328 ( .A(n2191), .Y(n2201) );
  INVX1 U13329 ( .A(n2193), .Y(n2202) );
  INVX1 U13330 ( .A(top_core_KE_n914), .Y(n2203) );
  INVX1 U13331 ( .A(top_core_KE_n914), .Y(n2196) );
  INVX1 U13332 ( .A(top_core_EC_ss_in[86]), .Y(n2848) );
  INVX1 U13333 ( .A(top_core_EC_ss_in[6]), .Y(n3449) );
  INVX1 U13334 ( .A(top_core_EC_ss_in[118]), .Y(n2606) );
  INVX1 U13335 ( .A(top_core_EC_ss_in[38]), .Y(n3208) );
  INVX1 U13336 ( .A(top_core_EC_ss_in[46]), .Y(n3147) );
  INVX1 U13337 ( .A(top_core_EC_ss_in[126]), .Y(n2545) );
  INVX1 U13338 ( .A(top_core_EC_ss_in[78]), .Y(n2909) );
  INVX1 U13339 ( .A(top_core_EC_ss_in[70]), .Y(n2970) );
  INVX1 U13340 ( .A(top_core_EC_ss_in[110]), .Y(n2667) );
  INVX1 U13341 ( .A(top_core_EC_ss_in[22]), .Y(n3330) );
  INVX1 U13342 ( .A(top_core_EC_ss_in[62]), .Y(n3028) );
  INVX1 U13343 ( .A(top_core_EC_ss_in[102]), .Y(n2727) );
  INVX1 U13344 ( .A(top_core_EC_ss_in[14]), .Y(n3388) );
  INVX1 U13345 ( .A(top_core_EC_ss_in[54]), .Y(n3089) );
  INVX1 U13346 ( .A(top_core_EC_ss_in[94]), .Y(n2788) );
  INVX1 U13347 ( .A(top_core_EC_ss_in[30]), .Y(n3269) );
  INVX1 U13348 ( .A(n3480), .Y(n3474) );
  INVX1 U13349 ( .A(n2879), .Y(n2873) );
  INVX1 U13350 ( .A(n3480), .Y(n3475) );
  INVX1 U13351 ( .A(n2637), .Y(n2631) );
  INVX1 U13352 ( .A(n3239), .Y(n3234) );
  INVX1 U13353 ( .A(n3178), .Y(n3173) );
  INVX1 U13354 ( .A(n2576), .Y(n2570) );
  INVX1 U13355 ( .A(n2940), .Y(n2934) );
  INVX1 U13356 ( .A(n2698), .Y(n2692) );
  INVX1 U13357 ( .A(n3059), .Y(n3053) );
  INVX1 U13358 ( .A(n3419), .Y(n3413) );
  INVX1 U13359 ( .A(n3001), .Y(n2995) );
  INVX1 U13360 ( .A(n3361), .Y(n3356) );
  INVX1 U13361 ( .A(n2758), .Y(n2753) );
  INVX1 U13362 ( .A(n3120), .Y(n3114) );
  INVX1 U13363 ( .A(n3300), .Y(n3294) );
  INVX1 U13364 ( .A(n2819), .Y(n2813) );
  INVX1 U13365 ( .A(n3448), .Y(n3450) );
  INVX1 U13366 ( .A(n2847), .Y(n2849) );
  INVX1 U13367 ( .A(n2605), .Y(n2607) );
  INVX1 U13368 ( .A(n3207), .Y(n3209) );
  INVX1 U13369 ( .A(n3146), .Y(n3148) );
  INVX1 U13370 ( .A(n2544), .Y(n2546) );
  INVX1 U13371 ( .A(n2908), .Y(n2910) );
  INVX1 U13372 ( .A(n2666), .Y(n2668) );
  INVX1 U13373 ( .A(n3027), .Y(n3029) );
  INVX1 U13374 ( .A(n3387), .Y(n3389) );
  INVX1 U13375 ( .A(n2969), .Y(n2971) );
  INVX1 U13376 ( .A(n3329), .Y(n3331) );
  INVX1 U13377 ( .A(n2726), .Y(n2728) );
  INVX1 U13378 ( .A(n3088), .Y(n3090) );
  INVX1 U13379 ( .A(n2787), .Y(n2789) );
  INVX1 U13380 ( .A(n3268), .Y(n3270) );
  INVX1 U13381 ( .A(n3480), .Y(n3476) );
  INVX1 U13382 ( .A(n2879), .Y(n2874) );
  INVX1 U13383 ( .A(n2637), .Y(n2632) );
  INVX1 U13384 ( .A(n3239), .Y(n3235) );
  INVX1 U13385 ( .A(n3178), .Y(n3174) );
  INVX1 U13386 ( .A(n2576), .Y(n2571) );
  INVX1 U13387 ( .A(n2940), .Y(n2935) );
  INVX1 U13388 ( .A(n3001), .Y(n2996) );
  INVX1 U13389 ( .A(n2698), .Y(n2693) );
  INVX1 U13390 ( .A(n3361), .Y(n3357) );
  INVX1 U13391 ( .A(n3059), .Y(n3054) );
  INVX1 U13392 ( .A(n2758), .Y(n2754) );
  INVX1 U13393 ( .A(n3419), .Y(n3414) );
  INVX1 U13394 ( .A(n3120), .Y(n3115) );
  INVX1 U13395 ( .A(n3300), .Y(n3295) );
  INVX1 U13396 ( .A(n2819), .Y(n2814) );
  AND2X2 U13397 ( .A(n6305), .B(n2490), .Y(n617) );
  INVX1 U13398 ( .A(n3506), .Y(n3505) );
  INVX1 U13399 ( .A(n3492), .Y(n3490) );
  INVX1 U13400 ( .A(n3495), .Y(n3504) );
  INVX1 U13401 ( .A(n2905), .Y(n2902) );
  INVX1 U13402 ( .A(n2890), .Y(n2889) );
  INVX1 U13403 ( .A(n2905), .Y(n2903) );
  INVX1 U13404 ( .A(n3507), .Y(n3503) );
  INVX1 U13405 ( .A(n3265), .Y(n3262) );
  INVX1 U13406 ( .A(n2663), .Y(n2659) );
  INVX1 U13407 ( .A(n2663), .Y(n2660) );
  INVX1 U13408 ( .A(n3265), .Y(n3263) );
  INVX1 U13409 ( .A(n3086), .Y(n3083) );
  INVX1 U13410 ( .A(n2664), .Y(n2661) );
  INVX1 U13411 ( .A(n2648), .Y(n2647) );
  INVX1 U13412 ( .A(n3250), .Y(n3249) );
  INVX1 U13413 ( .A(n3204), .Y(n3201) );
  INVX1 U13414 ( .A(n2723), .Y(n2721) );
  INVX1 U13415 ( .A(n2723), .Y(n2720) );
  INVX1 U13416 ( .A(n3085), .Y(n3081) );
  INVX1 U13417 ( .A(n2966), .Y(n2963) );
  INVX1 U13418 ( .A(n3445), .Y(n3443) );
  INVX1 U13419 ( .A(n3445), .Y(n3442) );
  INVX1 U13420 ( .A(n2845), .Y(n2844) );
  INVX1 U13421 ( .A(n3085), .Y(n3082) );
  INVX1 U13422 ( .A(n2603), .Y(n2600) );
  INVX1 U13423 ( .A(n2602), .Y(n2599) );
  INVX1 U13424 ( .A(n3430), .Y(n3429) );
  INVX1 U13425 ( .A(n3327), .Y(n3326) );
  INVX1 U13426 ( .A(n3012), .Y(n3011) );
  INVX1 U13427 ( .A(n3190), .Y(n3189) );
  INVX1 U13428 ( .A(n3373), .Y(n3372) );
  INVX1 U13429 ( .A(n2588), .Y(n2587) );
  INVX1 U13430 ( .A(n2602), .Y(n2598) );
  INVX1 U13431 ( .A(n2785), .Y(n2784) );
  INVX1 U13432 ( .A(n2770), .Y(n2769) );
  INVX1 U13433 ( .A(n2774), .Y(n2783) );
  INVX1 U13434 ( .A(n3132), .Y(n3131) );
  INVX1 U13435 ( .A(n3311), .Y(n3310) );
  INVX1 U13436 ( .A(n3315), .Y(n3324) );
  INVX1 U13437 ( .A(n3204), .Y(n3202) );
  INVX1 U13438 ( .A(n3070), .Y(n3069) );
  INVX1 U13439 ( .A(n2966), .Y(n2964) );
  INVX1 U13440 ( .A(n2951), .Y(n2950) );
  INVX1 U13441 ( .A(n3327), .Y(n3325) );
  INVX1 U13442 ( .A(n2830), .Y(n2829) );
  INVX1 U13443 ( .A(n2366), .Y(n2494) );
  INVX1 U13444 ( .A(n2525), .Y(n2516) );
  INVX1 U13445 ( .A(n2522), .Y(n2520) );
  INVX1 U13446 ( .A(n2525), .Y(n2515) );
  INVX1 U13447 ( .A(n2524), .Y(n2517) );
  INVX1 U13448 ( .A(n2522), .Y(n2519) );
  INVX1 U13449 ( .A(n2524), .Y(n2518) );
  INVX1 U13450 ( .A(n2534), .Y(n2496) );
  INVX1 U13451 ( .A(n2540), .Y(n2514) );
  INVX1 U13452 ( .A(n2534), .Y(n2495) );
  INVX1 U13453 ( .A(top_core_EC_ss_in[6]), .Y(n3451) );
  INVX1 U13454 ( .A(top_core_EC_ss_in[86]), .Y(n2850) );
  INVX1 U13455 ( .A(top_core_EC_ss_in[118]), .Y(n2608) );
  INVX1 U13456 ( .A(top_core_EC_ss_in[38]), .Y(n3210) );
  INVX1 U13457 ( .A(top_core_EC_ss_in[110]), .Y(n2669) );
  INVX1 U13458 ( .A(top_core_EC_ss_in[62]), .Y(n3030) );
  INVX1 U13459 ( .A(top_core_EC_ss_in[14]), .Y(n3390) );
  INVX1 U13460 ( .A(top_core_EC_ss_in[70]), .Y(n2972) );
  INVX1 U13461 ( .A(top_core_EC_ss_in[46]), .Y(n3149) );
  INVX1 U13462 ( .A(top_core_EC_ss_in[22]), .Y(n3332) );
  INVX1 U13463 ( .A(top_core_EC_ss_in[126]), .Y(n2547) );
  INVX1 U13464 ( .A(top_core_EC_ss_in[102]), .Y(n2729) );
  INVX1 U13465 ( .A(top_core_EC_ss_in[78]), .Y(n2911) );
  INVX1 U13466 ( .A(top_core_EC_ss_in[54]), .Y(n3091) );
  INVX1 U13467 ( .A(top_core_EC_ss_in[94]), .Y(n2790) );
  INVX1 U13468 ( .A(top_core_EC_ss_in[30]), .Y(n3271) );
  INVX1 U13469 ( .A(n3680), .Y(n3672) );
  INVX1 U13470 ( .A(n3680), .Y(n3671) );
  INVX1 U13471 ( .A(n3680), .Y(n3670) );
  INVX1 U13472 ( .A(n3681), .Y(n3669) );
  INVX1 U13473 ( .A(n3681), .Y(n3668) );
  INVX1 U13474 ( .A(n3681), .Y(n3667) );
  INVX1 U13475 ( .A(top_core_c_ready), .Y(n3666) );
  INVX1 U13476 ( .A(n3682), .Y(n3665) );
  INVX1 U13477 ( .A(n3682), .Y(n3664) );
  INVX1 U13478 ( .A(n3682), .Y(n3663) );
  INVX1 U13479 ( .A(n3683), .Y(n3662) );
  INVX1 U13480 ( .A(n3683), .Y(n3661) );
  INVX1 U13481 ( .A(n3683), .Y(n3660) );
  INVX1 U13482 ( .A(n3684), .Y(n3659) );
  INVX1 U13483 ( .A(n3684), .Y(n3658) );
  INVX1 U13484 ( .A(n3684), .Y(n3657) );
  INVX1 U13485 ( .A(n3647), .Y(n3656) );
  INVX1 U13486 ( .A(n3648), .Y(n3655) );
  INVX1 U13487 ( .A(n3685), .Y(n3654) );
  INVX1 U13488 ( .A(n3685), .Y(n3653) );
  INVX1 U13489 ( .A(n3685), .Y(n3652) );
  INVX1 U13490 ( .A(n3627), .Y(n3626) );
  INVX1 U13491 ( .A(top_core_EC_ss_in[4]), .Y(n3469) );
  INVX1 U13492 ( .A(top_core_EC_ss_in[84]), .Y(n2868) );
  INVX1 U13493 ( .A(top_core_EC_ss_in[4]), .Y(n3470) );
  INVX1 U13494 ( .A(top_core_EC_ss_in[116]), .Y(n2626) );
  INVX1 U13495 ( .A(top_core_EC_ss_in[36]), .Y(n3228) );
  INVX1 U13496 ( .A(top_core_EC_ss_in[44]), .Y(n3167) );
  INVX1 U13497 ( .A(n2686), .Y(n2687) );
  INVX1 U13498 ( .A(top_core_EC_ss_in[76]), .Y(n2929) );
  INVX1 U13499 ( .A(top_core_EC_ss_in[124]), .Y(n2565) );
  INVX1 U13500 ( .A(top_core_EC_ss_in[28]), .Y(n3289) );
  INVX1 U13501 ( .A(top_core_EC_ss_in[68]), .Y(n2990) );
  INVX1 U13502 ( .A(top_core_EC_ss_in[20]), .Y(n3350) );
  INVX1 U13503 ( .A(top_core_EC_ss_in[60]), .Y(n3048) );
  INVX1 U13504 ( .A(top_core_EC_ss_in[100]), .Y(n2747) );
  INVX1 U13505 ( .A(top_core_EC_ss_in[12]), .Y(n3408) );
  INVX1 U13506 ( .A(top_core_EC_ss_in[52]), .Y(n3109) );
  INVX1 U13507 ( .A(top_core_EC_ss_in[92]), .Y(n2808) );
  INVX1 U13508 ( .A(top_core_EC_ss_in[100]), .Y(n2748) );
  INVX1 U13509 ( .A(n3454), .Y(n3464) );
  INVX1 U13510 ( .A(n2853), .Y(n2863) );
  INVX1 U13511 ( .A(n3213), .Y(n3223) );
  INVX1 U13512 ( .A(n2609), .Y(n2621) );
  INVX1 U13513 ( .A(n3152), .Y(n3162) );
  INVX1 U13514 ( .A(n2914), .Y(n2924) );
  INVX1 U13515 ( .A(n2562), .Y(n2560) );
  INVX1 U13516 ( .A(n3274), .Y(n3284) );
  INVX1 U13517 ( .A(n2975), .Y(n2985) );
  INVX1 U13518 ( .A(n2672), .Y(n2682) );
  INVX1 U13519 ( .A(n3333), .Y(n3345) );
  INVX1 U13520 ( .A(n3031), .Y(n3043) );
  INVX1 U13521 ( .A(n2732), .Y(n2742) );
  INVX1 U13522 ( .A(n3391), .Y(n3403) );
  INVX1 U13523 ( .A(n3094), .Y(n3104) );
  INVX1 U13524 ( .A(n2793), .Y(n2803) );
  INVX1 U13525 ( .A(top_core_EC_ss_in[108]), .Y(n2688) );
  INVX1 U13526 ( .A(n3650), .Y(n3673) );
  INVX1 U13527 ( .A(top_core_EC_ss_in[81]), .Y(n2888) );
  INVX1 U13528 ( .A(n2647), .Y(n2646) );
  INVX1 U13529 ( .A(n3249), .Y(n3248) );
  INVX1 U13530 ( .A(n3189), .Y(n3188) );
  INVX1 U13531 ( .A(top_core_EC_ss_in[105]), .Y(n2708) );
  INVX1 U13532 ( .A(n2587), .Y(n2586) );
  INVX1 U13533 ( .A(top_core_EC_ss_in[57]), .Y(n3068) );
  INVX1 U13534 ( .A(top_core_EC_ss_in[73]), .Y(n2949) );
  INVX1 U13535 ( .A(n3429), .Y(n3428) );
  INVX1 U13536 ( .A(n3310), .Y(n3309) );
  INVX1 U13537 ( .A(n3011), .Y(n3010) );
  INVX1 U13538 ( .A(n3372), .Y(n3371) );
  INVX1 U13539 ( .A(n2769), .Y(n2768) );
  INVX1 U13540 ( .A(n3131), .Y(n3130) );
  INVX1 U13541 ( .A(top_core_EC_ss_in[89]), .Y(n2828) );
  INVX1 U13542 ( .A(top_core_EC_ss_in[1]), .Y(n3489) );
  INVX1 U13543 ( .A(top_core_Addr[1]), .Y(n4022) );
  INVX1 U13544 ( .A(n4030), .Y(n4025) );
  INVX1 U13545 ( .A(n3988), .Y(n4024) );
  INVX1 U13546 ( .A(n4029), .Y(n4023) );
  INVX1 U13547 ( .A(n3988), .Y(n4021) );
  INVX1 U13548 ( .A(top_core_EC_ss_in[85]), .Y(n2864) );
  INVX1 U13549 ( .A(top_core_EC_ss_in[37]), .Y(n3224) );
  INVX1 U13550 ( .A(top_core_EC_ss_in[117]), .Y(n2622) );
  INVX1 U13551 ( .A(n3988), .Y(n4026) );
  INVX1 U13552 ( .A(n4029), .Y(n4027) );
  INVX1 U13553 ( .A(top_core_EC_ss_in[5]), .Y(n3465) );
  INVX1 U13554 ( .A(n2620), .Y(n2623) );
  INVX1 U13555 ( .A(top_core_EC_ss_in[109]), .Y(n2683) );
  INVX1 U13556 ( .A(top_core_EC_ss_in[45]), .Y(n3163) );
  INVX1 U13557 ( .A(top_core_EC_ss_in[61]), .Y(n3044) );
  INVX1 U13558 ( .A(top_core_EC_ss_in[13]), .Y(n3404) );
  INVX1 U13559 ( .A(top_core_EC_ss_in[77]), .Y(n2925) );
  INVX1 U13560 ( .A(n2379), .Y(n2527) );
  INVX1 U13561 ( .A(top_core_EC_ss_in[29]), .Y(n3285) );
  INVX1 U13562 ( .A(top_core_EC_ss_in[69]), .Y(n2986) );
  INVX1 U13563 ( .A(top_core_EC_ss_in[21]), .Y(n3346) );
  INVX1 U13564 ( .A(top_core_EC_ss_in[101]), .Y(n2743) );
  INVX1 U13565 ( .A(top_core_EC_ss_in[53]), .Y(n3105) );
  INVX1 U13566 ( .A(top_core_EC_ss_in[93]), .Y(n2804) );
  INVX1 U13567 ( .A(n3042), .Y(n3045) );
  INVX1 U13568 ( .A(n2560), .Y(n2561) );
  INVX1 U13569 ( .A(n2536), .Y(n2530) );
  INVX1 U13570 ( .A(n3402), .Y(n3405) );
  INVX1 U13571 ( .A(n2365), .Y(n2526) );
  INVX1 U13572 ( .A(n3344), .Y(n3347) );
  INVX1 U13573 ( .A(n2537), .Y(n2528) );
  INVX1 U13574 ( .A(n2537), .Y(n2529) );
  INVX1 U13575 ( .A(n2535), .Y(n2532) );
  INVX1 U13576 ( .A(n2536), .Y(n2531) );
  INVX1 U13577 ( .A(top_core_KE_n915), .Y(n2211) );
  INVX1 U13578 ( .A(n2535), .Y(n2533) );
  INVX1 U13579 ( .A(n2355), .Y(n2364) );
  INVX1 U13580 ( .A(n767), .Y(n2363) );
  INVX1 U13581 ( .A(n2315), .Y(n2316) );
  INVX1 U13582 ( .A(top_core_KE_n2179), .Y(n2325) );
  INVX1 U13583 ( .A(top_core_KE_n2179), .Y(n2326) );
  INVX1 U13584 ( .A(top_core_EC_n733), .Y(n3542) );
  INVX1 U13585 ( .A(n3650), .Y(n3674) );
  INVX1 U13586 ( .A(n3651), .Y(n3675) );
  INVX1 U13587 ( .A(n3679), .Y(n3676) );
  INVX1 U13588 ( .A(n3679), .Y(n3677) );
  INVX1 U13589 ( .A(n3679), .Y(n3678) );
  INVX1 U13590 ( .A(n1841), .Y(n1856) );
  INVX1 U13591 ( .A(n1840), .Y(n1855) );
  INVX1 U13592 ( .A(top_core_KE_n873), .Y(n1876) );
  INVX1 U13593 ( .A(top_core_KE_n743), .Y(n1854) );
  INVX1 U13594 ( .A(top_core_KE_n876), .Y(n1916) );
  INVX1 U13595 ( .A(top_core_KE_n879), .Y(n1956) );
  INVX1 U13596 ( .A(top_core_KE_n881), .Y(n1996) );
  INVX1 U13597 ( .A(top_core_KE_n888), .Y(n2076) );
  INVX1 U13598 ( .A(top_core_KE_n890), .Y(n2116) );
  INVX1 U13599 ( .A(top_core_KE_n873), .Y(n1873) );
  INVX1 U13600 ( .A(n1844), .Y(n1853) );
  INVX1 U13601 ( .A(n1899), .Y(n1913) );
  INVX1 U13602 ( .A(n1939), .Y(n1953) );
  INVX1 U13603 ( .A(n1979), .Y(n1993) );
  INVX1 U13604 ( .A(n2059), .Y(n2073) );
  INVX1 U13605 ( .A(n2099), .Y(n2113) );
  INVX1 U13606 ( .A(n1898), .Y(n1915) );
  INVX1 U13607 ( .A(n1947), .Y(n1955) );
  INVX1 U13608 ( .A(n1977), .Y(n1995) );
  INVX1 U13609 ( .A(n2057), .Y(n2075) );
  INVX1 U13610 ( .A(n2097), .Y(n2115) );
  INVX1 U13611 ( .A(top_core_KE_n873), .Y(n1874) );
  INVX1 U13612 ( .A(top_core_KE_n873), .Y(n1875) );
  INVX1 U13613 ( .A(top_core_KE_n876), .Y(n1914) );
  INVX1 U13614 ( .A(top_core_KE_n879), .Y(n1954) );
  INVX1 U13615 ( .A(top_core_KE_n881), .Y(n1994) );
  INVX1 U13616 ( .A(top_core_KE_n888), .Y(n2074) );
  INVX1 U13617 ( .A(top_core_KE_n890), .Y(n2114) );
  INVX1 U13618 ( .A(top_core_KE_n885), .Y(n2036) );
  INVX1 U13619 ( .A(n2019), .Y(n2033) );
  INVX1 U13620 ( .A(n2027), .Y(n2035) );
  INVX1 U13621 ( .A(top_core_KE_n885), .Y(n2034) );
  INVX1 U13622 ( .A(top_core_EC_ss_in[84]), .Y(n2869) );
  INVX1 U13623 ( .A(top_core_EC_ss_in[116]), .Y(n2627) );
  INVX1 U13624 ( .A(top_core_EC_ss_in[36]), .Y(n3229) );
  INVX1 U13625 ( .A(top_core_EC_ss_in[44]), .Y(n3168) );
  INVX1 U13626 ( .A(top_core_EC_ss_in[76]), .Y(n2930) );
  INVX1 U13627 ( .A(top_core_EC_ss_in[124]), .Y(n2566) );
  INVX1 U13628 ( .A(top_core_EC_ss_in[28]), .Y(n3290) );
  INVX1 U13629 ( .A(top_core_EC_ss_in[68]), .Y(n2991) );
  INVX1 U13630 ( .A(top_core_EC_ss_in[20]), .Y(n3351) );
  INVX1 U13631 ( .A(top_core_EC_ss_in[60]), .Y(n3049) );
  INVX1 U13632 ( .A(top_core_EC_ss_in[100]), .Y(n2749) );
  INVX1 U13633 ( .A(top_core_EC_ss_in[12]), .Y(n3409) );
  INVX1 U13634 ( .A(top_core_EC_ss_in[52]), .Y(n3110) );
  INVX1 U13635 ( .A(top_core_EC_ss_in[92]), .Y(n2809) );
  INVX1 U13636 ( .A(n4097), .Y(n4091) );
  INVX1 U13637 ( .A(n4105), .Y(n4073) );
  INVX1 U13638 ( .A(n4096), .Y(n4094) );
  INVX1 U13639 ( .A(n4102), .Y(n4079) );
  INVX1 U13640 ( .A(n4107), .Y(n4068) );
  INVX1 U13641 ( .A(n4097), .Y(n4090) );
  INVX1 U13642 ( .A(n4106), .Y(n4072) );
  INVX1 U13643 ( .A(n4100), .Y(n4082) );
  INVX1 U13644 ( .A(n4099), .Y(n4083) );
  INVX1 U13645 ( .A(n4101), .Y(n4087) );
  INVX1 U13646 ( .A(n4096), .Y(n4095) );
  INVX1 U13647 ( .A(n4109), .Y(n4089) );
  INVX1 U13648 ( .A(n4106), .Y(n4071) );
  INVX1 U13649 ( .A(n4098), .Y(n4086) );
  INVX1 U13650 ( .A(n4105), .Y(n4075) );
  INVX1 U13651 ( .A(n4103), .Y(n4078) );
  INVX1 U13652 ( .A(n4100), .Y(n4067) );
  INVX1 U13653 ( .A(n4096), .Y(n4093) );
  INVX1 U13654 ( .A(n4098), .Y(n4085) );
  INVX1 U13655 ( .A(n4103), .Y(n4077) );
  INVX1 U13656 ( .A(n4108), .Y(n4066) );
  INVX1 U13657 ( .A(n4031), .Y(n4088) );
  INVX1 U13658 ( .A(n4106), .Y(n4070) );
  INVX1 U13659 ( .A(n4102), .Y(n4081) );
  INVX1 U13660 ( .A(n4107), .Y(n4069) );
  INVX1 U13661 ( .A(n4105), .Y(n4074) );
  INVX1 U13662 ( .A(n4098), .Y(n4084) );
  INVX1 U13663 ( .A(n4103), .Y(n4076) );
  INVX1 U13664 ( .A(n4097), .Y(n4092) );
  INVX1 U13665 ( .A(n4102), .Y(n4080) );
  INVX1 U13666 ( .A(n2204), .Y(n2219) );
  NOR2X1 U13667 ( .A(n4128), .B(n4124), .Y(top_core_io_n188) );
  INVX1 U13668 ( .A(top_core_io_n177), .Y(n4194) );
  CLKINVX3 U13669 ( .A(n_DIN[0]), .Y(n1578) );
  CLKINVX3 U13670 ( .A(n_DIN[0]), .Y(n1579) );
  CLKINVX3 U13671 ( .A(n_DIN[0]), .Y(n1580) );
  OAI22X2 U13672 ( .A0(n2461), .A1(top_core_EC_ss_n226), .B0(n2368), .B1(n5042), .Y(top_core_EC_mc_mix_in_8[15]) );
  OAI22X2 U13673 ( .A0(n2432), .A1(top_core_EC_ss_n191), .B0(n2370), .B1(n5394), .Y(top_core_EC_mc_mix_in_8[47]) );
  OAI22X2 U13674 ( .A0(n2423), .A1(top_core_EC_ss_n214), .B0(n2369), .B1(n5309), .Y(top_core_EC_mc_mix_in_2_16_) );
  OAI22X2 U13675 ( .A0(n2430), .A1(top_core_EC_ss_n197), .B0(n2370), .B1(n5781), .Y(top_core_EC_mc_mix_in_2_32_) );
  OAI22X2 U13676 ( .A0(n2406), .A1(top_core_EC_ss_n212), .B0(n2369), .B1(n4850), .Y(top_core_EC_mc_mix_in_2_26_) );
  OAI22X2 U13677 ( .A0(n2437), .A1(top_core_EC_ss_n177), .B0(n2371), .B1(n5232), .Y(top_core_EC_mc_mix_in_2_58_) );
  NOR2X2 U13678 ( .A(n1676), .B(n1666), .Y(n13229) );
  NOR2X2 U13679 ( .A(n1705), .B(n1695), .Y(n12914) );
  NOR2X2 U13680 ( .A(n1734), .B(n1724), .Y(n12599) );
  OAI22X2 U13681 ( .A0(n2522), .A1(top_core_EC_ss_n130), .B0(n2375), .B1(n5046), .Y(top_core_EC_mc_mix_in_2_10_) );
  OAI22X2 U13682 ( .A0(n2431), .A1(top_core_EC_ss_n194), .B0(n2370), .B1(n5404), .Y(top_core_EC_mc_mix_in_2_42_) );
  OAI22X2 U13683 ( .A0(n2434), .A1(top_core_EC_ss_n185), .B0(n2371), .B1(n6094), .Y(top_core_EC_mc_mix_in_8[7]) );
  OAI22X2 U13684 ( .A0(n2435), .A1(top_core_EC_ss_n182), .B0(n2371), .B1(n4958), .Y(top_core_EC_mc_mix_in_8[55]) );
  OAI22X2 U13685 ( .A0(n2429), .A1(top_core_EC_ss_n200), .B0(n2370), .B1(n5784), .Y(top_core_EC_mc_mix_in_8[39]) );
  OAI22X2 U13686 ( .A0(n2425), .A1(top_core_EC_ss_n217), .B0(n2368), .B1(n5312), .Y(top_core_EC_mc_mix_in_8[23]) );
  NOR2X2 U13687 ( .A(n17153), .B(n17167), .Y(n17205) );
  NOR2X2 U13688 ( .A(n14003), .B(n14017), .Y(n14055) );
  NOR2X2 U13689 ( .A(n18413), .B(n18427), .Y(n18465) );
  NOR2X2 U13690 ( .A(n15263), .B(n15277), .Y(n15315) );
  NOR2X2 U13691 ( .A(n15578), .B(n15592), .Y(n15630) );
  NOR2X2 U13692 ( .A(n16838), .B(n16852), .Y(n16890) );
  NOR2X2 U13693 ( .A(n18728), .B(n18742), .Y(n18780) );
  NOR2X2 U13694 ( .A(n14948), .B(n14962), .Y(n15000) );
  NOR2X2 U13695 ( .A(n16523), .B(n16537), .Y(n16575) );
  NOR2X2 U13696 ( .A(n18098), .B(n18112), .Y(n18150) );
  NOR2X2 U13697 ( .A(n14633), .B(n14647), .Y(n14685) );
  NOR2X2 U13698 ( .A(n16208), .B(n16222), .Y(n16260) );
  NOR2X2 U13699 ( .A(n17783), .B(n17797), .Y(n17835) );
  NOR2X2 U13700 ( .A(n14318), .B(n14332), .Y(n14370) );
  NOR2X2 U13701 ( .A(n15893), .B(n15907), .Y(n15945) );
  NOR2X2 U13702 ( .A(n17468), .B(n17482), .Y(n17520) );
  OAI221XL U13703 ( .A0(n1246), .A1(n9917), .B0(n2898), .B1(n9886), .C0(n9944), 
        .Y(n9902) );
  OAI221XL U13704 ( .A0(n1328), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n101), 
        .B0(n3500), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n68), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n129), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n85) );
  OAI221XL U13705 ( .A0(n1234), .A1(n8165), .B0(n3258), .B1(n8134), .C0(n8192), 
        .Y(n8150) );
  OAI221XL U13706 ( .A0(n1254), .A1(n11085), .B0(n2655), .B1(n11054), .C0(
        n11112), .Y(n11070) );
  OAI221XL U13707 ( .A0(n1252), .A1(n10793), .B0(n2716), .B1(n10762), .C0(
        n10820), .Y(n10778) );
  OAI221XL U13708 ( .A0(n1240), .A1(n9041), .B0(n3077), .B1(n9010), .C0(n9068), 
        .Y(n9026) );
  OAI221XL U13709 ( .A0(n1228), .A1(n7289), .B0(n3438), .B1(n7258), .C0(n7316), 
        .Y(n7274) );
  OAI221XL U13710 ( .A0(n1248), .A1(n10209), .B0(n2841), .B1(n10178), .C0(
        n10236), .Y(n10194) );
  OAI221XL U13711 ( .A0(n1242), .A1(n9333), .B0(n3022), .B1(n9302), .C0(n9360), 
        .Y(n9318) );
  OAI221XL U13712 ( .A0(n1236), .A1(n8457), .B0(n3197), .B1(n8426), .C0(n8484), 
        .Y(n8442) );
  OAI221XL U13713 ( .A0(n1230), .A1(n7581), .B0(n3382), .B1(n7550), .C0(n7608), 
        .Y(n7566) );
  OAI221XL U13714 ( .A0(n1256), .A1(n11377), .B0(n2594), .B1(n11346), .C0(
        n11404), .Y(n11362) );
  OAI221XL U13715 ( .A0(n1250), .A1(n10501), .B0(n2780), .B1(n10470), .C0(
        n10528), .Y(n10486) );
  OAI221XL U13716 ( .A0(n1244), .A1(n9625), .B0(n2959), .B1(n9594), .C0(n9652), 
        .Y(n9610) );
  OAI221XL U13717 ( .A0(n1238), .A1(n8749), .B0(n3141), .B1(n8718), .C0(n8776), 
        .Y(n8734) );
  OAI221XL U13718 ( .A0(n1232), .A1(n7873), .B0(n3321), .B1(n7842), .C0(n7900), 
        .Y(n7858) );
  NAND2X2 U13719 ( .A(n1666), .B(n1677), .Y(n13256) );
  NAND2X2 U13720 ( .A(n1724), .B(n1736), .Y(n12626) );
  NAND2X2 U13721 ( .A(n1695), .B(n1707), .Y(n12941) );
  NAND2X2 U13722 ( .A(n1000), .B(n2868), .Y(n9893) );
  NAND2X2 U13723 ( .A(n1140), .B(n3471), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n76) );
  NAND2X2 U13724 ( .A(n944), .B(n2626), .Y(n11061) );
  NAND2X2 U13725 ( .A(n1084), .B(n3228), .Y(n8141) );
  NAND2X2 U13726 ( .A(n958), .B(n2687), .Y(n10769) );
  NAND2X2 U13727 ( .A(n1042), .B(n3050), .Y(n9017) );
  NAND2X2 U13728 ( .A(n1126), .B(n3410), .Y(n7265) );
  NAND2X2 U13729 ( .A(n986), .B(n2808), .Y(n10185) );
  NAND2X2 U13730 ( .A(n1028), .B(n2990), .Y(n9309) );
  NAND2X2 U13731 ( .A(n1070), .B(n3167), .Y(n8433) );
  NAND2X2 U13732 ( .A(n1112), .B(n3350), .Y(n7557) );
  NAND2X2 U13733 ( .A(n930), .B(n2565), .Y(n11353) );
  NAND2X2 U13734 ( .A(n972), .B(n2748), .Y(n10477) );
  NAND2X2 U13735 ( .A(n1014), .B(n2929), .Y(n9601) );
  NAND2X2 U13736 ( .A(n1056), .B(n3109), .Y(n8725) );
  NAND2X2 U13737 ( .A(n1098), .B(n3289), .Y(n7849) );
  NAND2X2 U13738 ( .A(n1203), .B(n1211), .Y(n11852) );
  NAND2X2 U13739 ( .A(n1194), .B(n1210), .Y(top_core_KE_sb1_n281) );
  NAND2X2 U13740 ( .A(n1149), .B(n1679), .Y(n13428) );
  NAND2X2 U13741 ( .A(n1154), .B(n1170), .Y(n12168) );
  NAND2X2 U13742 ( .A(n1189), .B(n1735), .Y(n12798) );
  NAND2X2 U13743 ( .A(n1198), .B(n1706), .Y(n13113) );
  NAND2X2 U13744 ( .A(n1158), .B(n1644), .Y(n13743) );
  NAND2X2 U13745 ( .A(n6964), .B(n1795), .Y(n11674) );
  NAND2X2 U13746 ( .A(n6958), .B(n1816), .Y(top_core_KE_sb1_n99) );
  NAND2X2 U13747 ( .A(n1675), .B(n1671), .Y(n13251) );
  NAND2X2 U13748 ( .A(n6670), .B(n1774), .Y(n11990) );
  NAND2X2 U13749 ( .A(n1706), .B(n1700), .Y(n12936) );
  NAND2X2 U13750 ( .A(n1643), .B(n1635), .Y(n13566) );
  NAND2X2 U13751 ( .A(n1735), .B(n1729), .Y(n12621) );
  NOR2X1 U13752 ( .A(n17075), .B(n17035), .Y(n17068) );
  NOR2X1 U13753 ( .A(n13925), .B(n13885), .Y(n13918) );
  NOR2X1 U13754 ( .A(n18335), .B(n18295), .Y(n18328) );
  NOR2X1 U13755 ( .A(n15185), .B(n15145), .Y(n15178) );
  NOR2X1 U13756 ( .A(n15500), .B(n15460), .Y(n15493) );
  NOR2X1 U13757 ( .A(n18650), .B(n18610), .Y(n18643) );
  NOR2X1 U13758 ( .A(n16760), .B(n16720), .Y(n16753) );
  NOR2X1 U13759 ( .A(n14870), .B(n14830), .Y(n14863) );
  NOR2X1 U13760 ( .A(n16445), .B(n16405), .Y(n16438) );
  NOR2X1 U13761 ( .A(n18020), .B(n17980), .Y(n18013) );
  NOR2X1 U13762 ( .A(n14555), .B(n14515), .Y(n14548) );
  NOR2X1 U13763 ( .A(n16130), .B(n16090), .Y(n16123) );
  NOR2X1 U13764 ( .A(n17705), .B(n17665), .Y(n17698) );
  NOR2X1 U13765 ( .A(n14240), .B(n14200), .Y(n14233) );
  NOR2X1 U13766 ( .A(n15815), .B(n15775), .Y(n15808) );
  NOR2X1 U13767 ( .A(n17390), .B(n17350), .Y(n17383) );
  OAI22X1 U13768 ( .A0(n2483), .A1(top_core_EC_ss_n207), .B0(n2369), .B1(n6100), .Y(top_core_EC_mix_in[2]) );
  OAI22X1 U13769 ( .A0(n2431), .A1(top_core_EC_ss_n196), .B0(n2370), .B1(n6098), .Y(top_core_EC_mix_in[3]) );
  AOI22X1 U13770 ( .A0(n1675), .A1(n1692), .B0(n1673), .B1(n629), .Y(n13294)
         );
  AOI22X1 U13771 ( .A0(n1733), .A1(n1750), .B0(n1731), .B1(n630), .Y(n12664)
         );
  AOI22X1 U13772 ( .A0(n1704), .A1(n1721), .B0(n1702), .B1(n632), .Y(n12979)
         );
  OAI22X1 U13773 ( .A0(n2435), .A1(top_core_EC_ss_n141), .B0(n2374), .B1(n5047), .Y(top_core_EC_mix_in[8]) );
  OAI22X1 U13774 ( .A0(n2431), .A1(top_core_EC_ss_n195), .B0(n2370), .B1(n5395), .Y(top_core_EC_mix_in[40]) );
  OAI22X1 U13775 ( .A0(n2432), .A1(top_core_EC_ss_n193), .B0(n2370), .B1(n5402), .Y(top_core_EC_mix_in[42]) );
  OAI22X1 U13776 ( .A0(n2432), .A1(top_core_EC_ss_n192), .B0(n2370), .B1(n5401), .Y(top_core_EC_mix_in[43]) );
  OAI22X1 U13777 ( .A0(n2435), .A1(top_core_EC_ss_n184), .B0(n2371), .B1(n4962), .Y(top_core_EC_mix_in[50]) );
  OAI22X1 U13778 ( .A0(n2404), .A1(top_core_EC_ss_n222), .B0(n2368), .B1(n5314), .Y(top_core_EC_mix_in[16]) );
  OAI22X1 U13779 ( .A0(n2434), .A1(top_core_EC_ss_n187), .B0(n2371), .B1(n4960), .Y(top_core_EC_mix_in[48]) );
  OAI22X1 U13780 ( .A0(n2435), .A1(top_core_EC_ss_n183), .B0(n2371), .B1(n4959), .Y(top_core_EC_mix_in[51]) );
  OAI22X1 U13781 ( .A0(n2402), .A1(top_core_EC_ss_n220), .B0(n2368), .B1(n5316), .Y(top_core_EC_mix_in[18]) );
  OAI22X1 U13782 ( .A0(n2400), .A1(top_core_EC_ss_n202), .B0(n2370), .B1(n5788), .Y(top_core_EC_mix_in[34]) );
  OAI22X1 U13783 ( .A0(n2481), .A1(top_core_EC_ss_n257), .B0(n2370), .B1(n6095), .Y(top_core_EC_mix_in[0]) );
  OAI22X1 U13784 ( .A0(n2476), .A1(top_core_EC_ss_n219), .B0(n2368), .B1(n5313), .Y(top_core_EC_mix_in[19]) );
  OAI22X1 U13785 ( .A0(n2436), .A1(top_core_EC_ss_n204), .B0(n2369), .B1(n5786), .Y(top_core_EC_mix_in[32]) );
  OAI22X1 U13786 ( .A0(n2429), .A1(top_core_EC_ss_n201), .B0(n2370), .B1(n5785), .Y(top_core_EC_mix_in[35]) );
  OAI22X1 U13787 ( .A0(n2426), .A1(top_core_EC_ss_n246), .B0(n2367), .B1(n5045), .Y(top_core_EC_mix_in[10]) );
  OAI22X1 U13788 ( .A0(n2529), .A1(top_core_EC_ss_n235), .B0(n2368), .B1(n5043), .Y(top_core_EC_mix_in[11]) );
  NOR2X1 U13789 ( .A(n1000), .B(n2873), .Y(n17167) );
  NOR2X1 U13790 ( .A(n1140), .B(n3475), .Y(n14017) );
  NOR2X1 U13791 ( .A(n944), .B(n2631), .Y(n18427) );
  NOR2X1 U13792 ( .A(n1084), .B(n3234), .Y(n15277) );
  NOR2X1 U13793 ( .A(n1070), .B(n3173), .Y(n15592) );
  NOR2X1 U13794 ( .A(n1014), .B(n2934), .Y(n16852) );
  NOR2X1 U13795 ( .A(n930), .B(n2570), .Y(n18742) );
  NOR2X1 U13796 ( .A(n1098), .B(n3294), .Y(n14962) );
  NOR2X1 U13797 ( .A(n1028), .B(n2995), .Y(n16537) );
  NOR2X1 U13798 ( .A(n958), .B(n2692), .Y(n18112) );
  NOR2X1 U13799 ( .A(n1112), .B(n3356), .Y(n14647) );
  NOR2X1 U13800 ( .A(n1042), .B(n3053), .Y(n16222) );
  NOR2X1 U13801 ( .A(n972), .B(n2753), .Y(n17797) );
  NOR2X1 U13802 ( .A(n1126), .B(n3413), .Y(n14332) );
  NOR2X1 U13803 ( .A(n1056), .B(n3114), .Y(n15907) );
  NOR2X1 U13804 ( .A(n986), .B(n2813), .Y(n17482) );
  NAND2X1 U13805 ( .A(n681), .B(n745), .Y(n11808) );
  NAND2X1 U13806 ( .A(n682), .B(n746), .Y(top_core_KE_sb1_n236) );
  NAND2X1 U13807 ( .A(n683), .B(n744), .Y(n12439) );
  NAND2X1 U13808 ( .A(n684), .B(n747), .Y(n12124) );
  NOR2X1 U13809 ( .A(n12483), .B(n1266), .Y(n12372) );
  NOR2X1 U13810 ( .A(n2871), .B(n1000), .Y(n17060) );
  NOR2X1 U13811 ( .A(n3472), .B(n1140), .Y(n13910) );
  NOR2X1 U13812 ( .A(n2629), .B(n944), .Y(n18320) );
  NOR2X1 U13813 ( .A(n3231), .B(n1084), .Y(n15170) );
  NOR2X1 U13814 ( .A(n3292), .B(n1098), .Y(n14855) );
  NOR2X1 U13815 ( .A(n2993), .B(n1028), .Y(n16430) );
  NOR2X1 U13816 ( .A(n2690), .B(n958), .Y(n18005) );
  NOR2X1 U13817 ( .A(n3353), .B(n1112), .Y(n14540) );
  NOR2X1 U13818 ( .A(n3051), .B(n1042), .Y(n16115) );
  NOR2X1 U13819 ( .A(n2750), .B(n972), .Y(n17690) );
  NOR2X1 U13820 ( .A(n3411), .B(n1126), .Y(n14225) );
  NOR2X1 U13821 ( .A(n3112), .B(n1056), .Y(n15800) );
  NOR2X1 U13822 ( .A(n2811), .B(n986), .Y(n17375) );
  NOR2X1 U13823 ( .A(n3170), .B(n1070), .Y(n15485) );
  NOR2X1 U13824 ( .A(n2568), .B(n930), .Y(n18635) );
  NOR2X1 U13825 ( .A(n2932), .B(n1014), .Y(n16745) );
  NOR2X1 U13826 ( .A(n13597), .B(n183), .Y(n13573) );
  NOR2X1 U13827 ( .A(n6), .B(n685), .Y(n13556) );
  NAND2X1 U13828 ( .A(n761), .B(n1211), .Y(n11706) );
  NAND2X1 U13829 ( .A(n762), .B(n1210), .Y(top_core_KE_sb1_n131) );
  NAND2X1 U13830 ( .A(n756), .B(n1676), .Y(n13283) );
  NAND2X1 U13831 ( .A(n763), .B(n1170), .Y(n12022) );
  NAND2X1 U13832 ( .A(n757), .B(n1735), .Y(n12653) );
  NAND2X1 U13833 ( .A(n759), .B(n1643), .Y(n13598) );
  NAND2X1 U13834 ( .A(n758), .B(n1706), .Y(n12968) );
  NOR2BX1 U13835 ( .AN(n13858), .B(n1140), .Y(n14033) );
  NOR2BX1 U13836 ( .AN(n17008), .B(n1000), .Y(n17183) );
  NOR2BX1 U13837 ( .AN(n18268), .B(n944), .Y(n18443) );
  NOR2BX1 U13838 ( .AN(n15118), .B(n1084), .Y(n15293) );
  NOR2BX1 U13839 ( .AN(n15433), .B(n1070), .Y(n15608) );
  NOR2BX1 U13840 ( .AN(n16693), .B(n1014), .Y(n16868) );
  NOR2BX1 U13841 ( .AN(n18583), .B(n930), .Y(n18758) );
  NOR2BX1 U13842 ( .AN(n14803), .B(n1098), .Y(n14978) );
  NOR2BX1 U13843 ( .AN(n16378), .B(n1028), .Y(n16553) );
  NOR2BX1 U13844 ( .AN(n17953), .B(n958), .Y(n18128) );
  NOR2BX1 U13845 ( .AN(n14488), .B(n1112), .Y(n14663) );
  NOR2BX1 U13846 ( .AN(n16063), .B(n1042), .Y(n16238) );
  NOR2BX1 U13847 ( .AN(n17638), .B(n972), .Y(n17813) );
  NOR2BX1 U13848 ( .AN(n14173), .B(n1126), .Y(n14348) );
  NOR2BX1 U13849 ( .AN(n15748), .B(n1056), .Y(n15923) );
  NOR2BX1 U13850 ( .AN(n17323), .B(n986), .Y(n17498) );
  NOR3XL U13851 ( .A(n13256), .B(n1174), .C(n52), .Y(n13230) );
  NOR3XL U13852 ( .A(n11679), .B(n605), .C(n50), .Y(n11653) );
  NOR3XL U13853 ( .A(top_core_KE_sb1_n104), .B(n606), .C(n51), .Y(
        top_core_KE_sb1_n78) );
  NOR3XL U13854 ( .A(n12310), .B(n607), .C(n89), .Y(n12285) );
  NOR3XL U13855 ( .A(n11995), .B(n608), .C(n53), .Y(n11969) );
  NOR3XL U13856 ( .A(n12626), .B(n1214), .C(n54), .Y(n12600) );
  NOR3XL U13857 ( .A(n13571), .B(n1179), .C(n55), .Y(n13545) );
  NOR3XL U13858 ( .A(n12941), .B(n1220), .C(n56), .Y(n12915) );
  AOI22X1 U13859 ( .A0(top_core_EC_ss_sbox_out_r[84]), .A1(n2462), .B0(
        top_core_EC_ss_sbox_out[84]), .B1(n2380), .Y(top_core_EC_ss_n217) );
  OAI21XL U13860 ( .A0(n17138), .A1(n992), .B0(n17139), .Y(
        top_core_EC_ss_sbox_out[84]) );
  OAI222XL U13861 ( .A0(n10022), .A1(n9932), .B0(n10023), .B1(n9934), .C0(
        n10024), .C1(n992), .Y(top_core_EC_ss_sbox_out_r[84]) );
  AOI222X1 U13862 ( .A0(n2847), .A1(n17157), .B0(n5321), .B1(n17158), .C0(
        n17051), .C1(n17159), .Y(n17138) );
  AOI22X1 U13863 ( .A0(top_core_EC_ss_sbox_out_r[4]), .A1(n2446), .B0(
        top_core_EC_ss_sbox_out[4]), .B1(n2497), .Y(top_core_EC_ss_n185) );
  OAI21XL U13864 ( .A0(n13988), .A1(n1132), .B0(n13989), .Y(
        top_core_EC_ss_sbox_out[4]) );
  OAI222XL U13865 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n208), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n117), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n209), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n119), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n210), .C1(n1132), .Y(
        top_core_EC_ss_sbox_out_r[4]) );
  AOI222X1 U13866 ( .A0(n3448), .A1(n14007), .B0(n6105), .B1(n14008), .C0(
        n13901), .C1(n14009), .Y(n13988) );
  AOI22X1 U13867 ( .A0(top_core_EC_ss_sbox_out_r[116]), .A1(n2447), .B0(
        top_core_EC_ss_sbox_out[116]), .B1(n2384), .Y(top_core_EC_ss_n182) );
  OAI21XL U13868 ( .A0(n18398), .A1(n936), .B0(n18399), .Y(
        top_core_EC_ss_sbox_out[116]) );
  OAI222XL U13869 ( .A0(n11190), .A1(n11100), .B0(n11191), .B1(n11102), .C0(
        n11192), .C1(n936), .Y(top_core_EC_ss_sbox_out_r[116]) );
  AOI222X1 U13870 ( .A0(n2605), .A1(n18417), .B0(n4967), .B1(n18418), .C0(
        n18311), .C1(n18419), .Y(n18398) );
  AOI22X1 U13871 ( .A0(top_core_EC_ss_sbox_out_r[36]), .A1(n2442), .B0(
        top_core_EC_ss_sbox_out[36]), .B1(n2370), .Y(top_core_EC_ss_n200) );
  OAI21XL U13872 ( .A0(n15248), .A1(n1076), .B0(n15249), .Y(
        top_core_EC_ss_sbox_out[36]) );
  OAI222XL U13873 ( .A0(n8270), .A1(n8180), .B0(n8271), .B1(n8182), .C0(n8272), 
        .C1(n1076), .Y(top_core_EC_ss_sbox_out_r[36]) );
  AOI222X1 U13874 ( .A0(n3207), .A1(n15267), .B0(n5793), .B1(n15268), .C0(
        n15161), .C1(n15269), .Y(n15248) );
  AOI22X1 U13875 ( .A0(top_core_EC_ss_sbox_out_r[108]), .A1(n2465), .B0(
        top_core_EC_ss_sbox_out[44]), .B1(n2368), .Y(top_core_EC_ss_n226) );
  OAI21XL U13876 ( .A0(n15563), .A1(n1062), .B0(n15564), .Y(
        top_core_EC_ss_sbox_out[44]) );
  OAI222XL U13877 ( .A0(n10898), .A1(n10808), .B0(n10899), .B1(n10810), .C0(
        n10900), .C1(n950), .Y(top_core_EC_ss_sbox_out_r[108]) );
  AOI222X1 U13878 ( .A0(n3146), .A1(n15582), .B0(n5709), .B1(n15583), .C0(
        n15476), .C1(n15584), .Y(n15563) );
  AOI22X1 U13879 ( .A0(top_core_EC_ss_sbox_out_r[60]), .A1(n2397), .B0(
        top_core_EC_ss_sbox_out[124]), .B1(n2514), .Y(top_core_EC_ss_n209) );
  OAI21XL U13880 ( .A0(n18713), .A1(n922), .B0(n18714), .Y(
        top_core_EC_ss_sbox_out[124]) );
  OAI222XL U13881 ( .A0(n9146), .A1(n9056), .B0(n9147), .B1(n9058), .C0(n9148), 
        .C1(n1034), .Y(top_core_EC_ss_sbox_out_r[60]) );
  AOI222X1 U13882 ( .A0(n2544), .A1(n18732), .B0(n4851), .B1(n18733), .C0(
        n18626), .C1(n18734), .Y(n18713) );
  AOI22X1 U13883 ( .A0(top_core_EC_ss_sbox_out_r[12]), .A1(n2523), .B0(
        top_core_EC_ss_sbox_out[76]), .B1(n2539), .Y(top_core_EC_ss_n191) );
  OAI21XL U13884 ( .A0(n16823), .A1(n1006), .B0(n16824), .Y(
        top_core_EC_ss_sbox_out[76]) );
  OAI222XL U13885 ( .A0(n7394), .A1(n7304), .B0(n7395), .B1(n7306), .C0(n7396), 
        .C1(n1118), .Y(top_core_EC_ss_sbox_out_r[12]) );
  AOI222X1 U13886 ( .A0(n2908), .A1(n16842), .B0(n5405), .B1(n16843), .C0(
        n16736), .C1(n16844), .Y(n16823) );
  AOI22X1 U13887 ( .A0(top_core_EC_ss_sbox_out_r[92]), .A1(n2532), .B0(
        top_core_EC_ss_sbox_out[28]), .B1(n2517), .Y(top_core_EC_ss_n173) );
  OAI21XL U13888 ( .A0(n14933), .A1(n1090), .B0(n14934), .Y(
        top_core_EC_ss_sbox_out[28]) );
  OAI222XL U13889 ( .A0(n10314), .A1(n10224), .B0(n10315), .B1(n10226), .C0(
        n10316), .C1(n978), .Y(top_core_EC_ss_sbox_out_r[92]) );
  AOI222X1 U13890 ( .A0(n3268), .A1(n14952), .B0(n5869), .B1(n14953), .C0(
        n14846), .C1(n14954), .Y(n14933) );
  AOI22X1 U13891 ( .A0(top_core_EC_ss_sbox_out_r[68]), .A1(n2450), .B0(
        top_core_EC_ss_sbox_out[68]), .B1(n2504), .Y(top_core_EC_ss_n165) );
  OAI21XL U13892 ( .A0(n16508), .A1(n1020), .B0(n16509), .Y(
        top_core_EC_ss_sbox_out[68]) );
  OAI222XL U13893 ( .A0(n9438), .A1(n9348), .B0(n9439), .B1(n9350), .C0(n9440), 
        .C1(n1020), .Y(top_core_EC_ss_sbox_out_r[68]) );
  AOI222X1 U13894 ( .A0(n2969), .A1(n16527), .B0(n5481), .B1(n16528), .C0(
        n16421), .C1(n16529), .Y(n16508) );
  AOI22X1 U13895 ( .A0(top_core_EC_ss_sbox_out_r[44]), .A1(n2453), .B0(
        top_core_EC_ss_sbox_out[108]), .B1(n2501), .Y(top_core_EC_ss_n156) );
  OAI21XL U13896 ( .A0(n18083), .A1(n950), .B0(n18084), .Y(
        top_core_EC_ss_sbox_out[108]) );
  OAI222XL U13897 ( .A0(n8562), .A1(n8472), .B0(n8563), .B1(n8474), .C0(n8564), 
        .C1(n1062), .Y(top_core_EC_ss_sbox_out_r[44]) );
  AOI222X1 U13898 ( .A0(n2666), .A1(n18102), .B0(n5051), .B1(n18103), .C0(
        n17996), .C1(n18104), .Y(n18083) );
  AOI22X1 U13899 ( .A0(top_core_EC_ss_sbox_out_r[20]), .A1(n2456), .B0(
        top_core_EC_ss_sbox_out[20]), .B1(n2394), .Y(top_core_EC_ss_n147) );
  OAI21XL U13900 ( .A0(n14618), .A1(n1104), .B0(n14619), .Y(
        top_core_EC_ss_sbox_out[20]) );
  OAI222XL U13901 ( .A0(n7686), .A1(n7596), .B0(n7687), .B1(n7598), .C0(n7688), 
        .C1(n1104), .Y(top_core_EC_ss_sbox_out_r[20]) );
  AOI222X1 U13902 ( .A0(n3329), .A1(n14637), .B0(n5945), .B1(n14638), .C0(
        n14531), .C1(n14639), .Y(n14618) );
  AOI22X1 U13903 ( .A0(top_core_EC_ss_sbox_out_r[124]), .A1(n2459), .B0(
        top_core_EC_ss_sbox_out[60]), .B1(n2394), .Y(top_core_EC_ss_n138) );
  OAI21XL U13904 ( .A0(n16193), .A1(n1034), .B0(n16194), .Y(
        top_core_EC_ss_sbox_out[60]) );
  OAI222XL U13905 ( .A0(n11482), .A1(n11392), .B0(n11483), .B1(n11394), .C0(
        n11484), .C1(n922), .Y(top_core_EC_ss_sbox_out_r[124]) );
  AOI222X1 U13906 ( .A0(n3027), .A1(n16212), .B0(n5557), .B1(n16213), .C0(
        n16106), .C1(n16214), .Y(n16193) );
  AOI22X1 U13907 ( .A0(top_core_EC_ss_sbox_out_r[100]), .A1(n2475), .B0(
        top_core_EC_ss_sbox_out[100]), .B1(n2373), .Y(top_core_EC_ss_n256) );
  OAI21XL U13908 ( .A0(n17768), .A1(n964), .B0(n17769), .Y(
        top_core_EC_ss_sbox_out[100]) );
  OAI222XL U13909 ( .A0(n10606), .A1(n10516), .B0(n10607), .B1(n10518), .C0(
        n10608), .C1(n964), .Y(top_core_EC_ss_sbox_out_r[100]) );
  AOI222X1 U13910 ( .A0(n2726), .A1(n17787), .B0(n5159), .B1(n17788), .C0(
        n17681), .C1(n17789), .Y(n17768) );
  AOI22X1 U13911 ( .A0(top_core_EC_ss_sbox_out_r[76]), .A1(n2473), .B0(
        top_core_EC_ss_sbox_out[12]), .B1(n2390), .Y(top_core_EC_ss_n248) );
  OAI21XL U13912 ( .A0(n14303), .A1(n1118), .B0(n14304), .Y(
        top_core_EC_ss_sbox_out[12]) );
  OAI222XL U13913 ( .A0(n9730), .A1(n9640), .B0(n9731), .B1(n9642), .C0(n9732), 
        .C1(n1006), .Y(top_core_EC_ss_sbox_out_r[76]) );
  AOI222X1 U13914 ( .A0(n3387), .A1(n14322), .B0(n6021), .B1(n14323), .C0(
        n14216), .C1(n14324), .Y(n14303) );
  AOI22X1 U13915 ( .A0(top_core_EC_ss_sbox_out_r[52]), .A1(n2470), .B0(
        top_core_EC_ss_sbox_out[52]), .B1(n2386), .Y(top_core_EC_ss_n239) );
  OAI21XL U13916 ( .A0(n15878), .A1(n1048), .B0(n15879), .Y(
        top_core_EC_ss_sbox_out[52]) );
  OAI222XL U13917 ( .A0(n8854), .A1(n8764), .B0(n8855), .B1(n8766), .C0(n8856), 
        .C1(n1048), .Y(top_core_EC_ss_sbox_out_r[52]) );
  AOI222X1 U13918 ( .A0(n3088), .A1(n15897), .B0(n5633), .B1(n15898), .C0(
        n15791), .C1(n15899), .Y(n15878) );
  AOI22X1 U13919 ( .A0(top_core_EC_ss_sbox_out_r[28]), .A1(n2467), .B0(
        top_core_EC_ss_sbox_out[92]), .B1(n2373), .Y(top_core_EC_ss_n230) );
  OAI21XL U13920 ( .A0(n17453), .A1(n978), .B0(n17454), .Y(
        top_core_EC_ss_sbox_out[92]) );
  OAI222XL U13921 ( .A0(n7978), .A1(n7888), .B0(n7979), .B1(n7890), .C0(n7980), 
        .C1(n1090), .Y(top_core_EC_ss_sbox_out_r[28]) );
  AOI222X1 U13922 ( .A0(n2787), .A1(n17472), .B0(n5237), .B1(n17473), .C0(
        n17366), .C1(n17474), .Y(n17453) );
  NAND2X1 U13923 ( .A(n3467), .B(n1140), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n131) );
  NAND2X1 U13924 ( .A(n2866), .B(n1000), .Y(n9946) );
  NAND2X1 U13925 ( .A(n2624), .B(n944), .Y(n11114) );
  NAND2X1 U13926 ( .A(n3226), .B(n1084), .Y(n8194) );
  NAND2X1 U13927 ( .A(n2685), .B(n958), .Y(n10822) );
  NAND2X1 U13928 ( .A(n3046), .B(n1042), .Y(n9070) );
  NAND2X1 U13929 ( .A(n3406), .B(n1126), .Y(n7318) );
  NAND2X1 U13930 ( .A(n2806), .B(n986), .Y(n10238) );
  NAND2X1 U13931 ( .A(n2988), .B(n1028), .Y(n9362) );
  NAND2X1 U13932 ( .A(n3165), .B(n1070), .Y(n8486) );
  NAND2X1 U13933 ( .A(n3348), .B(n1112), .Y(n7610) );
  NAND2X1 U13934 ( .A(n2563), .B(n930), .Y(n11406) );
  NAND2X1 U13935 ( .A(n2745), .B(n972), .Y(n10530) );
  NAND2X1 U13936 ( .A(n2927), .B(n1014), .Y(n9654) );
  NAND2X1 U13937 ( .A(n3107), .B(n1056), .Y(n8778) );
  NAND2X1 U13938 ( .A(n3287), .B(n1098), .Y(n7902) );
  OAI222XL U13939 ( .A0(n1222), .A1(n11677), .B0(n11678), .B1(n1796), .C0(
        n11679), .C1(n11680), .Y(n11665) );
  OAI222XL U13940 ( .A0(n1216), .A1(top_core_KE_sb1_n102), .B0(
        top_core_KE_sb1_n103), .B1(n1817), .C0(top_core_KE_sb1_n104), .C1(
        top_core_KE_sb1_n105), .Y(top_core_KE_sb1_n90) );
  OAI222XL U13941 ( .A0(n1176), .A1(n11993), .B0(n11994), .B1(n1775), .C0(
        n11995), .C1(n11996), .Y(n11981) );
  OAI222XL U13942 ( .A0(n1181), .A1(n12308), .B0(n12309), .B1(n1753), .C0(
        n12310), .C1(n12311), .Y(n12296) );
  OAI222XL U13943 ( .A0(n1178), .A1(n13569), .B0(n13570), .B1(n1636), .C0(
        n13571), .C1(n13572), .Y(n13557) );
  OAI222XL U13944 ( .A0(n1173), .A1(n13254), .B0(n13255), .B1(n1670), .C0(
        n13256), .C1(n13257), .Y(n13242) );
  OAI222XL U13945 ( .A0(n1219), .A1(n12939), .B0(n12940), .B1(n1699), .C0(
        n12941), .C1(n12942), .Y(n12927) );
  OAI222XL U13946 ( .A0(n1213), .A1(n12624), .B0(n12625), .B1(n1728), .C0(
        n12626), .C1(n12627), .Y(n12612) );
  AOI22X1 U13947 ( .A0(n1680), .A1(n1673), .B0(n1675), .B1(n629), .Y(n13313)
         );
  AOI22X1 U13948 ( .A0(n1738), .A1(n1731), .B0(n1733), .B1(n630), .Y(n12683)
         );
  AOI22X1 U13949 ( .A0(n1709), .A1(n1702), .B0(n1704), .B1(n632), .Y(n12998)
         );
  XOR2X1 U13950 ( .A(n1536), .B(top_core_EC_mix_in[74]), .Y(
        top_core_EC_mc_mix_in_2_75_) );
  XOR2X1 U13951 ( .A(n1554), .B(top_core_EC_mix_in[106]), .Y(
        top_core_EC_mc_mix_in_2_107_) );
  OAI222XL U13952 ( .A0(n17075), .A1(n17074), .B0(n17208), .B1(n2900), .C0(n57), .C1(n17007), .Y(n17206) );
  OAI222XL U13953 ( .A0(n13925), .A1(n13924), .B0(n14058), .B1(n3501), .C0(n58), .C1(n13857), .Y(n14056) );
  OAI222XL U13954 ( .A0(n18335), .A1(n18334), .B0(n18468), .B1(n2657), .C0(n59), .C1(n18267), .Y(n18466) );
  OAI222XL U13955 ( .A0(n15185), .A1(n15184), .B0(n15318), .B1(n3260), .C0(n60), .C1(n15117), .Y(n15316) );
  OAI222XL U13956 ( .A0(n15500), .A1(n15499), .B0(n15633), .B1(n3199), .C0(n61), .C1(n15432), .Y(n15631) );
  OAI222XL U13957 ( .A0(n16760), .A1(n16759), .B0(n16893), .B1(n2961), .C0(n62), .C1(n16692), .Y(n16891) );
  OAI222XL U13958 ( .A0(n18650), .A1(n18649), .B0(n18783), .B1(n2596), .C0(n63), .C1(n18582), .Y(n18781) );
  OAI222XL U13959 ( .A0(n14870), .A1(n14869), .B0(n15003), .B1(n3323), .C0(n64), .C1(n14802), .Y(n15001) );
  OAI222XL U13960 ( .A0(n16445), .A1(n16444), .B0(n16578), .B1(n3021), .C0(n65), .C1(n16377), .Y(n16576) );
  OAI222XL U13961 ( .A0(n18020), .A1(n18019), .B0(n18153), .B1(n2718), .C0(n66), .C1(n17952), .Y(n18151) );
  OAI222XL U13962 ( .A0(n14555), .A1(n14554), .B0(n14688), .B1(n3381), .C0(n67), .C1(n14487), .Y(n14686) );
  OAI222XL U13963 ( .A0(n16130), .A1(n16129), .B0(n16263), .B1(n3079), .C0(n68), .C1(n16062), .Y(n16261) );
  OAI222XL U13964 ( .A0(n17705), .A1(n17704), .B0(n17838), .B1(n2781), .C0(n69), .C1(n17637), .Y(n17836) );
  OAI222XL U13965 ( .A0(n14240), .A1(n14239), .B0(n14373), .B1(n3440), .C0(n70), .C1(n14172), .Y(n14371) );
  OAI222XL U13966 ( .A0(n15815), .A1(n15814), .B0(n15948), .B1(n3140), .C0(n71), .C1(n15747), .Y(n15946) );
  OAI222XL U13967 ( .A0(n17390), .A1(n17389), .B0(n17523), .B1(n2843), .C0(n72), .C1(n17322), .Y(n17521) );
  NOR2X1 U13968 ( .A(n11852), .B(n1807), .Y(n11642) );
  NOR2X1 U13969 ( .A(top_core_KE_sb1_n281), .B(n1828), .Y(top_core_KE_sb1_n67)
         );
  NOR2X1 U13970 ( .A(n12483), .B(n1762), .Y(n12274) );
  NOR2X1 U13971 ( .A(n13428), .B(n1684), .Y(n13219) );
  NOR2X1 U13972 ( .A(n12168), .B(n1786), .Y(n11958) );
  NOR2X1 U13973 ( .A(n12798), .B(n1742), .Y(n12589) );
  NOR2X1 U13974 ( .A(n13743), .B(n1654), .Y(n13534) );
  NOR2X1 U13975 ( .A(n13113), .B(n1713), .Y(n12904) );
  NOR3XL U13976 ( .A(n13312), .B(n1666), .C(n52), .Y(n13409) );
  NOR3XL U13977 ( .A(n12682), .B(n1724), .C(n54), .Y(n12779) );
  NOR3XL U13978 ( .A(n12997), .B(n1695), .C(n56), .Y(n13094) );
  OAI221XL U13979 ( .A0(n1615), .A1(n9886), .B0(n9895), .B1(n9889), .C0(n10148), .Y(n10147) );
  AOI22X1 U13980 ( .A0(n10149), .A1(n2851), .B0(n2855), .B1(n10150), .Y(n10148) );
  NAND3X1 U13981 ( .A(n10152), .B(n10013), .C(n10153), .Y(n10149) );
  OAI221XL U13982 ( .A0(n1001), .A1(n9918), .B0(n2884), .B1(n9896), .C0(n10151), .Y(n10150) );
  OAI221XL U13983 ( .A0(n1625), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n68), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n78), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n71), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n334), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n333) );
  AOI22X1 U13984 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n335), .A1(n3452), 
        .B0(n3456), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n336), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n334) );
  NAND3X1 U13985 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n338), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n199), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n339), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n335) );
  OAI221XL U13986 ( .A0(n1143), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n102), 
        .B0(n3488), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n337), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n336) );
  OAI221XL U13987 ( .A0(n1621), .A1(n8134), .B0(n8143), .B1(n8137), .C0(n8396), 
        .Y(n8395) );
  AOI22X1 U13988 ( .A0(n8397), .A1(n3211), .B0(n3215), .B1(n8398), .Y(n8396)
         );
  NAND3X1 U13989 ( .A(n8400), .B(n8261), .C(n8401), .Y(n8397) );
  OAI221XL U13990 ( .A0(n1085), .A1(n8166), .B0(n3243), .B1(n8144), .C0(n8399), 
        .Y(n8398) );
  OAI221XL U13991 ( .A0(n1611), .A1(n11054), .B0(n11063), .B1(n11057), .C0(
        n11316), .Y(n11315) );
  AOI22X1 U13992 ( .A0(n11317), .A1(n2609), .B0(n2613), .B1(n11318), .Y(n11316) );
  NAND3X1 U13993 ( .A(n11320), .B(n11181), .C(n11321), .Y(n11317) );
  OAI221XL U13994 ( .A0(n945), .A1(n11086), .B0(n2646), .B1(n11064), .C0(
        n11319), .Y(n11318) );
  OAI221XL U13995 ( .A0(n1612), .A1(n10762), .B0(n10771), .B1(n10765), .C0(
        n11024), .Y(n11023) );
  AOI22X1 U13996 ( .A0(n11025), .A1(n2670), .B0(n2674), .B1(n11026), .Y(n11024) );
  NAND3X1 U13997 ( .A(n11028), .B(n10889), .C(n11029), .Y(n11025) );
  OAI221XL U13998 ( .A0(n959), .A1(n10794), .B0(n2706), .B1(n10772), .C0(
        n11027), .Y(n11026) );
  OAI221XL U13999 ( .A0(n1624), .A1(n7258), .B0(n7267), .B1(n7261), .C0(n7520), 
        .Y(n7519) );
  AOI22X1 U14000 ( .A0(n7521), .A1(n3391), .B0(n3395), .B1(n7522), .Y(n7520)
         );
  NAND3X1 U14001 ( .A(n7524), .B(n7385), .C(n7525), .Y(n7521) );
  OAI221XL U14002 ( .A0(n1127), .A1(n7290), .B0(n3428), .B1(n7268), .C0(n7523), 
        .Y(n7522) );
  OAI221XL U14003 ( .A0(n1618), .A1(n9010), .B0(n9019), .B1(n9013), .C0(n9272), 
        .Y(n9271) );
  AOI22X1 U14004 ( .A0(n9273), .A1(n3031), .B0(n3035), .B1(n9274), .Y(n9272)
         );
  NAND3X1 U14005 ( .A(n9276), .B(n9137), .C(n9277), .Y(n9273) );
  OAI221XL U14006 ( .A0(n1043), .A1(n9042), .B0(n3064), .B1(n9020), .C0(n9275), 
        .Y(n9274) );
  OAI221XL U14007 ( .A0(n1614), .A1(n10178), .B0(n10187), .B1(n10181), .C0(
        n10440), .Y(n10439) );
  AOI22X1 U14008 ( .A0(n10441), .A1(n2791), .B0(n2795), .B1(n10442), .Y(n10440) );
  NAND3X1 U14009 ( .A(n10444), .B(n10305), .C(n10445), .Y(n10441) );
  OAI221XL U14010 ( .A0(n987), .A1(n10210), .B0(n2824), .B1(n10188), .C0(
        n10443), .Y(n10442) );
  OAI221XL U14011 ( .A0(n1617), .A1(n9302), .B0(n9311), .B1(n9305), .C0(n9564), 
        .Y(n9563) );
  AOI22X1 U14012 ( .A0(n9565), .A1(n2973), .B0(n2977), .B1(n9566), .Y(n9564)
         );
  NAND3X1 U14013 ( .A(n9568), .B(n9429), .C(n9569), .Y(n9565) );
  OAI221XL U14014 ( .A0(n1029), .A1(n9334), .B0(n3005), .B1(n9312), .C0(n9567), 
        .Y(n9566) );
  OAI221XL U14015 ( .A0(n1620), .A1(n8426), .B0(n8435), .B1(n8429), .C0(n8688), 
        .Y(n8687) );
  AOI22X1 U14016 ( .A0(n8689), .A1(n3150), .B0(n3154), .B1(n8690), .Y(n8688)
         );
  NAND3X1 U14017 ( .A(n8692), .B(n8553), .C(n8693), .Y(n8689) );
  OAI221XL U14018 ( .A0(n1071), .A1(n8458), .B0(n3186), .B1(n8436), .C0(n8691), 
        .Y(n8690) );
  OAI221XL U14019 ( .A0(n1623), .A1(n7550), .B0(n7559), .B1(n7553), .C0(n7812), 
        .Y(n7811) );
  AOI22X1 U14020 ( .A0(n7813), .A1(n3333), .B0(n3337), .B1(n7814), .Y(n7812)
         );
  NAND3X1 U14021 ( .A(n7816), .B(n7677), .C(n7817), .Y(n7813) );
  OAI221XL U14022 ( .A0(n1113), .A1(n7582), .B0(n3369), .B1(n7560), .C0(n7815), 
        .Y(n7814) );
  OAI221XL U14023 ( .A0(n1610), .A1(n11346), .B0(n11355), .B1(n11349), .C0(
        n11608), .Y(n11607) );
  AOI22X1 U14024 ( .A0(n11609), .A1(n2548), .B0(n2552), .B1(n11610), .Y(n11608) );
  NAND3X1 U14025 ( .A(n11612), .B(n11473), .C(n11613), .Y(n11609) );
  OAI221XL U14026 ( .A0(n931), .A1(n11378), .B0(n2584), .B1(n11356), .C0(
        n11611), .Y(n11610) );
  OAI221XL U14027 ( .A0(n1613), .A1(n10470), .B0(n10479), .B1(n10473), .C0(
        n10732), .Y(n10731) );
  AOI22X1 U14028 ( .A0(n10733), .A1(n2730), .B0(n2734), .B1(n10734), .Y(n10732) );
  NAND3X1 U14029 ( .A(n10736), .B(n10597), .C(n10737), .Y(n10733) );
  OAI221XL U14030 ( .A0(n973), .A1(n10502), .B0(n2766), .B1(n10480), .C0(
        n10735), .Y(n10734) );
  OAI221XL U14031 ( .A0(n1616), .A1(n9594), .B0(n9603), .B1(n9597), .C0(n9856), 
        .Y(n9855) );
  AOI22X1 U14032 ( .A0(n9857), .A1(n2912), .B0(n2916), .B1(n9858), .Y(n9856)
         );
  NAND3X1 U14033 ( .A(n9860), .B(n9721), .C(n9861), .Y(n9857) );
  OAI221XL U14034 ( .A0(n1015), .A1(n9626), .B0(n2945), .B1(n9604), .C0(n9859), 
        .Y(n9858) );
  OAI221XL U14035 ( .A0(n1619), .A1(n8718), .B0(n8727), .B1(n8721), .C0(n8980), 
        .Y(n8979) );
  AOI22X1 U14036 ( .A0(n8981), .A1(n3092), .B0(n3096), .B1(n8982), .Y(n8980)
         );
  NAND3X1 U14037 ( .A(n8984), .B(n8845), .C(n8985), .Y(n8981) );
  OAI221XL U14038 ( .A0(n1057), .A1(n8750), .B0(n3128), .B1(n8728), .C0(n8983), 
        .Y(n8982) );
  OAI221XL U14039 ( .A0(n1622), .A1(n7842), .B0(n7851), .B1(n7845), .C0(n8104), 
        .Y(n8103) );
  AOI22X1 U14040 ( .A0(n8105), .A1(n3272), .B0(n3276), .B1(n8106), .Y(n8104)
         );
  NAND3X1 U14041 ( .A(n8108), .B(n7969), .C(n8109), .Y(n8105) );
  OAI221XL U14042 ( .A0(n1099), .A1(n7874), .B0(n3304), .B1(n7852), .C0(n8107), 
        .Y(n8106) );
  NOR2X1 U14043 ( .A(n1205), .B(n6909), .Y(n11867) );
  NOR2X1 U14044 ( .A(n1196), .B(n6863), .Y(top_core_KE_sb1_n296) );
  NOR2X1 U14045 ( .A(n1165), .B(n6616), .Y(n12498) );
  NOR2X1 U14046 ( .A(n1156), .B(n6569), .Y(n12183) );
  OAI222XL U14047 ( .A0(n9893), .A1(n9913), .B0(n1615), .B1(n9886), .C0(n10032), .C1(n9900), .Y(n10167) );
  OAI222XL U14048 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n76), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .B0(n1625), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n68), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n218), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n83), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n353) );
  OAI222XL U14049 ( .A0(n8141), .A1(n8161), .B0(n1621), .B1(n8134), .C0(n8280), 
        .C1(n8148), .Y(n8415) );
  OAI222XL U14050 ( .A0(n11061), .A1(n11081), .B0(n1611), .B1(n11054), .C0(
        n11200), .C1(n11068), .Y(n11335) );
  OAI222XL U14051 ( .A0(n10769), .A1(n10789), .B0(n1612), .B1(n10762), .C0(
        n10908), .C1(n10776), .Y(n11043) );
  OAI222XL U14052 ( .A0(n7265), .A1(n7285), .B0(n1624), .B1(n7258), .C0(n7404), 
        .C1(n7272), .Y(n7539) );
  OAI222XL U14053 ( .A0(n9017), .A1(n9037), .B0(n1618), .B1(n9010), .C0(n9156), 
        .C1(n9024), .Y(n9291) );
  OAI222XL U14054 ( .A0(n10185), .A1(n10205), .B0(n1614), .B1(n10178), .C0(
        n10324), .C1(n10192), .Y(n10459) );
  OAI222XL U14055 ( .A0(n9309), .A1(n9329), .B0(n1617), .B1(n9302), .C0(n9448), 
        .C1(n9316), .Y(n9583) );
  OAI222XL U14056 ( .A0(n8433), .A1(n8453), .B0(n1620), .B1(n8426), .C0(n8572), 
        .C1(n8440), .Y(n8707) );
  OAI222XL U14057 ( .A0(n7557), .A1(n7577), .B0(n1623), .B1(n7550), .C0(n7696), 
        .C1(n7564), .Y(n7831) );
  OAI222XL U14058 ( .A0(n11353), .A1(n11373), .B0(n1610), .B1(n11346), .C0(
        n11492), .C1(n11360), .Y(n11627) );
  OAI222XL U14059 ( .A0(n10477), .A1(n10497), .B0(n1613), .B1(n10470), .C0(
        n10616), .C1(n10484), .Y(n10751) );
  OAI222XL U14060 ( .A0(n9601), .A1(n9621), .B0(n1616), .B1(n9594), .C0(n9740), 
        .C1(n9608), .Y(n9875) );
  OAI222XL U14061 ( .A0(n8725), .A1(n8745), .B0(n1619), .B1(n8718), .C0(n8864), 
        .C1(n8732), .Y(n8999) );
  OAI222XL U14062 ( .A0(n7849), .A1(n7869), .B0(n1622), .B1(n7842), .C0(n7988), 
        .C1(n7856), .Y(n8123) );
  OAI222XL U14063 ( .A0(n13388), .A1(n1665), .B0(n13389), .B1(n13256), .C0(
        n1666), .C1(n13390), .Y(n13377) );
  AOI211X1 U14064 ( .A0(n6544), .A1(n1683), .B0(n13391), .C0(n13392), .Y(
        n13390) );
  AOI221X1 U14065 ( .A0(n6552), .A1(n692), .B0(n1172), .B1(n756), .C0(n13394), 
        .Y(n13388) );
  AOI21XL U14066 ( .A0(n6550), .A1(n1274), .B0(n6538), .Y(n13389) );
  OAI222XL U14067 ( .A0(n12758), .A1(n1723), .B0(n12759), .B1(n12626), .C0(
        n1724), .C1(n12760), .Y(n12747) );
  AOI211X1 U14068 ( .A0(n6839), .A1(n1741), .B0(n12761), .C0(n12762), .Y(
        n12760) );
  AOI221X1 U14069 ( .A0(n6847), .A1(n694), .B0(n1212), .B1(n757), .C0(n12764), 
        .Y(n12758) );
  AOI21XL U14070 ( .A0(n6845), .A1(n1268), .B0(n6833), .Y(n12759) );
  OAI222XL U14071 ( .A0(n13073), .A1(n1694), .B0(n13074), .B1(n12941), .C0(
        n1695), .C1(n13075), .Y(n13062) );
  AOI211X1 U14072 ( .A0(n6885), .A1(n1712), .B0(n13076), .C0(n13077), .Y(
        n13075) );
  AOI221X1 U14073 ( .A0(n6893), .A1(n696), .B0(n1218), .B1(n758), .C0(n13079), 
        .Y(n13073) );
  AOI21XL U14074 ( .A0(n6891), .A1(n1271), .B0(n6879), .Y(n13074) );
  XOR2X1 U14075 ( .A(n1539), .B(top_core_EC_mix_in[58]), .Y(
        top_core_EC_mc_mix_in_2_59_) );
  XOR2X1 U14076 ( .A(n1533), .B(top_core_EC_mix_in[90]), .Y(
        top_core_EC_mc_mix_in_2_91_) );
  XOR2X1 U14077 ( .A(n1551), .B(top_core_EC_mix_in[122]), .Y(
        top_core_EC_mc_mix_in_2_123_) );
  OAI221XL U14078 ( .A0(n1172), .A1(n13428), .B0(n1692), .B1(n73), .C0(n13515), 
        .Y(n13514) );
  AOI22X1 U14079 ( .A0(n692), .A1(n1151), .B0(n6549), .B1(n1682), .Y(n13515)
         );
  NOR2X1 U14080 ( .A(n12290), .B(n1181), .Y(n12333) );
  OAI221XL U14081 ( .A0(n11766), .A1(n11674), .B0(n11767), .B1(n1796), .C0(
        n11768), .Y(n11754) );
  AOI211X1 U14082 ( .A0(n6909), .A1(n1803), .B0(n11770), .C0(n11771), .Y(
        n11767) );
  OAI221XL U14083 ( .A0(top_core_KE_sb1_n194), .A1(top_core_KE_sb1_n99), .B0(
        top_core_KE_sb1_n195), .B1(n1817), .C0(top_core_KE_sb1_n196), .Y(
        top_core_KE_sb1_n182) );
  AOI211X1 U14084 ( .A0(n6863), .A1(n1824), .B0(top_core_KE_sb1_n198), .C0(
        top_core_KE_sb1_n199), .Y(top_core_KE_sb1_n195) );
  OAI221XL U14085 ( .A0(n12082), .A1(n11990), .B0(n12083), .B1(n1775), .C0(
        n12084), .Y(n12070) );
  AOI211X1 U14086 ( .A0(n6569), .A1(n1782), .B0(n12086), .C0(n12087), .Y(
        n12083) );
  OAI221XL U14087 ( .A0(n12397), .A1(n12305), .B0(n12398), .B1(n1753), .C0(
        n12399), .Y(n12385) );
  AOI211X1 U14088 ( .A0(n6616), .A1(n1761), .B0(n12401), .C0(n12402), .Y(
        n12398) );
  OAI221XL U14089 ( .A0(n13658), .A1(n13566), .B0(n13659), .B1(n1636), .C0(
        n13660), .Y(n13646) );
  AOI211X1 U14090 ( .A0(n6592), .A1(n1652), .B0(n13662), .C0(n13663), .Y(
        n13659) );
  OAI221XL U14091 ( .A0(n13343), .A1(n13251), .B0(n13344), .B1(n1669), .C0(
        n13345), .Y(n13331) );
  AOI211X1 U14092 ( .A0(n6544), .A1(n1681), .B0(n13347), .C0(n13348), .Y(
        n13344) );
  OAI221XL U14093 ( .A0(n12713), .A1(n12621), .B0(n12714), .B1(n1727), .C0(
        n12715), .Y(n12701) );
  AOI211X1 U14094 ( .A0(n6839), .A1(n1739), .B0(n12717), .C0(n12718), .Y(
        n12714) );
  OAI221XL U14095 ( .A0(n13028), .A1(n12936), .B0(n13029), .B1(n1698), .C0(
        n13030), .Y(n13016) );
  AOI211X1 U14096 ( .A0(n6885), .A1(n1710), .B0(n13032), .C0(n13033), .Y(
        n13029) );
  NAND2X1 U14097 ( .A(n1205), .B(n1222), .Y(n11757) );
  NAND2X1 U14098 ( .A(n1196), .B(n1216), .Y(top_core_KE_sb1_n185) );
  NAND2X1 U14099 ( .A(n1165), .B(n1181), .Y(n12388) );
  NAND2X1 U14100 ( .A(n1156), .B(n1176), .Y(n12073) );
  NOR2X1 U14101 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n104), .B(n3489), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n112) );
  NOR2X1 U14102 ( .A(n9919), .B(n2886), .Y(n9927) );
  NOR2X1 U14103 ( .A(n11087), .B(n2648), .Y(n11095) );
  NOR2X1 U14104 ( .A(n8167), .B(n3244), .Y(n8175) );
  NOR2X1 U14105 ( .A(n10795), .B(n2702), .Y(n10803) );
  NOR2X1 U14106 ( .A(n9043), .B(n3064), .Y(n9051) );
  NOR2X1 U14107 ( .A(n7291), .B(n3430), .Y(n7299) );
  NOR2X1 U14108 ( .A(n10211), .B(n2824), .Y(n10219) );
  NOR2X1 U14109 ( .A(n9335), .B(n3006), .Y(n9343) );
  NOR2X1 U14110 ( .A(n8459), .B(n3182), .Y(n8467) );
  NOR2X1 U14111 ( .A(n7583), .B(n3365), .Y(n7591) );
  NOR2X1 U14112 ( .A(n11379), .B(n2580), .Y(n11387) );
  NOR2X1 U14113 ( .A(n10503), .B(n2762), .Y(n10511) );
  NOR2X1 U14114 ( .A(n9627), .B(n2945), .Y(n9635) );
  NOR2X1 U14115 ( .A(n8751), .B(n3124), .Y(n8759) );
  NOR2X1 U14116 ( .A(n7875), .B(n3305), .Y(n7883) );
  NAND2X1 U14117 ( .A(n1205), .B(n1809), .Y(n11734) );
  NAND2X1 U14118 ( .A(n1196), .B(n1830), .Y(top_core_KE_sb1_n161) );
  NAND2X1 U14119 ( .A(n1165), .B(n1767), .Y(n12365) );
  NAND2X1 U14120 ( .A(n1156), .B(n1788), .Y(n12050) );
  NOR2XL U14121 ( .A(n6), .B(n583), .Y(n13656) );
  CLKINVX3 U14122 ( .A(n9919), .Y(n5388) );
  CLKINVX3 U14123 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n104), .Y(n6175) );
  CLKINVX3 U14124 ( .A(n11087), .Y(n5034) );
  CLKINVX3 U14125 ( .A(n8167), .Y(n5860) );
  CLKINVX3 U14126 ( .A(n10795), .Y(n5118) );
  CLKINVX3 U14127 ( .A(n7291), .Y(n6088) );
  CLKINVX3 U14128 ( .A(n9043), .Y(n5624) );
  CLKINVX3 U14129 ( .A(n10211), .Y(n5304) );
  CLKINVX3 U14130 ( .A(n9335), .Y(n5548) );
  CLKINVX3 U14131 ( .A(n8459), .Y(n5776) );
  CLKINVX3 U14132 ( .A(n7583), .Y(n6012) );
  CLKINVX3 U14133 ( .A(n11379), .Y(n4918) );
  CLKINVX3 U14134 ( .A(n10503), .Y(n5226) );
  CLKINVX3 U14135 ( .A(n9627), .Y(n5472) );
  CLKINVX3 U14136 ( .A(n8751), .Y(n5700) );
  CLKINVX3 U14137 ( .A(n7875), .Y(n5936) );
  OAI211XL U14138 ( .A0(n52), .A1(n1681), .B0(n13297), .C0(n13247), .Y(n13296)
         );
  OAI211XL U14139 ( .A0(n54), .A1(n1739), .B0(n12667), .C0(n12617), .Y(n12666)
         );
  OAI211XL U14140 ( .A0(n56), .A1(n1710), .B0(n12982), .C0(n12932), .Y(n12981)
         );
  OAI211XL U14141 ( .A0(n55), .A1(n1652), .B0(n13612), .C0(n13562), .Y(n13611)
         );
  OAI211XL U14142 ( .A0(n89), .A1(n1761), .B0(n12351), .C0(n12301), .Y(n12350)
         );
  OAI211XL U14143 ( .A0(n50), .A1(n1803), .B0(n11720), .C0(n11670), .Y(n11719)
         );
  OAI211XL U14144 ( .A0(n51), .A1(n1824), .B0(top_core_KE_sb1_n147), .C0(
        top_core_KE_sb1_n95), .Y(top_core_KE_sb1_n146) );
  OAI211XL U14145 ( .A0(n53), .A1(n1782), .B0(n12036), .C0(n11986), .Y(n12035)
         );
  NAND2X1 U14146 ( .A(n6598), .B(n1643), .Y(n13550) );
  NAND2X1 U14147 ( .A(n6915), .B(n1211), .Y(n11658) );
  NAND2X1 U14148 ( .A(n6869), .B(n1210), .Y(top_core_KE_sb1_n83) );
  NAND2X1 U14149 ( .A(n6575), .B(n1170), .Y(n11974) );
  AOI32XL U14150 ( .A0(n17135), .A1(n2872), .A2(n1615), .B0(n17153), .B1(n1002), .Y(n17225) );
  AOI32XL U14151 ( .A0(n13985), .A1(n3473), .A2(n1625), .B0(n14003), .B1(n1141), .Y(n14075) );
  AOI32XL U14152 ( .A0(n15245), .A1(n3232), .A2(n1621), .B0(n15263), .B1(n1086), .Y(n15335) );
  AOI32XL U14153 ( .A0(n18395), .A1(n2630), .A2(n1611), .B0(n18413), .B1(n946), 
        .Y(n18485) );
  AOI32XL U14154 ( .A0(n15560), .A1(n3171), .A2(n1620), .B0(n15578), .B1(n1072), .Y(n15650) );
  AOI32XL U14155 ( .A0(n16820), .A1(n2933), .A2(n1616), .B0(n16838), .B1(n1016), .Y(n16910) );
  AOI32XL U14156 ( .A0(n18710), .A1(n2569), .A2(n1610), .B0(n18728), .B1(n932), 
        .Y(n18800) );
  AOI32XL U14157 ( .A0(n14930), .A1(n3293), .A2(n1622), .B0(n14948), .B1(n1100), .Y(n15020) );
  AOI32XL U14158 ( .A0(n16505), .A1(n2994), .A2(n1617), .B0(n16523), .B1(n1030), .Y(n16595) );
  AOI32XL U14159 ( .A0(n18080), .A1(n2691), .A2(n1612), .B0(n18098), .B1(n960), 
        .Y(n18170) );
  AOI32XL U14160 ( .A0(n14615), .A1(n3354), .A2(n1623), .B0(n14633), .B1(n1114), .Y(n14705) );
  AOI32XL U14161 ( .A0(n16190), .A1(n3052), .A2(n1618), .B0(n16208), .B1(n1044), .Y(n16280) );
  AOI32XL U14162 ( .A0(n17765), .A1(n2751), .A2(n1613), .B0(n17783), .B1(n974), 
        .Y(n17855) );
  AOI32XL U14163 ( .A0(n14300), .A1(n3412), .A2(n1624), .B0(n14318), .B1(n1128), .Y(n14390) );
  AOI32XL U14164 ( .A0(n15875), .A1(n3113), .A2(n1619), .B0(n15893), .B1(n1058), .Y(n15965) );
  AOI32XL U14165 ( .A0(n17450), .A1(n2812), .A2(n1614), .B0(n17468), .B1(n988), 
        .Y(n17540) );
  NAND2X1 U14166 ( .A(n6550), .B(n1675), .Y(n13235) );
  NAND2X1 U14167 ( .A(n6845), .B(n1733), .Y(n12605) );
  NAND2X1 U14168 ( .A(n6891), .B(n1704), .Y(n12920) );
  OAI22X1 U14169 ( .A0(top_core_EC_mc_n541), .A1(n2480), .B0(n2379), .B1(
        top_core_EC_mc_n542), .Y(top_core_EC_mix_out_34_) );
  XOR2X1 U14170 ( .A(top_core_EC_mc_n543), .B(top_core_EC_mc_n544), .Y(
        top_core_EC_mc_n542) );
  XNOR2X1 U14171 ( .A(top_core_EC_mix_in[58]), .B(top_core_EC_mc_n545), .Y(
        top_core_EC_mc_n541) );
  XNOR2X1 U14172 ( .A(top_core_EC_mix_in[58]), .B(top_core_EC_mc_n424), .Y(
        top_core_EC_mc_n543) );
  OAI22X1 U14173 ( .A0(top_core_EC_mc_n533), .A1(n2481), .B0(n2379), .B1(
        top_core_EC_mc_n534), .Y(top_core_EC_mix_out_35_) );
  XOR2X1 U14174 ( .A(top_core_EC_mc_n535), .B(top_core_EC_mc_n536), .Y(
        top_core_EC_mc_n534) );
  XNOR2X1 U14175 ( .A(top_core_EC_mix_in[59]), .B(top_core_EC_mc_n537), .Y(
        top_core_EC_mc_n533) );
  XNOR2X1 U14176 ( .A(top_core_EC_mix_in[59]), .B(top_core_EC_mc_n416), .Y(
        top_core_EC_mc_n535) );
  OAI22X1 U14177 ( .A0(top_core_EC_mc_n525), .A1(n2481), .B0(n2379), .B1(
        top_core_EC_mc_n526), .Y(top_core_EC_mix_out_36_) );
  XOR2X1 U14178 ( .A(top_core_EC_mc_n527), .B(top_core_EC_mc_n528), .Y(
        top_core_EC_mc_n526) );
  XNOR2X1 U14179 ( .A(top_core_EC_mc_mix_in_8[63]), .B(top_core_EC_mc_n529), 
        .Y(top_core_EC_mc_n525) );
  XNOR2X1 U14180 ( .A(top_core_EC_mc_mix_in_8[63]), .B(top_core_EC_mc_n408), 
        .Y(top_core_EC_mc_n527) );
  OAI22X1 U14181 ( .A0(top_core_EC_mc_n517), .A1(n2481), .B0(n2379), .B1(
        top_core_EC_mc_n518), .Y(top_core_EC_mix_out_37_) );
  XOR2X1 U14182 ( .A(top_core_EC_mc_n519), .B(top_core_EC_mc_n520), .Y(
        top_core_EC_mc_n518) );
  XNOR2X1 U14183 ( .A(n1541), .B(top_core_EC_mc_n521), .Y(top_core_EC_mc_n517)
         );
  XNOR2X1 U14184 ( .A(n1541), .B(top_core_EC_mc_n400), .Y(top_core_EC_mc_n519)
         );
  OAI22X1 U14185 ( .A0(top_core_EC_mc_n509), .A1(n2482), .B0(n2380), .B1(
        top_core_EC_mc_n510), .Y(top_core_EC_mix_out_38_) );
  XOR2X1 U14186 ( .A(top_core_EC_mc_n511), .B(top_core_EC_mc_n512), .Y(
        top_core_EC_mc_n510) );
  XNOR2X1 U14187 ( .A(n1540), .B(top_core_EC_mc_n513), .Y(top_core_EC_mc_n509)
         );
  XNOR2X1 U14188 ( .A(n1540), .B(top_core_EC_mc_n392), .Y(top_core_EC_mc_n511)
         );
  OAI22X1 U14189 ( .A0(top_core_EC_mc_n501), .A1(n2482), .B0(n2380), .B1(
        top_core_EC_mc_n502), .Y(top_core_EC_mix_out_39_) );
  XOR2X1 U14190 ( .A(top_core_EC_mc_n503), .B(top_core_EC_mc_n504), .Y(
        top_core_EC_mc_n502) );
  XNOR2X1 U14191 ( .A(n1539), .B(top_core_EC_mc_n505), .Y(top_core_EC_mc_n501)
         );
  XNOR2X1 U14192 ( .A(n1539), .B(top_core_EC_mc_n384), .Y(top_core_EC_mc_n503)
         );
  OAI22X1 U14193 ( .A0(top_core_EC_mc_n444), .A1(n2470), .B0(n2380), .B1(
        top_core_EC_mc_n445), .Y(top_core_EC_mix_out_48_) );
  XOR2X1 U14194 ( .A(top_core_EC_mc_n373), .B(top_core_EC_mc_n446), .Y(
        top_core_EC_mc_n445) );
  XNOR2X1 U14195 ( .A(n1539), .B(top_core_EC_mc_n447), .Y(top_core_EC_mc_n444)
         );
  XOR2X1 U14196 ( .A(top_core_EC_mc_n447), .B(top_core_EC_mc_n448), .Y(
        top_core_EC_mc_n446) );
  OAI22X1 U14197 ( .A0(top_core_EC_mc_n395), .A1(n2464), .B0(n2381), .B1(
        top_core_EC_mc_n396), .Y(top_core_EC_mix_out_53_) );
  XOR2X1 U14198 ( .A(top_core_EC_mc_n324), .B(top_core_EC_mc_n397), .Y(
        top_core_EC_mc_n396) );
  XNOR2X1 U14199 ( .A(top_core_EC_mc_mix_in_8[63]), .B(top_core_EC_mc_n398), 
        .Y(top_core_EC_mc_n395) );
  XOR2X1 U14200 ( .A(top_core_EC_mc_n398), .B(top_core_EC_mc_n399), .Y(
        top_core_EC_mc_n397) );
  OAI22X1 U14201 ( .A0(top_core_EC_mc_n387), .A1(n2445), .B0(n2381), .B1(
        top_core_EC_mc_n388), .Y(top_core_EC_mix_out_54_) );
  XOR2X1 U14202 ( .A(top_core_EC_mc_n316), .B(top_core_EC_mc_n389), .Y(
        top_core_EC_mc_n388) );
  XNOR2X1 U14203 ( .A(n1541), .B(top_core_EC_mc_n390), .Y(top_core_EC_mc_n387)
         );
  XOR2X1 U14204 ( .A(top_core_EC_mc_n390), .B(top_core_EC_mc_n391), .Y(
        top_core_EC_mc_n389) );
  OAI22X1 U14205 ( .A0(top_core_EC_mc_n379), .A1(n2444), .B0(n2381), .B1(
        top_core_EC_mc_n380), .Y(top_core_EC_mix_out_55_) );
  XOR2X1 U14206 ( .A(top_core_EC_mc_n308), .B(top_core_EC_mc_n381), .Y(
        top_core_EC_mc_n380) );
  XNOR2X1 U14207 ( .A(n1540), .B(top_core_EC_mc_n382), .Y(top_core_EC_mc_n379)
         );
  XOR2X1 U14208 ( .A(top_core_EC_mc_n382), .B(top_core_EC_mc_n383), .Y(
        top_core_EC_mc_n381) );
  OAI22X1 U14209 ( .A0(top_core_EC_mc_n371), .A1(n2439), .B0(n2381), .B1(
        top_core_EC_mc_n372), .Y(top_core_EC_mix_out_56_) );
  XOR2X1 U14210 ( .A(top_core_EC_mc_n373), .B(top_core_EC_mc_n374), .Y(
        top_core_EC_mc_n372) );
  XNOR2X1 U14211 ( .A(n1539), .B(top_core_EC_mc_n375), .Y(top_core_EC_mc_n371)
         );
  XOR2X1 U14212 ( .A(top_core_EC_mc_n375), .B(top_core_EC_mc_n376), .Y(
        top_core_EC_mc_n374) );
  NAND2X1 U14213 ( .A(n577), .B(n761), .Y(n11673) );
  NAND2X1 U14214 ( .A(n578), .B(n762), .Y(top_core_KE_sb1_n98) );
  NAND2X1 U14215 ( .A(n579), .B(n760), .Y(n12304) );
  NAND2X1 U14216 ( .A(n580), .B(n756), .Y(n13250) );
  NAND2X1 U14217 ( .A(n581), .B(n763), .Y(n11989) );
  NAND2X1 U14218 ( .A(n582), .B(n758), .Y(n12935) );
  NAND2X1 U14219 ( .A(n583), .B(n759), .Y(n13565) );
  NAND2X1 U14220 ( .A(n584), .B(n757), .Y(n12620) );
  OAI221XL U14221 ( .A0(n3482), .A1(n91), .B0(n1143), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n104), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n105), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n94) );
  OAI221XL U14222 ( .A0(n2882), .A1(n90), .B0(n1001), .B1(n9919), .C0(n9920), 
        .Y(n9910) );
  OAI221XL U14223 ( .A0(n2640), .A1(n92), .B0(n945), .B1(n11087), .C0(n11088), 
        .Y(n11078) );
  OAI221XL U14224 ( .A0(n3242), .A1(n93), .B0(n1085), .B1(n8167), .C0(n8168), 
        .Y(n8158) );
  OAI221XL U14225 ( .A0(n2701), .A1(n94), .B0(n959), .B1(n10795), .C0(n10796), 
        .Y(n10786) );
  OAI221XL U14226 ( .A0(n3062), .A1(n96), .B0(n1043), .B1(n9043), .C0(n9044), 
        .Y(n9034) );
  OAI221XL U14227 ( .A0(n3422), .A1(n95), .B0(n1127), .B1(n7291), .C0(n7292), 
        .Y(n7282) );
  OAI221XL U14228 ( .A0(n2822), .A1(n97), .B0(n987), .B1(n10211), .C0(n10212), 
        .Y(n10202) );
  OAI221XL U14229 ( .A0(n3004), .A1(n98), .B0(n1029), .B1(n9335), .C0(n9336), 
        .Y(n9326) );
  OAI221XL U14230 ( .A0(n3181), .A1(n99), .B0(n1071), .B1(n8459), .C0(n8460), 
        .Y(n8450) );
  OAI221XL U14231 ( .A0(n3364), .A1(n100), .B0(n1113), .B1(n7583), .C0(n7584), 
        .Y(n7574) );
  OAI221XL U14232 ( .A0(n2579), .A1(n101), .B0(n931), .B1(n11379), .C0(n11380), 
        .Y(n11370) );
  OAI221XL U14233 ( .A0(n2761), .A1(n102), .B0(n973), .B1(n10503), .C0(n10504), 
        .Y(n10494) );
  OAI221XL U14234 ( .A0(n2943), .A1(n103), .B0(n1015), .B1(n9627), .C0(n9628), 
        .Y(n9618) );
  OAI221XL U14235 ( .A0(n3123), .A1(n104), .B0(n1057), .B1(n8751), .C0(n8752), 
        .Y(n8742) );
  OAI221XL U14236 ( .A0(n3303), .A1(n105), .B0(n1099), .B1(n7875), .C0(n7876), 
        .Y(n7866) );
  NAND2X1 U14237 ( .A(n751), .B(n1643), .Y(n13697) );
  NAND2X1 U14238 ( .A(n753), .B(n1211), .Y(n11806) );
  NAND2X1 U14239 ( .A(n754), .B(n1210), .Y(top_core_KE_sb1_n234) );
  NAND2X1 U14240 ( .A(n755), .B(n1170), .Y(n12122) );
  NAND2X1 U14241 ( .A(n745), .B(n1802), .Y(n11670) );
  NAND2X1 U14242 ( .A(n746), .B(n1823), .Y(top_core_KE_sb1_n95) );
  NAND2X1 U14243 ( .A(n744), .B(n1760), .Y(n12301) );
  NAND2X1 U14244 ( .A(n747), .B(n1781), .Y(n11986) );
  NAND2X1 U14245 ( .A(n748), .B(n1677), .Y(n13382) );
  NAND2X1 U14246 ( .A(n750), .B(n1707), .Y(n13067) );
  NAND2X1 U14247 ( .A(n749), .B(n1736), .Y(n12752) );
  INVX1 U14248 ( .A(n13979), .Y(n6126) );
  INVX1 U14249 ( .A(n17129), .Y(n5358) );
  INVX1 U14250 ( .A(n18389), .Y(n5004) );
  INVX1 U14251 ( .A(n15239), .Y(n5830) );
  INVX1 U14252 ( .A(n15554), .Y(n5746) );
  INVX1 U14253 ( .A(n18704), .Y(n4888) );
  INVX1 U14254 ( .A(n16814), .Y(n5442) );
  INVX1 U14255 ( .A(n14924), .Y(n5906) );
  INVX1 U14256 ( .A(n16499), .Y(n5518) );
  INVX1 U14257 ( .A(n18074), .Y(n5088) );
  INVX1 U14258 ( .A(n14609), .Y(n5982) );
  INVX1 U14259 ( .A(n16184), .Y(n5594) );
  INVX1 U14260 ( .A(n17759), .Y(n5196) );
  INVX1 U14261 ( .A(n14294), .Y(n6058) );
  INVX1 U14262 ( .A(n15869), .Y(n5670) );
  INVX1 U14263 ( .A(n17444), .Y(n5274) );
  AOI31X1 U14264 ( .A0(n12303), .A1(n12304), .A2(n12282), .B0(n12305), .Y(
        n12298) );
  OAI221XL U14265 ( .A0(n1667), .A1(n13516), .B0(n13268), .B1(n13428), .C0(
        n13517), .Y(n13508) );
  AOI21X1 U14266 ( .A0(n6472), .A1(n13518), .B0(n13519), .Y(n13517) );
  OAI32X1 U14267 ( .A0(n1675), .A1(n13520), .A2(n1672), .B0(n1172), .B1(n13252), .Y(n13519) );
  OAI221XL U14268 ( .A0(n1725), .A1(n12886), .B0(n12638), .B1(n12798), .C0(
        n12887), .Y(n12878) );
  AOI21X1 U14269 ( .A0(n6775), .A1(n12888), .B0(n12889), .Y(n12887) );
  OAI32X1 U14270 ( .A0(n1733), .A1(n12890), .A2(n1730), .B0(n1212), .B1(n12622), .Y(n12889) );
  OAI221XL U14271 ( .A0(n1696), .A1(n13201), .B0(n12953), .B1(n13113), .C0(
        n13202), .Y(n13193) );
  AOI21X1 U14272 ( .A0(n6815), .A1(n13203), .B0(n13204), .Y(n13202) );
  OAI32X1 U14273 ( .A0(n1704), .A1(n13205), .A2(n1701), .B0(n1218), .B1(n12937), .Y(n13204) );
  CLKINVX2 U14274 ( .A(n50), .Y(n6915) );
  CLKINVX2 U14275 ( .A(n51), .Y(n6869) );
  CLKINVX2 U14276 ( .A(n89), .Y(n6622) );
  CLKINVX2 U14277 ( .A(n52), .Y(n6550) );
  CLKINVX2 U14278 ( .A(n53), .Y(n6575) );
  CLKINVX2 U14279 ( .A(n54), .Y(n6845) );
  CLKINVX2 U14280 ( .A(n55), .Y(n6598) );
  CLKINVX2 U14281 ( .A(n56), .Y(n6891) );
  OAI211X1 U14282 ( .A0(n1173), .A1(n13495), .B0(n13496), .C0(n13497), .Y(
        n13494) );
  AOI31XL U14283 ( .A0(n1173), .A1(n13346), .A2(n13229), .B0(n6474), .Y(n13496) );
  NAND4X1 U14284 ( .A(n13460), .B(n13384), .C(n13499), .D(n13500), .Y(n13498)
         );
  OAI211X1 U14285 ( .A0(n1213), .A1(n12865), .B0(n12866), .C0(n12867), .Y(
        n12864) );
  AOI31XL U14286 ( .A0(n1213), .A1(n12716), .A2(n12599), .B0(n6777), .Y(n12866) );
  NAND4X1 U14287 ( .A(n12830), .B(n12754), .C(n12869), .D(n12870), .Y(n12868)
         );
  OAI211X1 U14288 ( .A0(n1219), .A1(n13180), .B0(n13181), .C0(n13182), .Y(
        n13179) );
  AOI31XL U14289 ( .A0(n1219), .A1(n13031), .A2(n12914), .B0(n6817), .Y(n13181) );
  NAND4X1 U14290 ( .A(n13145), .B(n13069), .C(n13184), .D(n13185), .Y(n13183)
         );
  NAND2X1 U14291 ( .A(n753), .B(n6830), .Y(n11675) );
  NAND2X1 U14292 ( .A(n754), .B(n6809), .Y(top_core_KE_sb1_n100) );
  NAND2X1 U14293 ( .A(n752), .B(n6534), .Y(n12306) );
  NAND2X1 U14294 ( .A(n755), .B(n6512), .Y(n11991) );
  NAND2X1 U14295 ( .A(n749), .B(n6780), .Y(n12622) );
  NAND2X1 U14296 ( .A(n751), .B(n6523), .Y(n13567) );
  NAND2X1 U14297 ( .A(n750), .B(n6819), .Y(n12937) );
  NAND2X1 U14298 ( .A(n748), .B(n6477), .Y(n13252) );
  AOI31X1 U14299 ( .A0(n1813), .A1(n1796), .A2(n745), .B0(n11656), .Y(n11913)
         );
  AOI31X1 U14300 ( .A0(n1834), .A1(n1817), .A2(n746), .B0(top_core_KE_sb1_n81), 
        .Y(top_core_KE_sb1_n342) );
  AOI31X1 U14301 ( .A0(n1771), .A1(n1752), .A2(n744), .B0(n12288), .Y(n12544)
         );
  AOI31X1 U14302 ( .A0(n1689), .A1(n1670), .A2(n1151), .B0(n13233), .Y(n13489)
         );
  AOI31X1 U14303 ( .A0(n1792), .A1(n1775), .A2(n747), .B0(n11972), .Y(n12229)
         );
  AOI31X1 U14304 ( .A0(n1747), .A1(n1728), .A2(n1191), .B0(n12603), .Y(n12859)
         );
  AOI31X1 U14305 ( .A0(n1661), .A1(n1635), .A2(n1160), .B0(n13548), .Y(n13804)
         );
  AOI31X1 U14306 ( .A0(n1718), .A1(n1699), .A2(n1200), .B0(n12918), .Y(n13174)
         );
  XOR2X1 U14307 ( .A(top_core_EC_mc_mix_in_2_112_), .B(top_core_EC_mix_in[112]), .Y(top_core_EC_mc_mix_in_4_114_) );
  XOR2X1 U14308 ( .A(top_core_EC_mc_mix_in_2_64_), .B(top_core_EC_mix_in[64]), 
        .Y(top_core_EC_mc_mix_in_4_66_) );
  XOR2X1 U14309 ( .A(top_core_EC_mc_mix_in_2_64_), .B(top_core_EC_mix_in[67]), 
        .Y(top_core_EC_mc_mix_in_8[70]) );
  XOR2X1 U14310 ( .A(top_core_EC_mc_mix_in_2_96_), .B(top_core_EC_mix_in[99]), 
        .Y(top_core_EC_mc_mix_in_8[102]) );
  XNOR2X1 U14311 ( .A(top_core_EC_mc_n562), .B(top_core_EC_mc_n563), .Y(
        top_core_EC_mc_n449) );
  XNOR2X1 U14312 ( .A(n1544), .B(top_core_EC_mc_mix_in_8[32]), .Y(
        top_core_EC_mc_n562) );
  XOR2X1 U14313 ( .A(n1541), .B(top_core_EC_mc_mix_in_8[48]), .Y(
        top_core_EC_mc_n563) );
  XNOR2X1 U14314 ( .A(top_core_EC_mc_n506), .B(top_core_EC_mc_n507), .Y(
        top_core_EC_mc_n384) );
  XNOR2X1 U14315 ( .A(top_core_EC_mc_mix_in_8[47]), .B(
        top_core_EC_mc_mix_in_8[39]), .Y(top_core_EC_mc_n506) );
  XOR2X1 U14316 ( .A(top_core_EC_mc_mix_in_8[63]), .B(
        top_core_EC_mc_mix_in_8[55]), .Y(top_core_EC_mc_n507) );
  XNOR2X1 U14317 ( .A(top_core_EC_mc_n303), .B(top_core_EC_mc_n304), .Y(
        top_core_EC_mc_n181) );
  XNOR2X1 U14318 ( .A(n1538), .B(top_core_EC_mc_mix_in_8[64]), .Y(
        top_core_EC_mc_n303) );
  XOR2X1 U14319 ( .A(n1535), .B(top_core_EC_mc_mix_in_8[80]), .Y(
        top_core_EC_mc_n304) );
  XNOR2X1 U14320 ( .A(top_core_EC_mc_n295), .B(top_core_EC_mc_n296), .Y(
        top_core_EC_mc_n173) );
  XNOR2X1 U14321 ( .A(top_core_EC_mc_mix_in_8[73]), .B(
        top_core_EC_mc_mix_in_8[65]), .Y(top_core_EC_mc_n295) );
  XOR2X1 U14322 ( .A(top_core_EC_mc_mix_in_8[89]), .B(
        top_core_EC_mc_mix_in_8[81]), .Y(top_core_EC_mc_n296) );
  XOR2X1 U14323 ( .A(n1538), .B(n1537), .Y(top_core_EC_mc_mix_in_8[73]) );
  XNOR2X1 U14324 ( .A(top_core_EC_mc_n279), .B(top_core_EC_mc_n280), .Y(
        top_core_EC_mc_n157) );
  XNOR2X1 U14325 ( .A(top_core_EC_mc_mix_in_8[75]), .B(
        top_core_EC_mc_mix_in_8[67]), .Y(top_core_EC_mc_n279) );
  XOR2X1 U14326 ( .A(top_core_EC_mc_mix_in_8[91]), .B(
        top_core_EC_mc_mix_in_8[83]), .Y(top_core_EC_mc_n280) );
  XOR2X1 U14327 ( .A(n1538), .B(top_core_EC_mc_mix_in_4_74_), .Y(
        top_core_EC_mc_mix_in_8[75]) );
  XNOR2X1 U14328 ( .A(top_core_EC_mc_n271), .B(top_core_EC_mc_n272), .Y(
        top_core_EC_mc_n149) );
  XNOR2X1 U14329 ( .A(top_core_EC_mc_mix_in_8[76]), .B(
        top_core_EC_mc_mix_in_8[68]), .Y(top_core_EC_mc_n271) );
  XOR2X1 U14330 ( .A(top_core_EC_mc_mix_in_8[92]), .B(
        top_core_EC_mc_mix_in_8[84]), .Y(top_core_EC_mc_n272) );
  XOR2X1 U14331 ( .A(n1538), .B(top_core_EC_mc_mix_in_4_75_), .Y(
        top_core_EC_mc_mix_in_8[76]) );
  XNOR2X1 U14332 ( .A(top_core_EC_mc_n238), .B(top_core_EC_mc_n239), .Y(
        top_core_EC_mc_n125) );
  XNOR2X1 U14333 ( .A(top_core_EC_mc_mix_in_8[79]), .B(
        top_core_EC_mc_mix_in_8[71]), .Y(top_core_EC_mc_n238) );
  XOR2X1 U14334 ( .A(top_core_EC_mc_mix_in_8[95]), .B(
        top_core_EC_mc_mix_in_8[87]), .Y(top_core_EC_mc_n239) );
  XNOR2X1 U14335 ( .A(top_core_EC_mc_n888), .B(top_core_EC_mc_n889), .Y(
        top_core_EC_mc_n44) );
  XNOR2X1 U14336 ( .A(top_core_EC_mc_mix_in_8[112]), .B(n1556), .Y(
        top_core_EC_mc_n888) );
  XOR2X1 U14337 ( .A(top_core_EC_mc_mix_in_8[96]), .B(n1553), .Y(
        top_core_EC_mc_n889) );
  XNOR2X1 U14338 ( .A(top_core_EC_mc_n881), .B(top_core_EC_mc_n882), .Y(
        top_core_EC_mc_n35) );
  XNOR2X1 U14339 ( .A(top_core_EC_mc_mix_in_8[113]), .B(
        top_core_EC_mc_mix_in_8[105]), .Y(top_core_EC_mc_n881) );
  XOR2X1 U14340 ( .A(top_core_EC_mc_mix_in_8[97]), .B(
        top_core_EC_mc_mix_in_8[121]), .Y(top_core_EC_mc_n882) );
  XOR2X1 U14341 ( .A(top_core_EC_mc_mix_in_8[112]), .B(
        top_core_EC_mc_mix_in_4_112_), .Y(top_core_EC_mc_mix_in_8[113]) );
  XNOR2X1 U14342 ( .A(top_core_EC_mc_n867), .B(top_core_EC_mc_n868), .Y(
        top_core_EC_mc_n17) );
  XNOR2X1 U14343 ( .A(top_core_EC_mc_mix_in_8[115]), .B(
        top_core_EC_mc_mix_in_8[107]), .Y(top_core_EC_mc_n867) );
  XOR2X1 U14344 ( .A(top_core_EC_mc_mix_in_8[99]), .B(
        top_core_EC_mc_mix_in_8[123]), .Y(top_core_EC_mc_n868) );
  XOR2X1 U14345 ( .A(top_core_EC_mc_mix_in_8[112]), .B(
        top_core_EC_mc_mix_in_4_114_), .Y(top_core_EC_mc_mix_in_8[115]) );
  XNOR2X1 U14346 ( .A(top_core_EC_mc_n919), .B(top_core_EC_mc_n920), .Y(
        top_core_EC_mc_n808) );
  XNOR2X1 U14347 ( .A(top_core_EC_mc_mix_in_8[108]), .B(
        top_core_EC_mc_mix_in_8[100]), .Y(top_core_EC_mc_n919) );
  XOR2X1 U14348 ( .A(top_core_EC_mc_mix_in_8[124]), .B(
        top_core_EC_mc_mix_in_8[116]), .Y(top_core_EC_mc_n920) );
  XOR2X1 U14349 ( .A(n1556), .B(top_core_EC_mc_mix_in_4_107_), .Y(
        top_core_EC_mc_mix_in_8[108]) );
  XNOR2X1 U14350 ( .A(top_core_EC_mc_n895), .B(top_core_EC_mc_n896), .Y(
        top_core_EC_mc_n784) );
  XNOR2X1 U14351 ( .A(top_core_EC_mc_mix_in_8[111]), .B(
        top_core_EC_mc_mix_in_8[103]), .Y(top_core_EC_mc_n895) );
  XOR2X1 U14352 ( .A(top_core_EC_mc_mix_in_8[127]), .B(
        top_core_EC_mc_mix_in_8[119]), .Y(top_core_EC_mc_n896) );
  AOI211X1 U14353 ( .A0(n6168), .A1(n1145), .B0(n6175), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n100), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n99) );
  AOI21X1 U14354 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n101), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n102), .B0(n530), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n100) );
  AOI211X1 U14355 ( .A0(n5383), .A1(n1004), .B0(n5388), .C0(n9916), .Y(n9915)
         );
  AOI21X1 U14356 ( .A0(n9917), .A1(n9918), .B0(n529), .Y(n9916) );
  AOI211X1 U14357 ( .A0(n5029), .A1(n948), .B0(n5034), .C0(n11084), .Y(n11083)
         );
  AOI21X1 U14358 ( .A0(n11085), .A1(n11086), .B0(n531), .Y(n11084) );
  AOI211X1 U14359 ( .A0(n5855), .A1(n1088), .B0(n5860), .C0(n8164), .Y(n8163)
         );
  AOI21X1 U14360 ( .A0(n8165), .A1(n8166), .B0(n532), .Y(n8164) );
  AOI211X1 U14361 ( .A0(n5113), .A1(n962), .B0(n5118), .C0(n10792), .Y(n10791)
         );
  AOI21X1 U14362 ( .A0(n10793), .A1(n10794), .B0(n533), .Y(n10792) );
  AOI211X1 U14363 ( .A0(n5619), .A1(n1046), .B0(n5624), .C0(n9040), .Y(n9039)
         );
  AOI21X1 U14364 ( .A0(n9041), .A1(n9042), .B0(n534), .Y(n9040) );
  AOI211X1 U14365 ( .A0(n6083), .A1(n1130), .B0(n6088), .C0(n7288), .Y(n7287)
         );
  AOI21X1 U14366 ( .A0(n7289), .A1(n7290), .B0(n535), .Y(n7288) );
  AOI211X1 U14367 ( .A0(n5299), .A1(n990), .B0(n5304), .C0(n10208), .Y(n10207)
         );
  AOI21X1 U14368 ( .A0(n10209), .A1(n10210), .B0(n536), .Y(n10208) );
  AOI211X1 U14369 ( .A0(n5543), .A1(n1032), .B0(n5548), .C0(n9332), .Y(n9331)
         );
  AOI21X1 U14370 ( .A0(n9333), .A1(n9334), .B0(n537), .Y(n9332) );
  AOI211X1 U14371 ( .A0(n5771), .A1(n1074), .B0(n5776), .C0(n8456), .Y(n8455)
         );
  AOI21X1 U14372 ( .A0(n8457), .A1(n8458), .B0(n538), .Y(n8456) );
  AOI211X1 U14373 ( .A0(n6007), .A1(n1116), .B0(n6012), .C0(n7580), .Y(n7579)
         );
  AOI21X1 U14374 ( .A0(n7581), .A1(n7582), .B0(n539), .Y(n7580) );
  AOI211X1 U14375 ( .A0(n4913), .A1(n934), .B0(n4918), .C0(n11376), .Y(n11375)
         );
  AOI21X1 U14376 ( .A0(n11377), .A1(n11378), .B0(n540), .Y(n11376) );
  AOI211X1 U14377 ( .A0(n5221), .A1(n976), .B0(n5226), .C0(n10500), .Y(n10499)
         );
  AOI21X1 U14378 ( .A0(n10501), .A1(n10502), .B0(n541), .Y(n10500) );
  AOI211X1 U14379 ( .A0(n5467), .A1(n1018), .B0(n5472), .C0(n9624), .Y(n9623)
         );
  AOI21X1 U14380 ( .A0(n9625), .A1(n9626), .B0(n542), .Y(n9624) );
  AOI211X1 U14381 ( .A0(n5695), .A1(n1060), .B0(n5700), .C0(n8748), .Y(n8747)
         );
  AOI21X1 U14382 ( .A0(n8749), .A1(n8750), .B0(n543), .Y(n8748) );
  AOI211X1 U14383 ( .A0(n5931), .A1(n1102), .B0(n5936), .C0(n7872), .Y(n7871)
         );
  AOI21X1 U14384 ( .A0(n7873), .A1(n7874), .B0(n544), .Y(n7872) );
  OAI22XL U14385 ( .A0(n1140), .A1(n3484), .B0(n3481), .B1(n13985), .Y(n14004)
         );
  OAI22XL U14386 ( .A0(n1000), .A1(n2883), .B0(n2880), .B1(n17135), .Y(n17154)
         );
  OAI22XL U14387 ( .A0(n944), .A1(n2643), .B0(n2638), .B1(n18395), .Y(n18414)
         );
  OAI22XL U14388 ( .A0(n1084), .A1(n3245), .B0(n3240), .B1(n15245), .Y(n15264)
         );
  OAI22XL U14389 ( .A0(n1070), .A1(n3190), .B0(n3179), .B1(n15560), .Y(n15579)
         );
  OAI22XL U14390 ( .A0(n930), .A1(n2588), .B0(n2577), .B1(n18710), .Y(n18729)
         );
  OAI22XL U14391 ( .A0(n1014), .A1(n2947), .B0(n2941), .B1(n16820), .Y(n16839)
         );
  OAI22XL U14392 ( .A0(n1098), .A1(n3306), .B0(n3301), .B1(n14930), .Y(n14949)
         );
  OAI22XL U14393 ( .A0(n1028), .A1(n3007), .B0(n3002), .B1(n16505), .Y(n16524)
         );
  OAI22XL U14394 ( .A0(n958), .A1(n2709), .B0(n2699), .B1(n18080), .Y(n18099)
         );
  OAI22XL U14395 ( .A0(n1112), .A1(n3373), .B0(n3362), .B1(n14615), .Y(n14634)
         );
  OAI22XL U14396 ( .A0(n1042), .A1(n3067), .B0(n3060), .B1(n16190), .Y(n16209)
         );
  OAI22XL U14397 ( .A0(n972), .A1(n2770), .B0(n2759), .B1(n17765), .Y(n17784)
         );
  OAI22XL U14398 ( .A0(n1126), .A1(n3425), .B0(n3420), .B1(n14300), .Y(n14319)
         );
  OAI22XL U14399 ( .A0(n1056), .A1(n3132), .B0(n3121), .B1(n15875), .Y(n15894)
         );
  OAI22XL U14400 ( .A0(n986), .A1(n2827), .B0(n2820), .B1(n17450), .Y(n17469)
         );
  XOR2X1 U14401 ( .A(top_core_EC_mc_mix_in_2_80_), .B(top_core_EC_mix_in[80]), 
        .Y(top_core_EC_mc_mix_in_4_82_) );
  XOR2X1 U14402 ( .A(top_core_EC_mc_mix_in_2_80_), .B(top_core_EC_mix_in[83]), 
        .Y(top_core_EC_mc_mix_in_8[86]) );
  XOR2X1 U14403 ( .A(top_core_EC_mc_mix_in_2_112_), .B(top_core_EC_mix_in[115]), .Y(top_core_EC_mc_mix_in_8[118]) );
  XOR2X1 U14404 ( .A(top_core_EC_mc_mix_in_2_96_), .B(top_core_EC_mix_in[96]), 
        .Y(top_core_EC_mc_mix_in_4_98_) );
  AOI21X1 U14405 ( .A0(n6539), .A1(n629), .B0(n13381), .Y(n13380) );
  AOI21X1 U14406 ( .A0(n6834), .A1(n630), .B0(n12751), .Y(n12750) );
  AOI21X1 U14407 ( .A0(n6880), .A1(n632), .B0(n13066), .Y(n13065) );
  AOI31X1 U14408 ( .A0(n5330), .A1(n1000), .A2(n450), .B0(n5329), .Y(n17292)
         );
  AOI31X1 U14409 ( .A0(n6114), .A1(n1140), .A2(n449), .B0(n6113), .Y(n14142)
         );
  AOI31X1 U14410 ( .A0(n5802), .A1(n1084), .A2(n452), .B0(n5801), .Y(n15402)
         );
  AOI31X1 U14411 ( .A0(n4976), .A1(n944), .A2(n451), .B0(n4975), .Y(n18552) );
  AOI31X1 U14412 ( .A0(n5718), .A1(n1070), .A2(n453), .B0(n5717), .Y(n15717)
         );
  AOI31X1 U14413 ( .A0(n5414), .A1(n1014), .A2(n455), .B0(n5413), .Y(n16977)
         );
  AOI31X1 U14414 ( .A0(n4860), .A1(n930), .A2(n454), .B0(n4859), .Y(n18867) );
  AOI31X1 U14415 ( .A0(n5878), .A1(n1098), .A2(n456), .B0(n5877), .Y(n15087)
         );
  AOI31X1 U14416 ( .A0(n5490), .A1(n1028), .A2(n457), .B0(n5489), .Y(n16662)
         );
  AOI31X1 U14417 ( .A0(n5060), .A1(n958), .A2(n458), .B0(n5059), .Y(n18237) );
  AOI31X1 U14418 ( .A0(n5954), .A1(n1112), .A2(n459), .B0(n5953), .Y(n14772)
         );
  AOI31X1 U14419 ( .A0(n5566), .A1(n1042), .A2(n460), .B0(n5565), .Y(n16347)
         );
  AOI31X1 U14420 ( .A0(n5168), .A1(n972), .A2(n461), .B0(n5167), .Y(n17922) );
  AOI31X1 U14421 ( .A0(n6030), .A1(n1126), .A2(n462), .B0(n6029), .Y(n14457)
         );
  AOI31X1 U14422 ( .A0(n5642), .A1(n1056), .A2(n463), .B0(n5641), .Y(n16032)
         );
  AOI31X1 U14423 ( .A0(n5246), .A1(n986), .A2(n464), .B0(n5245), .Y(n17607) );
  INVX1 U14424 ( .A(top_core_EC_n1024), .Y(n6305) );
  NOR4BX1 U14425 ( .AN(n12883), .B(n12884), .C(n6851), .D(n12628), .Y(n12881)
         );
  AOI21XL U14426 ( .A0(n12593), .A1(n6849), .B0(n12649), .Y(n12883) );
  OAI221XL U14427 ( .A0(n1212), .A1(n12798), .B0(n1750), .B1(n74), .C0(n12885), 
        .Y(n12884) );
  AOI22X1 U14428 ( .A0(n694), .A1(n1191), .B0(n6844), .B1(n1740), .Y(n12885)
         );
  NOR4BX1 U14429 ( .AN(n13828), .B(n13829), .C(n6604), .D(n13573), .Y(n13826)
         );
  AOI21XL U14430 ( .A0(n13538), .A1(n6602), .B0(n13594), .Y(n13828) );
  OAI221XL U14431 ( .A0(n1180), .A1(n13743), .B0(n1664), .B1(n76), .C0(n13830), 
        .Y(n13829) );
  AOI22X1 U14432 ( .A0(n695), .A1(n1160), .B0(n6597), .B1(n1653), .Y(n13830)
         );
  NOR4BX1 U14433 ( .AN(n13198), .B(n13199), .C(n6897), .D(n12943), .Y(n13196)
         );
  AOI21XL U14434 ( .A0(n12908), .A1(n6895), .B0(n12964), .Y(n13198) );
  OAI221XL U14435 ( .A0(n1218), .A1(n13113), .B0(n1721), .B1(n75), .C0(n13200), 
        .Y(n13199) );
  AOI22X1 U14436 ( .A0(n696), .A1(n1200), .B0(n6890), .B1(n1711), .Y(n13200)
         );
  NAND2X1 U14437 ( .A(n6914), .B(n1812), .Y(n11799) );
  NAND2X1 U14438 ( .A(n6868), .B(n1833), .Y(top_core_KE_sb1_n227) );
  NAND2X1 U14439 ( .A(n6621), .B(n1769), .Y(n12430) );
  NAND2X1 U14440 ( .A(n6549), .B(n1691), .Y(n13375) );
  NAND2X1 U14441 ( .A(n6574), .B(n1791), .Y(n12115) );
  NAND2X1 U14442 ( .A(n6844), .B(n1749), .Y(n12745) );
  NAND2X1 U14443 ( .A(n6597), .B(n1663), .Y(n13690) );
  NAND2X1 U14444 ( .A(n6890), .B(n1720), .Y(n13060) );
  NAND2X1 U14445 ( .A(n6914), .B(n1257), .Y(n11756) );
  NAND2X1 U14446 ( .A(n6868), .B(n1329), .Y(top_core_KE_sb1_n184) );
  NAND2X1 U14447 ( .A(n6621), .B(n1264), .Y(n12387) );
  NAND2X1 U14448 ( .A(n6574), .B(n1260), .Y(n12072) );
  NAND2X1 U14449 ( .A(n1202), .B(n1802), .Y(n11657) );
  NAND2X1 U14450 ( .A(n1193), .B(n1823), .Y(top_core_KE_sb1_n82) );
  NAND2X1 U14451 ( .A(n1153), .B(n1781), .Y(n11973) );
  NAND2X1 U14452 ( .A(n1162), .B(n1761), .Y(n12289) );
  NAND2X1 U14453 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n104), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n79), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n82) );
  NAND2X1 U14454 ( .A(n9919), .B(n9896), .Y(n9899) );
  NAND2X1 U14455 ( .A(n11087), .B(n11064), .Y(n11067) );
  NAND2X1 U14456 ( .A(n8167), .B(n8144), .Y(n8147) );
  NAND2X1 U14457 ( .A(n10795), .B(n10772), .Y(n10775) );
  NAND2X1 U14458 ( .A(n9043), .B(n9020), .Y(n9023) );
  NAND2X1 U14459 ( .A(n7291), .B(n7268), .Y(n7271) );
  NAND2X1 U14460 ( .A(n10211), .B(n10188), .Y(n10191) );
  NAND2X1 U14461 ( .A(n9335), .B(n9312), .Y(n9315) );
  NAND2X1 U14462 ( .A(n8459), .B(n8436), .Y(n8439) );
  NAND2X1 U14463 ( .A(n7583), .B(n7560), .Y(n7563) );
  NAND2X1 U14464 ( .A(n11379), .B(n11356), .Y(n11359) );
  NAND2X1 U14465 ( .A(n10503), .B(n10480), .Y(n10483) );
  NAND2X1 U14466 ( .A(n9627), .B(n9604), .Y(n9607) );
  NAND2X1 U14467 ( .A(n8751), .B(n8728), .Y(n8731) );
  NAND2X1 U14468 ( .A(n7875), .B(n7852), .Y(n7855) );
  AOI31XL U14469 ( .A0(n17099), .A1(n17072), .A2(n17042), .B0(n17035), .Y(
        n17118) );
  AOI31XL U14470 ( .A0(n13949), .A1(n13922), .A2(n13892), .B0(n13885), .Y(
        n13968) );
  AOI31XL U14471 ( .A0(n18359), .A1(n18332), .A2(n18302), .B0(n18295), .Y(
        n18378) );
  AOI31XL U14472 ( .A0(n15209), .A1(n15182), .A2(n15152), .B0(n15145), .Y(
        n15228) );
  AOI31XL U14473 ( .A0(n15524), .A1(n15497), .A2(n15467), .B0(n15460), .Y(
        n15543) );
  AOI31XL U14474 ( .A0(n18674), .A1(n18647), .A2(n18617), .B0(n18610), .Y(
        n18693) );
  AOI31XL U14475 ( .A0(n16784), .A1(n16757), .A2(n16727), .B0(n16720), .Y(
        n16803) );
  AOI31XL U14476 ( .A0(n14894), .A1(n14867), .A2(n14837), .B0(n14830), .Y(
        n14913) );
  AOI31XL U14477 ( .A0(n16469), .A1(n16442), .A2(n16412), .B0(n16405), .Y(
        n16488) );
  AOI31XL U14478 ( .A0(n18044), .A1(n18017), .A2(n17987), .B0(n17980), .Y(
        n18063) );
  AOI31XL U14479 ( .A0(n14579), .A1(n14552), .A2(n14522), .B0(n14515), .Y(
        n14598) );
  AOI31XL U14480 ( .A0(n16154), .A1(n16127), .A2(n16097), .B0(n16090), .Y(
        n16173) );
  AOI31XL U14481 ( .A0(n17729), .A1(n17702), .A2(n17672), .B0(n17665), .Y(
        n17748) );
  AOI31XL U14482 ( .A0(n14264), .A1(n14237), .A2(n14207), .B0(n14200), .Y(
        n14283) );
  AOI31XL U14483 ( .A0(n15839), .A1(n15812), .A2(n15782), .B0(n15775), .Y(
        n15858) );
  AOI31XL U14484 ( .A0(n17414), .A1(n17387), .A2(n17357), .B0(n17350), .Y(
        n17433) );
  NAND2X1 U14485 ( .A(n2875), .B(n1000), .Y(n10068) );
  NAND2X1 U14486 ( .A(n3479), .B(n1140), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n254) );
  NAND2X1 U14487 ( .A(n2633), .B(n944), .Y(n11236) );
  NAND2X1 U14488 ( .A(n3238), .B(n1084), .Y(n8316) );
  NAND2X1 U14489 ( .A(n2694), .B(n958), .Y(n10944) );
  NAND2X1 U14490 ( .A(n3055), .B(n1042), .Y(n9192) );
  NAND2X1 U14491 ( .A(n3415), .B(n1126), .Y(n7440) );
  NAND2X1 U14492 ( .A(n2818), .B(n986), .Y(n10360) );
  NAND2X1 U14493 ( .A(n2997), .B(n1028), .Y(n9484) );
  NAND2X1 U14494 ( .A(n3177), .B(n1070), .Y(n8608) );
  NAND2X1 U14495 ( .A(n3360), .B(n1112), .Y(n7732) );
  NAND2X1 U14496 ( .A(n2572), .B(n930), .Y(n11528) );
  NAND2X1 U14497 ( .A(n2757), .B(n972), .Y(n10652) );
  NAND2X1 U14498 ( .A(n2936), .B(n1014), .Y(n9776) );
  NAND2X1 U14499 ( .A(n3116), .B(n1056), .Y(n8900) );
  NAND2X1 U14500 ( .A(n3299), .B(n1098), .Y(n8024) );
  NOR2XL U14501 ( .A(n183), .B(n1658), .Y(n13770) );
  NOR2X1 U14502 ( .A(top_core_KE_n1870), .B(top_core_KE_n1871), .Y(
        top_core_KE_n2510) );
  AOI22XL U14503 ( .A0(n1802), .A1(n6914), .B0(n1259), .B1(n1202), .Y(n11864)
         );
  AOI22XL U14504 ( .A0(n1823), .A1(n6868), .B0(n1331), .B1(n1193), .Y(
        top_core_KE_sb1_n293) );
  AOI22XL U14505 ( .A0(n1760), .A1(n6621), .B0(n1266), .B1(n1162), .Y(n12495)
         );
  AOI22XL U14506 ( .A0(n1781), .A1(n6574), .B0(n1262), .B1(n1153), .Y(n12180)
         );
  AOI22XL U14507 ( .A0(n1259), .A1(n1202), .B0(n1221), .B1(n6917), .Y(n11720)
         );
  AOI22XL U14508 ( .A0(n1331), .A1(n1193), .B0(n1215), .B1(n6871), .Y(
        top_core_KE_sb1_n147) );
  AOI22XL U14509 ( .A0(n1266), .A1(n1162), .B0(n1183), .B1(n6624), .Y(n12351)
         );
  AOI22XL U14510 ( .A0(n1275), .A1(n1148), .B0(n1172), .B1(n6552), .Y(n13297)
         );
  AOI22XL U14511 ( .A0(n1262), .A1(n1153), .B0(n1175), .B1(n6577), .Y(n12036)
         );
  AOI22XL U14512 ( .A0(n1269), .A1(n1188), .B0(n1212), .B1(n6847), .Y(n12667)
         );
  AOI22XL U14513 ( .A0(n1272), .A1(n1197), .B0(n1218), .B1(n6893), .Y(n12982)
         );
  AOI22XL U14514 ( .A0(n1278), .A1(n1157), .B0(n1180), .B1(n6600), .Y(n13612)
         );
  AOI21X1 U14515 ( .A0(n1804), .A1(n761), .B0(n1205), .Y(n11727) );
  AOI21X1 U14516 ( .A0(n1825), .A1(n762), .B0(n1196), .Y(top_core_KE_sb1_n154)
         );
  AOI21X1 U14517 ( .A0(n1766), .A1(n760), .B0(n1165), .Y(n12358) );
  AOI21X1 U14518 ( .A0(n1682), .A1(n756), .B0(n1152), .Y(n13304) );
  AOI21X1 U14519 ( .A0(n1783), .A1(n763), .B0(n1156), .Y(n12043) );
  AOI21X1 U14520 ( .A0(n1740), .A1(n757), .B0(n1192), .Y(n12674) );
  AOI21X1 U14521 ( .A0(n1657), .A1(n759), .B0(n1161), .Y(n13619) );
  AOI21X1 U14522 ( .A0(n1711), .A1(n758), .B0(n1201), .Y(n12989) );
  NAND2X1 U14523 ( .A(n1809), .B(n753), .Y(n11650) );
  NAND2X1 U14524 ( .A(n1830), .B(n754), .Y(top_core_KE_sb1_n75) );
  NAND2X1 U14525 ( .A(n1767), .B(n752), .Y(n12282) );
  NAND2X1 U14526 ( .A(n1788), .B(n755), .Y(n11966) );
  NAND2X1 U14527 ( .A(n1716), .B(n750), .Y(n12912) );
  NAND2X1 U14528 ( .A(n1658), .B(n751), .Y(n13542) );
  NAND2X1 U14529 ( .A(n1745), .B(n749), .Y(n12597) );
  NAND2X1 U14530 ( .A(n1687), .B(n748), .Y(n13227) );
  NAND2X1 U14531 ( .A(n3473), .B(n1140), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n145) );
  NAND2X1 U14532 ( .A(n2872), .B(n1000), .Y(n9960) );
  NAND2X1 U14533 ( .A(n2630), .B(n944), .Y(n11128) );
  NAND2X1 U14534 ( .A(n3232), .B(n1084), .Y(n8208) );
  NAND2X1 U14535 ( .A(n2691), .B(n958), .Y(n10836) );
  NAND2X1 U14536 ( .A(n3052), .B(n1042), .Y(n9084) );
  NAND2X1 U14537 ( .A(n3412), .B(n1126), .Y(n7332) );
  NAND2X1 U14538 ( .A(n2812), .B(n986), .Y(n10252) );
  NAND2X1 U14539 ( .A(n2994), .B(n1028), .Y(n9376) );
  NAND2X1 U14540 ( .A(n3171), .B(n1070), .Y(n8500) );
  NAND2X1 U14541 ( .A(n3354), .B(n1112), .Y(n7624) );
  NAND2X1 U14542 ( .A(n2569), .B(n930), .Y(n11420) );
  NAND2X1 U14543 ( .A(n2751), .B(n972), .Y(n10544) );
  NAND2X1 U14544 ( .A(n2933), .B(n1014), .Y(n9668) );
  NAND2X1 U14545 ( .A(n3113), .B(n1056), .Y(n8792) );
  NAND2X1 U14546 ( .A(n3293), .B(n1098), .Y(n7916) );
  OAI211XL U14547 ( .A0(n3), .A1(n13238), .B0(n13349), .C0(n13356), .Y(n13353)
         );
  OAI211XL U14548 ( .A0(n11651), .A1(n50), .B0(n11686), .C0(n11648), .Y(n11749) );
  OAI211XL U14549 ( .A0(top_core_KE_sb1_n76), .A1(n51), .B0(
        top_core_KE_sb1_n111), .C0(top_core_KE_sb1_n73), .Y(
        top_core_KE_sb1_n177) );
  OAI211XL U14550 ( .A0(n12283), .A1(n89), .B0(n12317), .C0(n12280), .Y(n12380) );
  OAI211XL U14551 ( .A0(n13228), .A1(n52), .B0(n13263), .C0(n13225), .Y(n13326) );
  OAI211XL U14552 ( .A0(n11967), .A1(n53), .B0(n12002), .C0(n11964), .Y(n12065) );
  OAI211XL U14553 ( .A0(n12598), .A1(n54), .B0(n12633), .C0(n12595), .Y(n12696) );
  OAI211XL U14554 ( .A0(n13543), .A1(n55), .B0(n13578), .C0(n13540), .Y(n13641) );
  OAI211XL U14555 ( .A0(n12913), .A1(n56), .B0(n12948), .C0(n12910), .Y(n13011) );
  OAI211XL U14556 ( .A0(n1652), .A1(n6), .B0(n13626), .C0(n13755), .Y(n13771)
         );
  NAND2X1 U14557 ( .A(n681), .B(n6914), .Y(n11772) );
  NAND2X1 U14558 ( .A(n682), .B(n6868), .Y(top_core_KE_sb1_n200) );
  NAND2X1 U14559 ( .A(n683), .B(n6621), .Y(n12403) );
  NAND2X1 U14560 ( .A(n684), .B(n6574), .Y(n12088) );
  NAND2X1 U14561 ( .A(n1149), .B(n1687), .Y(n13350) );
  NAND2X1 U14562 ( .A(n1189), .B(n1745), .Y(n12720) );
  NAND2X1 U14563 ( .A(n1198), .B(n1716), .Y(n13035) );
  NAND2X1 U14564 ( .A(n1203), .B(n1809), .Y(n11773) );
  NAND2X1 U14565 ( .A(n1194), .B(n1830), .Y(top_core_KE_sb1_n201) );
  NAND2X1 U14566 ( .A(n1163), .B(n1767), .Y(n12404) );
  NAND2X1 U14567 ( .A(n1154), .B(n1788), .Y(n12089) );
  NAND2X1 U14568 ( .A(n1158), .B(n1658), .Y(n13665) );
  NAND2X1 U14569 ( .A(n1205), .B(n11651), .Y(n11669) );
  NAND2X1 U14570 ( .A(n1196), .B(top_core_KE_sb1_n76), .Y(top_core_KE_sb1_n94)
         );
  NAND2X1 U14571 ( .A(n1165), .B(n12283), .Y(n12300) );
  NAND2X1 U14572 ( .A(n1156), .B(n11967), .Y(n11985) );
  OAI21XL U14573 ( .A0(n996), .A1(n586), .B0(n1245), .Y(n10084) );
  OAI222XL U14574 ( .A0(n9891), .A1(n9918), .B0(n10003), .B1(n2887), .C0(n9970), .C1(n90), .Y(n10085) );
  OAI21XL U14575 ( .A0(n1139), .A1(n585), .B0(n1327), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n270) );
  OAI222XL U14576 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n74), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n102), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n189), .B1(n3485), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .C1(n91), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n271) );
  OAI21XL U14577 ( .A0(n940), .A1(n587), .B0(n1253), .Y(n11252) );
  OAI222XL U14578 ( .A0(n11059), .A1(n11086), .B0(n11171), .B1(n2645), .C0(
        n11138), .C1(n92), .Y(n11253) );
  OAI21XL U14579 ( .A0(n1080), .A1(n588), .B0(n1233), .Y(n8332) );
  OAI222XL U14580 ( .A0(n8139), .A1(n8166), .B0(n8251), .B1(n3247), .C0(n8218), 
        .C1(n93), .Y(n8333) );
  OAI21XL U14581 ( .A0(n954), .A1(n589), .B0(n1251), .Y(n10960) );
  OAI222XL U14582 ( .A0(n10767), .A1(n10794), .B0(n10879), .B1(n2707), .C0(
        n10846), .C1(n94), .Y(n10961) );
  OAI21XL U14583 ( .A0(n1122), .A1(n591), .B0(n1227), .Y(n7456) );
  OAI222XL U14584 ( .A0(n7263), .A1(n7290), .B0(n7375), .B1(n3427), .C0(n7342), 
        .C1(n95), .Y(n7457) );
  OAI21XL U14585 ( .A0(n1038), .A1(n590), .B0(n1239), .Y(n9208) );
  OAI222XL U14586 ( .A0(n9015), .A1(n9042), .B0(n9127), .B1(n3067), .C0(n9094), 
        .C1(n96), .Y(n9209) );
  OAI21XL U14587 ( .A0(n982), .A1(n592), .B0(n1247), .Y(n10376) );
  OAI222XL U14588 ( .A0(n10183), .A1(n10210), .B0(n10295), .B1(n2827), .C0(
        n10262), .C1(n97), .Y(n10377) );
  OAI21XL U14589 ( .A0(n1024), .A1(n593), .B0(n1241), .Y(n9500) );
  OAI222XL U14590 ( .A0(n9307), .A1(n9334), .B0(n9419), .B1(n3009), .C0(n9386), 
        .C1(n98), .Y(n9501) );
  OAI21XL U14591 ( .A0(n1066), .A1(n594), .B0(n1235), .Y(n8624) );
  OAI222XL U14592 ( .A0(n8431), .A1(n8458), .B0(n8543), .B1(n3187), .C0(n8510), 
        .C1(n99), .Y(n8625) );
  OAI21XL U14593 ( .A0(n1108), .A1(n595), .B0(n1229), .Y(n7748) );
  OAI222XL U14594 ( .A0(n7555), .A1(n7582), .B0(n7667), .B1(n3370), .C0(n7634), 
        .C1(n100), .Y(n7749) );
  OAI21XL U14595 ( .A0(n926), .A1(n596), .B0(n1255), .Y(n11544) );
  OAI222XL U14596 ( .A0(n11351), .A1(n11378), .B0(n11463), .B1(n2585), .C0(
        n11430), .C1(n101), .Y(n11545) );
  OAI21XL U14597 ( .A0(n968), .A1(n597), .B0(n1249), .Y(n10668) );
  OAI222XL U14598 ( .A0(n10475), .A1(n10502), .B0(n10587), .B1(n2767), .C0(
        n10554), .C1(n102), .Y(n10669) );
  OAI21XL U14599 ( .A0(n1010), .A1(n598), .B0(n1243), .Y(n9792) );
  OAI222XL U14600 ( .A0(n9599), .A1(n9626), .B0(n9711), .B1(n2948), .C0(n9678), 
        .C1(n103), .Y(n9793) );
  OAI21XL U14601 ( .A0(n1052), .A1(n599), .B0(n1237), .Y(n8916) );
  OAI222XL U14602 ( .A0(n8723), .A1(n8750), .B0(n8835), .B1(n3129), .C0(n8802), 
        .C1(n104), .Y(n8917) );
  OAI21XL U14603 ( .A0(n1094), .A1(n600), .B0(n1231), .Y(n8040) );
  OAI222XL U14604 ( .A0(n7847), .A1(n7874), .B0(n7959), .B1(n3308), .C0(n7926), 
        .C1(n105), .Y(n8041) );
  NAND2X1 U14605 ( .A(n1203), .B(n1805), .Y(n11672) );
  NAND2X1 U14606 ( .A(n1194), .B(n1826), .Y(top_core_KE_sb1_n97) );
  NAND2X1 U14607 ( .A(n1163), .B(n1763), .Y(n12303) );
  NAND2X1 U14608 ( .A(n1154), .B(n1784), .Y(n11988) );
  NAND2X1 U14609 ( .A(n1189), .B(n1740), .Y(n12619) );
  NAND2X1 U14610 ( .A(n1158), .B(n1655), .Y(n13564) );
  NAND2X1 U14611 ( .A(n1198), .B(n1711), .Y(n12934) );
  NAND2X1 U14612 ( .A(n1149), .B(n1682), .Y(n13249) );
  AOI22XL U14613 ( .A0(n13238), .A1(n1673), .B0(n1678), .B1(n13268), .Y(n13239) );
  AOI22XL U14614 ( .A0(n12923), .A1(n1702), .B0(n1706), .B1(n12953), .Y(n12924) );
  AOI22XL U14615 ( .A0(n12608), .A1(n1731), .B0(n1735), .B1(n12638), .Y(n12609) );
  NAND2X1 U14616 ( .A(n6826), .B(n761), .Y(n11919) );
  NAND2X1 U14617 ( .A(n6804), .B(n762), .Y(top_core_KE_sb1_n348) );
  NAND2X1 U14618 ( .A(n6530), .B(n760), .Y(n12550) );
  NAND2X1 U14619 ( .A(n6472), .B(n756), .Y(n13495) );
  NAND2X1 U14620 ( .A(n6507), .B(n763), .Y(n12235) );
  NAND2X1 U14621 ( .A(n6815), .B(n758), .Y(n13180) );
  NAND2X1 U14622 ( .A(n6519), .B(n759), .Y(n13810) );
  NAND2X1 U14623 ( .A(n6775), .B(n757), .Y(n12865) );
  NAND2X1 U14624 ( .A(n1202), .B(n1221), .Y(n11648) );
  NAND2X1 U14625 ( .A(n1193), .B(n1215), .Y(top_core_KE_sb1_n73) );
  NAND2X1 U14626 ( .A(n1162), .B(n1183), .Y(n12280) );
  NAND2X1 U14627 ( .A(n1153), .B(n1175), .Y(n11964) );
  NAND2X1 U14628 ( .A(n1221), .B(n6914), .Y(n11671) );
  NAND2X1 U14629 ( .A(n1215), .B(n6868), .Y(top_core_KE_sb1_n96) );
  NAND2X1 U14630 ( .A(n1183), .B(n6621), .Y(n12302) );
  NAND2X1 U14631 ( .A(n1175), .B(n6574), .Y(n11987) );
  NOR2X1 U14632 ( .A(n13601), .B(n695), .Y(n13627) );
  NAND3XL U14633 ( .A(n11646), .B(n1211), .C(n11769), .Y(n11884) );
  NAND3XL U14634 ( .A(top_core_KE_sb1_n71), .B(n1210), .C(top_core_KE_sb1_n197), .Y(top_core_KE_sb1_n313) );
  NAND3XL U14635 ( .A(n13223), .B(n1677), .C(n13346), .Y(n13460) );
  NAND3XL U14636 ( .A(n11962), .B(n1170), .C(n12085), .Y(n12200) );
  NAND3XL U14637 ( .A(n12593), .B(n1736), .C(n12716), .Y(n12830) );
  NAND3XL U14638 ( .A(n13538), .B(n1644), .C(n13661), .Y(n13775) );
  NAND3XL U14639 ( .A(n12908), .B(n1707), .C(n13031), .Y(n13145) );
  AOI31X1 U14640 ( .A0(n17081), .A1(n17082), .A2(n5356), .B0(n16997), .Y(
        n17080) );
  INVX1 U14641 ( .A(n17083), .Y(n5356) );
  OAI21XL U14642 ( .A0(n17072), .A1(n17074), .B0(n17084), .Y(n17083) );
  AOI31X1 U14643 ( .A0(n13931), .A1(n13932), .A2(n6124), .B0(n13847), .Y(
        n13930) );
  INVX1 U14644 ( .A(n13933), .Y(n6124) );
  OAI21XL U14645 ( .A0(n13922), .A1(n13924), .B0(n13934), .Y(n13933) );
  AOI31X1 U14646 ( .A0(n18341), .A1(n18342), .A2(n5002), .B0(n18257), .Y(
        n18340) );
  INVX1 U14647 ( .A(n18343), .Y(n5002) );
  OAI21XL U14648 ( .A0(n18332), .A1(n18334), .B0(n18344), .Y(n18343) );
  AOI31X1 U14649 ( .A0(n15191), .A1(n15192), .A2(n5828), .B0(n15107), .Y(
        n15190) );
  INVX1 U14650 ( .A(n15193), .Y(n5828) );
  OAI21XL U14651 ( .A0(n15182), .A1(n15184), .B0(n15194), .Y(n15193) );
  AOI31X1 U14652 ( .A0(n15506), .A1(n15507), .A2(n5744), .B0(n15422), .Y(
        n15505) );
  INVX1 U14653 ( .A(n15508), .Y(n5744) );
  OAI21XL U14654 ( .A0(n15497), .A1(n15499), .B0(n15509), .Y(n15508) );
  AOI31X1 U14655 ( .A0(n18656), .A1(n18657), .A2(n4886), .B0(n18572), .Y(
        n18655) );
  INVX1 U14656 ( .A(n18658), .Y(n4886) );
  OAI21XL U14657 ( .A0(n18647), .A1(n18649), .B0(n18659), .Y(n18658) );
  AOI31X1 U14658 ( .A0(n16766), .A1(n16767), .A2(n5440), .B0(n16682), .Y(
        n16765) );
  INVX1 U14659 ( .A(n16768), .Y(n5440) );
  OAI21XL U14660 ( .A0(n16757), .A1(n16759), .B0(n16769), .Y(n16768) );
  AOI31X1 U14661 ( .A0(n14876), .A1(n14877), .A2(n5904), .B0(n14792), .Y(
        n14875) );
  INVX1 U14662 ( .A(n14878), .Y(n5904) );
  OAI21XL U14663 ( .A0(n14867), .A1(n14869), .B0(n14879), .Y(n14878) );
  AOI31X1 U14664 ( .A0(n16451), .A1(n16452), .A2(n5516), .B0(n16367), .Y(
        n16450) );
  INVX1 U14665 ( .A(n16453), .Y(n5516) );
  OAI21XL U14666 ( .A0(n16442), .A1(n16444), .B0(n16454), .Y(n16453) );
  AOI31X1 U14667 ( .A0(n18026), .A1(n18027), .A2(n5086), .B0(n17942), .Y(
        n18025) );
  INVX1 U14668 ( .A(n18028), .Y(n5086) );
  OAI21XL U14669 ( .A0(n18017), .A1(n18019), .B0(n18029), .Y(n18028) );
  AOI31X1 U14670 ( .A0(n14561), .A1(n14562), .A2(n5980), .B0(n14477), .Y(
        n14560) );
  INVX1 U14671 ( .A(n14563), .Y(n5980) );
  OAI21XL U14672 ( .A0(n14552), .A1(n14554), .B0(n14564), .Y(n14563) );
  AOI31X1 U14673 ( .A0(n16136), .A1(n16137), .A2(n5592), .B0(n16052), .Y(
        n16135) );
  INVX1 U14674 ( .A(n16138), .Y(n5592) );
  OAI21XL U14675 ( .A0(n16127), .A1(n16129), .B0(n16139), .Y(n16138) );
  AOI31X1 U14676 ( .A0(n17711), .A1(n17712), .A2(n5194), .B0(n17627), .Y(
        n17710) );
  INVX1 U14677 ( .A(n17713), .Y(n5194) );
  OAI21XL U14678 ( .A0(n17702), .A1(n17704), .B0(n17714), .Y(n17713) );
  AOI31X1 U14679 ( .A0(n14246), .A1(n14247), .A2(n6056), .B0(n14162), .Y(
        n14245) );
  INVX1 U14680 ( .A(n14248), .Y(n6056) );
  OAI21XL U14681 ( .A0(n14237), .A1(n14239), .B0(n14249), .Y(n14248) );
  AOI31X1 U14682 ( .A0(n15821), .A1(n15822), .A2(n5668), .B0(n15737), .Y(
        n15820) );
  INVX1 U14683 ( .A(n15823), .Y(n5668) );
  OAI21XL U14684 ( .A0(n15812), .A1(n15814), .B0(n15824), .Y(n15823) );
  AOI31X1 U14685 ( .A0(n17396), .A1(n17397), .A2(n5272), .B0(n17312), .Y(
        n17395) );
  INVX1 U14686 ( .A(n17398), .Y(n5272) );
  OAI21XL U14687 ( .A0(n17387), .A1(n17389), .B0(n17399), .Y(n17398) );
  AOI31X1 U14688 ( .A0(n14103), .A1(n13934), .A2(n14104), .B0(n3462), .Y(
        n14101) );
  AOI222X1 U14689 ( .A0(n6172), .A1(n3476), .B0(n13869), .B1(n514), .C0(n6166), 
        .C1(n3491), .Y(n14104) );
  AOI31X1 U14690 ( .A0(n17253), .A1(n17084), .A2(n17254), .B0(n2862), .Y(
        n17251) );
  AOI222X1 U14691 ( .A0(n5390), .A1(n2878), .B0(n17019), .B1(n513), .C0(n5376), 
        .C1(n2888), .Y(n17254) );
  AOI31X1 U14692 ( .A0(n18513), .A1(n18344), .A2(n18514), .B0(n2619), .Y(
        n18511) );
  AOI222X1 U14693 ( .A0(n5036), .A1(n2636), .B0(n18279), .B1(n515), .C0(n5022), 
        .C1(n2646), .Y(n18514) );
  AOI31X1 U14694 ( .A0(n15363), .A1(n15194), .A2(n15364), .B0(n3222), .Y(
        n15361) );
  AOI222X1 U14695 ( .A0(n5862), .A1(n3238), .B0(n15129), .B1(n516), .C0(n5848), 
        .C1(n3248), .Y(n15364) );
  AOI31X1 U14696 ( .A0(n15678), .A1(n15509), .A2(n15679), .B0(n3160), .Y(
        n15676) );
  AOI222X1 U14697 ( .A0(n5778), .A1(n3177), .B0(n15444), .B1(n517), .C0(n5764), 
        .C1(n3188), .Y(n15679) );
  AOI31X1 U14698 ( .A0(n18828), .A1(n18659), .A2(n18829), .B0(n2557), .Y(
        n18826) );
  AOI222X1 U14699 ( .A0(n4920), .A1(n2575), .B0(n18594), .B1(n518), .C0(n4906), 
        .C1(n2586), .Y(n18829) );
  AOI31X1 U14700 ( .A0(n16938), .A1(n16769), .A2(n16939), .B0(n2922), .Y(
        n16936) );
  AOI222X1 U14701 ( .A0(n5474), .A1(n2939), .B0(n16704), .B1(n519), .C0(n5460), 
        .C1(n2949), .Y(n16939) );
  AOI31X1 U14702 ( .A0(n15048), .A1(n14879), .A2(n15049), .B0(n3282), .Y(
        n15046) );
  AOI222X1 U14703 ( .A0(n5938), .A1(n3299), .B0(n14814), .B1(n520), .C0(n5924), 
        .C1(n3309), .Y(n15049) );
  AOI31X1 U14704 ( .A0(n16623), .A1(n16454), .A2(n16624), .B0(n2983), .Y(
        n16621) );
  AOI222X1 U14705 ( .A0(n5550), .A1(n3000), .B0(n16389), .B1(n521), .C0(n5536), 
        .C1(n3010), .Y(n16624) );
  AOI31X1 U14706 ( .A0(n18198), .A1(n18029), .A2(n18199), .B0(n2681), .Y(
        n18196) );
  AOI222X1 U14707 ( .A0(n5120), .A1(n2697), .B0(n17964), .B1(n522), .C0(n5106), 
        .C1(n2708), .Y(n18199) );
  AOI31X1 U14708 ( .A0(n14733), .A1(n14564), .A2(n14734), .B0(n3343), .Y(
        n14731) );
  AOI222X1 U14709 ( .A0(n6014), .A1(n3360), .B0(n14499), .B1(n523), .C0(n6000), 
        .C1(n3371), .Y(n14734) );
  AOI31X1 U14710 ( .A0(n16308), .A1(n16139), .A2(n16309), .B0(n3041), .Y(
        n16306) );
  AOI222X1 U14711 ( .A0(n5626), .A1(n3058), .B0(n16074), .B1(n524), .C0(n5612), 
        .C1(n3068), .Y(n16309) );
  AOI31X1 U14712 ( .A0(n17883), .A1(n17714), .A2(n17884), .B0(n2741), .Y(
        n17881) );
  AOI222X1 U14713 ( .A0(n5228), .A1(n2757), .B0(n17649), .B1(n525), .C0(n5214), 
        .C1(n2768), .Y(n17884) );
  AOI31X1 U14714 ( .A0(n14418), .A1(n14249), .A2(n14419), .B0(n3401), .Y(
        n14416) );
  AOI222X1 U14715 ( .A0(n6090), .A1(n3418), .B0(n14184), .B1(n526), .C0(n6076), 
        .C1(n3428), .Y(n14419) );
  AOI31X1 U14716 ( .A0(n15993), .A1(n15824), .A2(n15994), .B0(n3103), .Y(
        n15991) );
  AOI222X1 U14717 ( .A0(n5702), .A1(n3119), .B0(n15759), .B1(n527), .C0(n5688), 
        .C1(n3130), .Y(n15994) );
  AOI31X1 U14718 ( .A0(n17568), .A1(n17399), .A2(n17569), .B0(n2801), .Y(
        n17566) );
  AOI222X1 U14719 ( .A0(n5306), .A1(n2818), .B0(n17334), .B1(n528), .C0(n5292), 
        .C1(n2828), .Y(n17569) );
  AOI31X1 U14720 ( .A0(n11648), .A1(n6922), .A2(n11649), .B0(n1796), .Y(n11647) );
  AOI21X1 U14721 ( .A0(n6914), .A1(n1802), .B0(n6918), .Y(n11649) );
  INVX1 U14722 ( .A(n11650), .Y(n6918) );
  AOI31X1 U14723 ( .A0(top_core_KE_sb1_n73), .A1(n6876), .A2(
        top_core_KE_sb1_n74), .B0(n1817), .Y(top_core_KE_sb1_n72) );
  AOI21X1 U14724 ( .A0(n6868), .A1(n1823), .B0(n6872), .Y(top_core_KE_sb1_n74)
         );
  INVX1 U14725 ( .A(top_core_KE_sb1_n75), .Y(n6872) );
  AOI31X1 U14726 ( .A0(n11964), .A1(n6582), .A2(n11965), .B0(n1775), .Y(n11963) );
  AOI21X1 U14727 ( .A0(n6574), .A1(n1781), .B0(n6578), .Y(n11965) );
  INVX1 U14728 ( .A(n11966), .Y(n6578) );
  AOI31X1 U14729 ( .A0(n12280), .A1(n6629), .A2(n12281), .B0(n1753), .Y(n12279) );
  AOI21X1 U14730 ( .A0(n6621), .A1(n1760), .B0(n6625), .Y(n12281) );
  INVX1 U14731 ( .A(n12282), .Y(n6625) );
  AOI31X1 U14732 ( .A0(n13225), .A1(n6558), .A2(n13226), .B0(n1672), .Y(n13224) );
  AOI21X1 U14733 ( .A0(n6549), .A1(n1680), .B0(n6553), .Y(n13226) );
  INVX1 U14734 ( .A(n13227), .Y(n6553) );
  AOI31X1 U14735 ( .A0(n12910), .A1(n6899), .A2(n12911), .B0(n1701), .Y(n12909) );
  AOI21X1 U14736 ( .A0(n6890), .A1(n1709), .B0(n6894), .Y(n12911) );
  INVX1 U14737 ( .A(n12912), .Y(n6894) );
  AOI31X1 U14738 ( .A0(n13540), .A1(n6606), .A2(n13541), .B0(n1636), .Y(n13539) );
  AOI21X1 U14739 ( .A0(n6597), .A1(n1651), .B0(n6601), .Y(n13541) );
  INVX1 U14740 ( .A(n13542), .Y(n6601) );
  AOI31X1 U14741 ( .A0(n12595), .A1(n6853), .A2(n12596), .B0(n1730), .Y(n12594) );
  AOI21X1 U14742 ( .A0(n6844), .A1(n1738), .B0(n6848), .Y(n12596) );
  INVX1 U14743 ( .A(n12597), .Y(n6848) );
  AOI31X1 U14744 ( .A0(n13418), .A1(n13419), .A2(n13420), .B0(n13277), .Y(
        n13417) );
  AOI222X1 U14745 ( .A0(n13313), .A1(n748), .B0(n1148), .B1(n1693), .C0(n677), 
        .C1(n1152), .Y(n13420) );
  AOI22X1 U14746 ( .A0(n6544), .A1(n1687), .B0(n6539), .B1(n1174), .Y(n13418)
         );
  AOI31X1 U14747 ( .A0(n12788), .A1(n12789), .A2(n12790), .B0(n12647), .Y(
        n12787) );
  AOI222X1 U14748 ( .A0(n12683), .A1(n749), .B0(n1188), .B1(n1751), .C0(n678), 
        .C1(n1192), .Y(n12790) );
  AOI22X1 U14749 ( .A0(n6839), .A1(n1745), .B0(n6834), .B1(n1214), .Y(n12788)
         );
  AOI31X1 U14750 ( .A0(n13103), .A1(n13104), .A2(n13105), .B0(n12962), .Y(
        n13102) );
  AOI222X1 U14751 ( .A0(n12998), .A1(n750), .B0(n1197), .B1(n1722), .C0(n680), 
        .C1(n1201), .Y(n13105) );
  AOI22X1 U14752 ( .A0(n6885), .A1(n1716), .B0(n6880), .B1(n1220), .Y(n13103)
         );
  AOI21XL U14753 ( .A0(n1258), .A1(n6914), .B0(n11879), .Y(n11689) );
  AOI21XL U14754 ( .A0(n1330), .A1(n6868), .B0(top_core_KE_sb1_n308), .Y(
        top_core_KE_sb1_n114) );
  AOI21XL U14755 ( .A0(n1265), .A1(n6621), .B0(n12510), .Y(n12320) );
  AOI21XL U14756 ( .A0(n1261), .A1(n6574), .B0(n12195), .Y(n12005) );
  NOR2X1 U14757 ( .A(n2291), .B(top_core_KE_n2695), .Y(top_core_KE_n2692) );
  NAND2X1 U14758 ( .A(n2846), .B(n992), .Y(n9932) );
  NAND2X1 U14759 ( .A(n3447), .B(n1132), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n117) );
  NAND2X1 U14760 ( .A(n2604), .B(n936), .Y(n11100) );
  NAND2X1 U14761 ( .A(n3206), .B(n1076), .Y(n8180) );
  NAND2X1 U14762 ( .A(n2665), .B(n950), .Y(n10808) );
  NAND2X1 U14763 ( .A(n3026), .B(n1034), .Y(n9056) );
  NAND2X1 U14764 ( .A(n3386), .B(n1118), .Y(n7304) );
  NAND2X1 U14765 ( .A(n2786), .B(n978), .Y(n10224) );
  NAND2X1 U14766 ( .A(n2968), .B(n1020), .Y(n9348) );
  NAND2X1 U14767 ( .A(n3145), .B(n1062), .Y(n8472) );
  NAND2X1 U14768 ( .A(n3328), .B(n1104), .Y(n7596) );
  NAND2X1 U14769 ( .A(n2543), .B(n922), .Y(n11392) );
  NAND2X1 U14770 ( .A(n2725), .B(n964), .Y(n10516) );
  NAND2X1 U14771 ( .A(n2907), .B(n1006), .Y(n9640) );
  NAND2X1 U14772 ( .A(n3087), .B(n1048), .Y(n8764) );
  NAND2X1 U14773 ( .A(n3267), .B(n1090), .Y(n7888) );
  NAND2X1 U14774 ( .A(n2849), .B(n992), .Y(n9934) );
  NAND2X1 U14775 ( .A(n3450), .B(n1132), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n119) );
  NAND2X1 U14776 ( .A(n2607), .B(n936), .Y(n11102) );
  NAND2X1 U14777 ( .A(n3209), .B(n1076), .Y(n8182) );
  NAND2X1 U14778 ( .A(n2668), .B(n950), .Y(n10810) );
  NAND2X1 U14779 ( .A(n3029), .B(n1034), .Y(n9058) );
  NAND2X1 U14780 ( .A(n3389), .B(n1118), .Y(n7306) );
  NAND2X1 U14781 ( .A(n2789), .B(n978), .Y(n10226) );
  NAND2X1 U14782 ( .A(n2971), .B(n1020), .Y(n9350) );
  NAND2X1 U14783 ( .A(n3148), .B(n1062), .Y(n8474) );
  NAND2X1 U14784 ( .A(n3331), .B(n1104), .Y(n7598) );
  NAND2X1 U14785 ( .A(n2546), .B(n922), .Y(n11394) );
  NAND2X1 U14786 ( .A(n2728), .B(n964), .Y(n10518) );
  NAND2X1 U14787 ( .A(n2910), .B(n1006), .Y(n9642) );
  NAND2X1 U14788 ( .A(n3090), .B(n1048), .Y(n8766) );
  NAND2X1 U14789 ( .A(n3270), .B(n1090), .Y(n7890) );
  NAND2X1 U14790 ( .A(n665), .B(n753), .Y(n11686) );
  NAND2X1 U14791 ( .A(n666), .B(n754), .Y(top_core_KE_sb1_n111) );
  NAND2X1 U14792 ( .A(n667), .B(n752), .Y(n12317) );
  NAND2X1 U14793 ( .A(n670), .B(n748), .Y(n13263) );
  NAND2X1 U14794 ( .A(n668), .B(n755), .Y(n12002) );
  NAND2X1 U14795 ( .A(n671), .B(n749), .Y(n12633) );
  NAND2X1 U14796 ( .A(n669), .B(n751), .Y(n13578) );
  NAND2X1 U14797 ( .A(n672), .B(n750), .Y(n12948) );
  INVX1 U14798 ( .A(n11679), .Y(n6830) );
  INVX1 U14799 ( .A(top_core_KE_sb1_n104), .Y(n6809) );
  INVX1 U14800 ( .A(n12310), .Y(n6534) );
  INVX1 U14801 ( .A(n11995), .Y(n6512) );
  INVX1 U14802 ( .A(n13571), .Y(n6523) );
  NOR2X1 U14803 ( .A(n618), .B(n625), .Y(n11929) );
  XNOR2X1 U14804 ( .A(n6964), .B(n1809), .Y(n618) );
  NOR2X1 U14805 ( .A(n619), .B(n626), .Y(top_core_KE_sb1_n358) );
  XNOR2X1 U14806 ( .A(n6958), .B(n1830), .Y(n619) );
  NOR2X1 U14807 ( .A(n620), .B(n629), .Y(n13505) );
  XNOR2X1 U14808 ( .A(n1676), .B(n1687), .Y(n620) );
  NOR2X1 U14809 ( .A(n621), .B(n628), .Y(n12245) );
  XNOR2X1 U14810 ( .A(n6670), .B(n1788), .Y(n621) );
  NOR2X1 U14811 ( .A(n622), .B(n630), .Y(n12875) );
  XNOR2X1 U14812 ( .A(n1734), .B(n1745), .Y(n622) );
  NOR2X1 U14813 ( .A(n623), .B(n631), .Y(n13820) );
  XNOR2X1 U14814 ( .A(n1643), .B(n1658), .Y(n623) );
  NOR2X1 U14815 ( .A(n624), .B(n632), .Y(n13190) );
  XNOR2X1 U14816 ( .A(n1705), .B(n1716), .Y(n624) );
  NAND2X1 U14817 ( .A(n17153), .B(n2893), .Y(n17224) );
  NAND2X1 U14818 ( .A(n14003), .B(n3494), .Y(n14074) );
  NAND2X1 U14819 ( .A(n15263), .B(n3253), .Y(n15334) );
  NAND2X1 U14820 ( .A(n18413), .B(n2650), .Y(n18484) );
  NAND2X1 U14821 ( .A(n15578), .B(n3192), .Y(n15649) );
  NAND2X1 U14822 ( .A(n16838), .B(n2954), .Y(n16909) );
  NAND2X1 U14823 ( .A(n18728), .B(n2600), .Y(n18799) );
  NAND2X1 U14824 ( .A(n14948), .B(n3314), .Y(n15019) );
  NAND2X1 U14825 ( .A(n16523), .B(n3015), .Y(n16594) );
  NAND2X1 U14826 ( .A(n18098), .B(n2711), .Y(n18169) );
  NAND2X1 U14827 ( .A(n14633), .B(n3375), .Y(n14704) );
  NAND2X1 U14828 ( .A(n16208), .B(n3072), .Y(n16279) );
  NAND2X1 U14829 ( .A(n17783), .B(n2772), .Y(n17854) );
  NAND2X1 U14830 ( .A(n14318), .B(n3433), .Y(n14389) );
  NAND2X1 U14831 ( .A(n15893), .B(n3134), .Y(n15964) );
  NAND2X1 U14832 ( .A(n17468), .B(n2833), .Y(n17539) );
  INVX1 U14833 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n218), .Y(n6174) );
  INVX1 U14834 ( .A(n8280), .Y(n5859) );
  INVX1 U14835 ( .A(n10032), .Y(n5387) );
  INVX1 U14836 ( .A(n11200), .Y(n5033) );
  INVX1 U14837 ( .A(n10908), .Y(n5117) );
  INVX1 U14838 ( .A(n9156), .Y(n5623) );
  INVX1 U14839 ( .A(n7404), .Y(n6087) );
  INVX1 U14840 ( .A(n10324), .Y(n5303) );
  INVX1 U14841 ( .A(n9448), .Y(n5547) );
  INVX1 U14842 ( .A(n8572), .Y(n5775) );
  INVX1 U14843 ( .A(n7696), .Y(n6011) );
  INVX1 U14844 ( .A(n11492), .Y(n4917) );
  INVX1 U14845 ( .A(n10616), .Y(n5225) );
  INVX1 U14846 ( .A(n9740), .Y(n5471) );
  INVX1 U14847 ( .A(n8864), .Y(n5699) );
  INVX1 U14848 ( .A(n7988), .Y(n5935) );
  XOR2X1 U14849 ( .A(top_core_EC_mc_mix_in_4_112_), .B(
        top_core_EC_mc_mix_in_2_114_), .Y(top_core_EC_mc_mix_in_4_115_) );
  XOR2X1 U14850 ( .A(top_core_EC_mc_mix_in_4_64_), .B(
        top_core_EC_mc_mix_in_2_66_), .Y(top_core_EC_mc_mix_in_4_67_) );
  XOR2X1 U14851 ( .A(top_core_EC_mc_mix_in_8[64]), .B(
        top_core_EC_mc_mix_in_8[80]), .Y(top_core_EC_mc_n70) );
  XOR2X1 U14852 ( .A(top_core_EC_mc_mix_in_4_64_), .B(
        top_core_EC_mc_mix_in_4_80_), .Y(top_core_EC_mc_n62) );
  XOR2X1 U14853 ( .A(top_core_EC_mc_mix_in_4_64_), .B(
        top_core_EC_mc_mix_in_2_64_), .Y(top_core_EC_mc_mix_in_8[66]) );
  XOR2X1 U14854 ( .A(top_core_EC_mc_mix_in_4_64_), .B(
        top_core_EC_mc_mix_in_2_67_), .Y(top_core_EC_mc_mix_in_8[69]) );
  XOR2X1 U14855 ( .A(top_core_EC_mc_mix_in_8[96]), .B(
        top_core_EC_mc_mix_in_8[112]), .Y(top_core_EC_mc_n735) );
  XOR2X1 U14856 ( .A(top_core_EC_mc_mix_in_4_96_), .B(
        top_core_EC_mc_mix_in_4_112_), .Y(top_core_EC_mc_n727) );
  XOR2X1 U14857 ( .A(top_core_EC_mc_mix_in_4_96_), .B(
        top_core_EC_mc_mix_in_2_99_), .Y(top_core_EC_mc_mix_in_8[101]) );
  CLKINVX3 U14858 ( .A(n12337), .Y(n6627) );
  XOR2X1 U14859 ( .A(top_core_EC_mc_mix_in_2_80_), .B(top_core_EC_mix_in[82]), 
        .Y(top_core_EC_mc_mix_in_2_83_) );
  XOR2X1 U14860 ( .A(top_core_EC_mc_mix_in_2_112_), .B(top_core_EC_mix_in[114]), .Y(top_core_EC_mc_mix_in_2_115_) );
  XOR2X1 U14861 ( .A(top_core_EC_mc_mix_in_2_64_), .B(top_core_EC_mix_in[66]), 
        .Y(top_core_EC_mc_mix_in_2_67_) );
  XOR2X1 U14862 ( .A(top_core_EC_mc_mix_in_2_96_), .B(top_core_EC_mix_in[98]), 
        .Y(top_core_EC_mc_mix_in_2_99_) );
  XOR2X1 U14863 ( .A(top_core_EC_mc_mix_in_2_64_), .B(
        top_core_EC_mc_mix_in_2_80_), .Y(top_core_EC_mc_n54) );
  XOR2X1 U14864 ( .A(top_core_EC_mc_mix_in_2_96_), .B(
        top_core_EC_mc_mix_in_2_112_), .Y(top_core_EC_mc_n719) );
  XOR2X1 U14865 ( .A(top_core_EC_mc_mix_in_2_106_), .B(
        top_core_EC_mc_mix_in_4_98_), .Y(top_core_EC_mc_n37) );
  XOR2X1 U14866 ( .A(top_core_EC_mc_mix_in_8[71]), .B(
        top_core_EC_mc_mix_in_8[87]), .Y(top_core_EC_mc_n78) );
  XOR2X1 U14867 ( .A(top_core_EC_mc_mix_in_8[103]), .B(
        top_core_EC_mc_mix_in_8[119]), .Y(top_core_EC_mc_n743) );
  XOR2X1 U14868 ( .A(top_core_EC_mix_in[104]), .B(top_core_EC_mc_mix_in_2_96_), 
        .Y(top_core_EC_mc_n46) );
  XOR2X1 U14869 ( .A(top_core_EC_mc_mix_in_2_66_), .B(
        top_core_EC_mc_mix_in_2_82_), .Y(top_core_EC_mc_n111) );
  XOR2X1 U14870 ( .A(n1537), .B(top_core_EC_mc_mix_in_2_74_), .Y(
        top_core_EC_mc_mix_in_4_75_) );
  XOR2X1 U14871 ( .A(n1555), .B(top_core_EC_mc_mix_in_2_106_), .Y(
        top_core_EC_mc_mix_in_4_107_) );
  XOR2X1 U14872 ( .A(top_core_EC_mix_in[64]), .B(top_core_EC_mix_in[80]), .Y(
        top_core_EC_mc_n119) );
  XOR2X1 U14873 ( .A(top_core_EC_mix_in[66]), .B(top_core_EC_mix_in[82]), .Y(
        top_core_EC_mc_n94) );
  XOR2X1 U14874 ( .A(top_core_EC_mix_in[67]), .B(top_core_EC_mix_in[83]), .Y(
        top_core_EC_mc_n86) );
  XOR2X1 U14875 ( .A(top_core_EC_mix_in[106]), .B(top_core_EC_mc_mix_in_2_98_), 
        .Y(top_core_EC_mc_n28) );
  XOR2X1 U14876 ( .A(top_core_EC_mix_in[107]), .B(top_core_EC_mc_mix_in_2_99_), 
        .Y(top_core_EC_mc_n19) );
  CLKINVX3 U14877 ( .A(n13608), .Y(n6597) );
  XNOR2X1 U14878 ( .A(top_core_EC_mc_n305), .B(top_core_EC_mc_n118), .Y(
        top_core_EC_mc_n302) );
  XNOR2X1 U14879 ( .A(top_core_EC_mix_in[80]), .B(n1536), .Y(
        top_core_EC_mc_n305) );
  XNOR2X1 U14880 ( .A(top_core_EC_mc_n297), .B(top_core_EC_mc_n110), .Y(
        top_core_EC_mc_n294) );
  XNOR2X1 U14881 ( .A(top_core_EC_mc_mix_in_2_82_), .B(
        top_core_EC_mc_mix_in_4_74_), .Y(top_core_EC_mc_n297) );
  XNOR2X1 U14882 ( .A(top_core_EC_mc_n289), .B(top_core_EC_mc_n93), .Y(
        top_core_EC_mc_n286) );
  XNOR2X1 U14883 ( .A(top_core_EC_mix_in[82]), .B(top_core_EC_mc_mix_in_2_74_), 
        .Y(top_core_EC_mc_n289) );
  XNOR2X1 U14884 ( .A(top_core_EC_mc_n281), .B(top_core_EC_mc_n85), .Y(
        top_core_EC_mc_n278) );
  XNOR2X1 U14885 ( .A(top_core_EC_mix_in[83]), .B(top_core_EC_mc_mix_in_2_75_), 
        .Y(top_core_EC_mc_n281) );
  XNOR2X1 U14886 ( .A(top_core_EC_mc_n273), .B(top_core_EC_mc_n77), .Y(
        top_core_EC_mc_n270) );
  XNOR2X1 U14887 ( .A(top_core_EC_mc_mix_in_8[87]), .B(
        top_core_EC_mc_mix_in_8[78]), .Y(top_core_EC_mc_n273) );
  XNOR2X1 U14888 ( .A(top_core_EC_mc_n265), .B(top_core_EC_mc_n69), .Y(
        top_core_EC_mc_n262) );
  XNOR2X1 U14889 ( .A(top_core_EC_mc_mix_in_8[80]), .B(
        top_core_EC_mc_mix_in_8[79]), .Y(top_core_EC_mc_n265) );
  XNOR2X1 U14890 ( .A(top_core_EC_mc_n248), .B(top_core_EC_mc_n61), .Y(
        top_core_EC_mc_n245) );
  XNOR2X1 U14891 ( .A(top_core_EC_mc_mix_in_4_80_), .B(n1538), .Y(
        top_core_EC_mc_n248) );
  XNOR2X1 U14892 ( .A(top_core_EC_mc_n240), .B(top_core_EC_mc_n53), .Y(
        top_core_EC_mc_n237) );
  XNOR2X1 U14893 ( .A(top_core_EC_mc_mix_in_2_80_), .B(n1537), .Y(
        top_core_EC_mc_n240) );
  XNOR2X1 U14894 ( .A(top_core_EC_mc_n921), .B(top_core_EC_mc_n742), .Y(
        top_core_EC_mc_n918) );
  XNOR2X1 U14895 ( .A(top_core_EC_mc_mix_in_8[119]), .B(
        top_core_EC_mc_mix_in_8[110]), .Y(top_core_EC_mc_n921) );
  XNOR2X1 U14896 ( .A(top_core_EC_mc_n913), .B(top_core_EC_mc_n734), .Y(
        top_core_EC_mc_n910) );
  XNOR2X1 U14897 ( .A(top_core_EC_mc_mix_in_8[112]), .B(
        top_core_EC_mc_mix_in_8[111]), .Y(top_core_EC_mc_n913) );
  XNOR2X1 U14898 ( .A(top_core_EC_mc_n905), .B(top_core_EC_mc_n726), .Y(
        top_core_EC_mc_n902) );
  XNOR2X1 U14899 ( .A(top_core_EC_mc_mix_in_4_112_), .B(n1556), .Y(
        top_core_EC_mc_n905) );
  XNOR2X1 U14900 ( .A(top_core_EC_mc_n897), .B(top_core_EC_mc_n718), .Y(
        top_core_EC_mc_n894) );
  XNOR2X1 U14901 ( .A(top_core_EC_mc_mix_in_2_112_), .B(n1555), .Y(
        top_core_EC_mc_n897) );
  XNOR2X1 U14902 ( .A(top_core_EC_mc_n833), .B(top_core_EC_mc_n834), .Y(
        top_core_EC_mc_n832) );
  XNOR2X1 U14903 ( .A(top_core_EC_mix_in[104]), .B(top_core_EC_mix_in[96]), 
        .Y(top_core_EC_mc_n833) );
  XNOR2X1 U14904 ( .A(top_core_EC_mc_n827), .B(top_core_EC_mc_n828), .Y(
        top_core_EC_mc_n826) );
  XNOR2X1 U14905 ( .A(top_core_EC_mc_mix_in_2_106_), .B(
        top_core_EC_mc_mix_in_2_98_), .Y(top_core_EC_mc_n827) );
  XNOR2X1 U14906 ( .A(top_core_EC_mc_n821), .B(top_core_EC_mc_n822), .Y(
        top_core_EC_mc_n820) );
  XNOR2X1 U14907 ( .A(top_core_EC_mix_in[106]), .B(top_core_EC_mix_in[98]), 
        .Y(top_core_EC_mc_n821) );
  XNOR2X1 U14908 ( .A(top_core_EC_mc_n815), .B(top_core_EC_mc_n816), .Y(
        top_core_EC_mc_n814) );
  XNOR2X1 U14909 ( .A(top_core_EC_mix_in[107]), .B(top_core_EC_mix_in[99]), 
        .Y(top_core_EC_mc_n815) );
  XOR2X1 U14910 ( .A(n1555), .B(n1554), .Y(top_core_EC_mc_mix_in_8[106]) );
  OAI22XL U14911 ( .A0(n1174), .A1(n180), .B0(n1689), .B1(n3), .Y(n13490) );
  NAND2X1 U14912 ( .A(n17019), .B(n1002), .Y(n17110) );
  NAND2X1 U14913 ( .A(n13869), .B(n1141), .Y(n13960) );
  NAND2X1 U14914 ( .A(n18279), .B(n946), .Y(n18370) );
  NAND2X1 U14915 ( .A(n15129), .B(n1086), .Y(n15220) );
  NAND2X1 U14916 ( .A(n15444), .B(n1072), .Y(n15535) );
  NAND2X1 U14917 ( .A(n18594), .B(n932), .Y(n18685) );
  NAND2X1 U14918 ( .A(n16704), .B(n1016), .Y(n16795) );
  NAND2X1 U14919 ( .A(n14814), .B(n1100), .Y(n14905) );
  NAND2X1 U14920 ( .A(n16389), .B(n1030), .Y(n16480) );
  NAND2X1 U14921 ( .A(n17964), .B(n960), .Y(n18055) );
  NAND2X1 U14922 ( .A(n14499), .B(n1114), .Y(n14590) );
  NAND2X1 U14923 ( .A(n16074), .B(n1044), .Y(n16165) );
  NAND2X1 U14924 ( .A(n17649), .B(n974), .Y(n17740) );
  NAND2X1 U14925 ( .A(n14184), .B(n1128), .Y(n14275) );
  NAND2X1 U14926 ( .A(n15759), .B(n1058), .Y(n15850) );
  NAND2X1 U14927 ( .A(n17334), .B(n988), .Y(n17425) );
  XOR2X1 U14928 ( .A(top_core_EC_mc_mix_in_4_112_), .B(
        top_core_EC_mc_mix_in_2_115_), .Y(top_core_EC_mc_mix_in_8[117]) );
  XOR2X1 U14929 ( .A(top_core_EC_mc_mix_in_4_80_), .B(
        top_core_EC_mc_mix_in_2_82_), .Y(top_core_EC_mc_mix_in_4_83_) );
  XOR2X1 U14930 ( .A(top_core_EC_mc_mix_in_4_80_), .B(
        top_core_EC_mc_mix_in_2_80_), .Y(top_core_EC_mc_mix_in_8[82]) );
  XOR2X1 U14931 ( .A(top_core_EC_mc_mix_in_4_80_), .B(
        top_core_EC_mc_mix_in_2_83_), .Y(top_core_EC_mc_mix_in_8[85]) );
  XOR2X1 U14932 ( .A(top_core_EC_mc_mix_in_4_80_), .B(
        top_core_EC_mc_mix_in_4_64_), .Y(top_core_EC_mc_n180) );
  XOR2X1 U14933 ( .A(top_core_EC_mc_mix_in_8[80]), .B(
        top_core_EC_mc_mix_in_8[64]), .Y(top_core_EC_mc_n124) );
  XOR2X1 U14934 ( .A(top_core_EC_mc_mix_in_4_96_), .B(
        top_core_EC_mc_mix_in_2_98_), .Y(top_core_EC_mc_mix_in_4_99_) );
  XOR2X1 U14935 ( .A(top_core_EC_mc_mix_in_4_96_), .B(
        top_core_EC_mc_mix_in_4_112_), .Y(top_core_EC_mc_n43) );
  XOR2X1 U14936 ( .A(top_core_EC_mc_mix_in_8[112]), .B(
        top_core_EC_mc_mix_in_8[96]), .Y(top_core_EC_mc_n783) );
  XOR2X1 U14937 ( .A(top_core_EC_mc_mix_in_8[63]), .B(
        top_core_EC_mc_mix_in_8[47]), .Y(top_core_EC_mc_n319) );
  XOR2X1 U14938 ( .A(top_core_EC_mc_mix_in_8[95]), .B(
        top_core_EC_mc_mix_in_8[79]), .Y(top_core_EC_mc_n60) );
  XOR2X1 U14939 ( .A(top_core_EC_mc_mix_in_8[127]), .B(
        top_core_EC_mc_mix_in_8[111]), .Y(top_core_EC_mc_n725) );
  XOR2X1 U14940 ( .A(top_core_EC_mc_mix_in_8[63]), .B(
        top_core_EC_mc_mix_in_8[54]), .Y(top_core_EC_mc_n410) );
  XOR2X1 U14941 ( .A(top_core_EC_mc_mix_in_8[95]), .B(
        top_core_EC_mc_mix_in_8[86]), .Y(top_core_EC_mc_n151) );
  XOR2X1 U14942 ( .A(top_core_EC_mc_mix_in_8[127]), .B(
        top_core_EC_mc_mix_in_8[118]), .Y(top_core_EC_mc_n810) );
  XOR2X1 U14943 ( .A(top_core_EC_mc_mix_in_4_112_), .B(
        top_core_EC_mc_mix_in_2_112_), .Y(top_core_EC_mc_mix_in_8[114]) );
  XOR2X1 U14944 ( .A(top_core_EC_mc_mix_in_8[79]), .B(
        top_core_EC_mc_mix_in_8[70]), .Y(top_core_EC_mc_n77) );
  XOR2X1 U14945 ( .A(top_core_EC_mc_mix_in_8[111]), .B(
        top_core_EC_mc_mix_in_8[102]), .Y(top_core_EC_mc_n742) );
  XOR2X1 U14946 ( .A(top_core_EC_mc_mix_in_2_90_), .B(
        top_core_EC_mc_mix_in_4_82_), .Y(top_core_EC_mc_n175) );
  XOR2X1 U14947 ( .A(top_core_EC_mc_mix_in_2_122_), .B(
        top_core_EC_mc_mix_in_4_114_), .Y(top_core_EC_mc_n828) );
  XOR2X1 U14948 ( .A(top_core_EC_mc_mix_in_2_74_), .B(
        top_core_EC_mc_mix_in_4_66_), .Y(top_core_EC_mc_n110) );
  XOR2X1 U14949 ( .A(n1551), .B(top_core_EC_mc_mix_in_4_112_), .Y(
        top_core_EC_mc_n786) );
  XOR2X1 U14950 ( .A(n1540), .B(top_core_EC_mc_mix_in_8[48]), .Y(
        top_core_EC_mc_n394) );
  XOR2X1 U14951 ( .A(n1539), .B(top_core_EC_mc_mix_in_4_48_), .Y(
        top_core_EC_mc_n386) );
  XOR2X1 U14952 ( .A(n1534), .B(top_core_EC_mc_mix_in_8[80]), .Y(
        top_core_EC_mc_n135) );
  XOR2X1 U14953 ( .A(n1533), .B(top_core_EC_mc_mix_in_4_80_), .Y(
        top_core_EC_mc_n127) );
  XOR2X1 U14954 ( .A(n1537), .B(top_core_EC_mc_mix_in_8[64]), .Y(
        top_core_EC_mc_n61) );
  XOR2X1 U14955 ( .A(n1536), .B(top_core_EC_mc_mix_in_4_64_), .Y(
        top_core_EC_mc_n53) );
  XOR2X1 U14956 ( .A(n1555), .B(top_core_EC_mc_mix_in_8[96]), .Y(
        top_core_EC_mc_n726) );
  XOR2X1 U14957 ( .A(n1554), .B(top_core_EC_mc_mix_in_4_96_), .Y(
        top_core_EC_mc_n718) );
  XOR2X1 U14958 ( .A(n1552), .B(top_core_EC_mc_mix_in_8[112]), .Y(
        top_core_EC_mc_n794) );
  XOR2X1 U14959 ( .A(top_core_EC_mc_mix_in_8[87]), .B(
        top_core_EC_mc_mix_in_8[71]), .Y(top_core_EC_mc_n132) );
  XOR2X1 U14960 ( .A(top_core_EC_mc_mix_in_8[119]), .B(
        top_core_EC_mc_mix_in_8[103]), .Y(top_core_EC_mc_n791) );
  XOR2X1 U14961 ( .A(top_core_EC_mix_in[88]), .B(top_core_EC_mc_mix_in_2_80_), 
        .Y(top_core_EC_mc_n183) );
  XOR2X1 U14962 ( .A(top_core_EC_mix_in[120]), .B(top_core_EC_mc_mix_in_2_112_), .Y(top_core_EC_mc_n834) );
  XOR2X1 U14963 ( .A(top_core_EC_mix_in[72]), .B(top_core_EC_mc_mix_in_2_64_), 
        .Y(top_core_EC_mc_n118) );
  XOR2X1 U14964 ( .A(n1540), .B(top_core_EC_mc_mix_in_2_58_), .Y(
        top_core_EC_mc_mix_in_4_59_) );
  XOR2X1 U14965 ( .A(n1534), .B(top_core_EC_mc_mix_in_2_90_), .Y(
        top_core_EC_mc_mix_in_4_91_) );
  XOR2X1 U14966 ( .A(n1552), .B(top_core_EC_mc_mix_in_2_122_), .Y(
        top_core_EC_mc_mix_in_4_123_) );
  XOR2X1 U14967 ( .A(top_core_EC_mc_mix_in_2_114_), .B(
        top_core_EC_mc_mix_in_2_98_), .Y(top_core_EC_mc_n764) );
  XOR2X1 U14968 ( .A(top_core_EC_mix_in[58]), .B(top_core_EC_mc_mix_in_2_50_), 
        .Y(top_core_EC_mc_n426) );
  XOR2X1 U14969 ( .A(top_core_EC_mix_in[59]), .B(top_core_EC_mc_mix_in_2_51_), 
        .Y(top_core_EC_mc_n418) );
  XOR2X1 U14970 ( .A(top_core_EC_mix_in[90]), .B(top_core_EC_mc_mix_in_2_82_), 
        .Y(top_core_EC_mc_n167) );
  XOR2X1 U14971 ( .A(top_core_EC_mix_in[91]), .B(top_core_EC_mc_mix_in_2_83_), 
        .Y(top_core_EC_mc_n159) );
  XOR2X1 U14972 ( .A(top_core_EC_mix_in[122]), .B(top_core_EC_mc_mix_in_2_114_), .Y(top_core_EC_mc_n822) );
  XOR2X1 U14973 ( .A(top_core_EC_mix_in[123]), .B(top_core_EC_mc_mix_in_2_115_), .Y(top_core_EC_mc_n816) );
  XOR2X1 U14974 ( .A(top_core_EC_mix_in[74]), .B(top_core_EC_mc_mix_in_2_66_), 
        .Y(top_core_EC_mc_n93) );
  XOR2X1 U14975 ( .A(top_core_EC_mix_in[75]), .B(top_core_EC_mc_mix_in_2_67_), 
        .Y(top_core_EC_mc_n85) );
  XOR2X1 U14976 ( .A(top_core_EC_mix_in[112]), .B(top_core_EC_mix_in[96]), .Y(
        top_core_EC_mc_n771) );
  XOR2X1 U14977 ( .A(top_core_EC_mix_in[114]), .B(top_core_EC_mix_in[98]), .Y(
        top_core_EC_mc_n757) );
  XOR2X1 U14978 ( .A(top_core_EC_mix_in[115]), .B(top_core_EC_mix_in[99]), .Y(
        top_core_EC_mc_n750) );
  XOR2X1 U14979 ( .A(n1541), .B(top_core_EC_mc_mix_in_8[55]), .Y(
        top_core_EC_mc_n402) );
  XOR2X1 U14980 ( .A(n1535), .B(top_core_EC_mc_mix_in_8[87]), .Y(
        top_core_EC_mc_n143) );
  XOR2X1 U14981 ( .A(n1538), .B(top_core_EC_mc_mix_in_8[71]), .Y(
        top_core_EC_mc_n69) );
  XOR2X1 U14982 ( .A(n1553), .B(top_core_EC_mc_mix_in_8[119]), .Y(
        top_core_EC_mc_n802) );
  XOR2X1 U14983 ( .A(n1556), .B(top_core_EC_mc_mix_in_8[103]), .Y(
        top_core_EC_mc_n734) );
  NAND2XL U14984 ( .A(n13415), .B(n13282), .Y(n13305) );
  NAND2XL U14985 ( .A(n11839), .B(n11705), .Y(n11728) );
  NAND2XL U14986 ( .A(top_core_KE_sb1_n268), .B(top_core_KE_sb1_n130), .Y(
        top_core_KE_sb1_n155) );
  NAND2XL U14987 ( .A(n12470), .B(n12336), .Y(n12359) );
  NAND2XL U14988 ( .A(n12155), .B(n12021), .Y(n12044) );
  NAND2XL U14989 ( .A(n12785), .B(n1269), .Y(n12675) );
  NAND2XL U14990 ( .A(n13100), .B(n1272), .Y(n12990) );
  NAND2XL U14991 ( .A(n13730), .B(n1278), .Y(n13620) );
  XNOR2X1 U14992 ( .A(top_core_EC_mc_n182), .B(top_core_EC_mc_n183), .Y(
        top_core_EC_mc_n179) );
  XNOR2X1 U14993 ( .A(top_core_EC_mix_in[64]), .B(top_core_EC_mix_in[72]), .Y(
        top_core_EC_mc_n182) );
  XNOR2X1 U14994 ( .A(top_core_EC_mc_n174), .B(top_core_EC_mc_n175), .Y(
        top_core_EC_mc_n171) );
  XNOR2X1 U14995 ( .A(top_core_EC_mc_mix_in_2_66_), .B(
        top_core_EC_mc_mix_in_2_74_), .Y(top_core_EC_mc_n174) );
  XNOR2X1 U14996 ( .A(top_core_EC_mc_n166), .B(top_core_EC_mc_n167), .Y(
        top_core_EC_mc_n163) );
  XNOR2X1 U14997 ( .A(top_core_EC_mix_in[66]), .B(top_core_EC_mix_in[74]), .Y(
        top_core_EC_mc_n166) );
  XNOR2X1 U14998 ( .A(top_core_EC_mc_n158), .B(top_core_EC_mc_n159), .Y(
        top_core_EC_mc_n155) );
  XNOR2X1 U14999 ( .A(top_core_EC_mix_in[67]), .B(top_core_EC_mix_in[75]), .Y(
        top_core_EC_mc_n158) );
  XNOR2X1 U15000 ( .A(top_core_EC_mc_n150), .B(top_core_EC_mc_n151), .Y(
        top_core_EC_mc_n147) );
  XNOR2X1 U15001 ( .A(top_core_EC_mc_mix_in_8[71]), .B(
        top_core_EC_mc_mix_in_8[79]), .Y(top_core_EC_mc_n150) );
  XNOR2X1 U15002 ( .A(top_core_EC_mc_n142), .B(top_core_EC_mc_n143), .Y(
        top_core_EC_mc_n139) );
  XNOR2X1 U15003 ( .A(top_core_EC_mc_mix_in_8[64]), .B(n1538), .Y(
        top_core_EC_mc_n142) );
  XNOR2X1 U15004 ( .A(top_core_EC_mc_n134), .B(top_core_EC_mc_n135), .Y(
        top_core_EC_mc_n131) );
  XNOR2X1 U15005 ( .A(top_core_EC_mc_mix_in_4_64_), .B(n1537), .Y(
        top_core_EC_mc_n134) );
  XNOR2X1 U15006 ( .A(top_core_EC_mc_n126), .B(top_core_EC_mc_n127), .Y(
        top_core_EC_mc_n123) );
  XNOR2X1 U15007 ( .A(top_core_EC_mc_mix_in_2_64_), .B(n1536), .Y(
        top_core_EC_mc_n126) );
  XNOR2X1 U15008 ( .A(top_core_EC_mc_n45), .B(top_core_EC_mc_n46), .Y(
        top_core_EC_mc_n42) );
  XNOR2X1 U15009 ( .A(top_core_EC_mix_in[112]), .B(n1554), .Y(
        top_core_EC_mc_n45) );
  XNOR2X1 U15010 ( .A(top_core_EC_mc_n36), .B(top_core_EC_mc_n37), .Y(
        top_core_EC_mc_n33) );
  XNOR2X1 U15011 ( .A(top_core_EC_mc_mix_in_2_114_), .B(
        top_core_EC_mc_mix_in_4_106_), .Y(top_core_EC_mc_n36) );
  XNOR2X1 U15012 ( .A(top_core_EC_mc_n27), .B(top_core_EC_mc_n28), .Y(
        top_core_EC_mc_n24) );
  XNOR2X1 U15013 ( .A(top_core_EC_mix_in[114]), .B(
        top_core_EC_mc_mix_in_2_106_), .Y(top_core_EC_mc_n27) );
  XNOR2X1 U15014 ( .A(top_core_EC_mc_n18), .B(top_core_EC_mc_n19), .Y(
        top_core_EC_mc_n15) );
  XNOR2X1 U15015 ( .A(top_core_EC_mix_in[115]), .B(
        top_core_EC_mc_mix_in_2_107_), .Y(top_core_EC_mc_n18) );
  XNOR2X1 U15016 ( .A(top_core_EC_mc_n809), .B(top_core_EC_mc_n810), .Y(
        top_core_EC_mc_n806) );
  XNOR2X1 U15017 ( .A(top_core_EC_mc_mix_in_8[103]), .B(
        top_core_EC_mc_mix_in_8[111]), .Y(top_core_EC_mc_n809) );
  XNOR2X1 U15018 ( .A(top_core_EC_mc_n801), .B(top_core_EC_mc_n802), .Y(
        top_core_EC_mc_n798) );
  XNOR2X1 U15019 ( .A(top_core_EC_mc_mix_in_8[96]), .B(n1556), .Y(
        top_core_EC_mc_n801) );
  XNOR2X1 U15020 ( .A(top_core_EC_mc_n793), .B(top_core_EC_mc_n794), .Y(
        top_core_EC_mc_n790) );
  XNOR2X1 U15021 ( .A(top_core_EC_mc_mix_in_4_96_), .B(n1555), .Y(
        top_core_EC_mc_n793) );
  XNOR2X1 U15022 ( .A(top_core_EC_mc_n785), .B(top_core_EC_mc_n786), .Y(
        top_core_EC_mc_n782) );
  XNOR2X1 U15023 ( .A(top_core_EC_mc_mix_in_2_96_), .B(n1554), .Y(
        top_core_EC_mc_n785) );
  XOR2X1 U15024 ( .A(n1552), .B(n1551), .Y(top_core_EC_mc_mix_in_8[122]) );
  XOR2X1 U15025 ( .A(n1540), .B(n1543), .Y(top_core_EC_mc_n376) );
  XOR2X1 U15026 ( .A(n1534), .B(n1537), .Y(top_core_EC_mc_n117) );
  XOR2X1 U15027 ( .A(n1552), .B(n1555), .Y(top_core_EC_mc_n770) );
  XOR2X1 U15028 ( .A(n1553), .B(n1556), .Y(top_core_EC_mc_n717) );
  XOR2X1 U15029 ( .A(n1541), .B(n1544), .Y(top_core_EC_mc_n311) );
  XOR2X1 U15030 ( .A(n1535), .B(n1538), .Y(top_core_EC_mc_n52) );
  NAND2X1 U15031 ( .A(n11839), .B(n1802), .Y(n11875) );
  NAND2X1 U15032 ( .A(top_core_KE_sb1_n268), .B(n1823), .Y(
        top_core_KE_sb1_n304) );
  NAND2X1 U15033 ( .A(n12470), .B(n1760), .Y(n12506) );
  NAND2X1 U15034 ( .A(n12155), .B(n1781), .Y(n12191) );
  NAND2X1 U15035 ( .A(n13730), .B(n1651), .Y(n13766) );
  NAND2X1 U15036 ( .A(n13415), .B(n1680), .Y(n13451) );
  NAND2X1 U15037 ( .A(n12785), .B(n1738), .Y(n12821) );
  NAND2X1 U15038 ( .A(n13100), .B(n1709), .Y(n13136) );
  XOR2X1 U15039 ( .A(n1537), .B(n1536), .Y(top_core_EC_mc_mix_in_8[74]) );
  XOR2X1 U15040 ( .A(n1537), .B(top_core_EC_mc_mix_in_2_75_), .Y(
        top_core_EC_mc_mix_in_8[77]) );
  XOR2X1 U15041 ( .A(n1555), .B(top_core_EC_mc_mix_in_2_107_), .Y(
        top_core_EC_mc_mix_in_8[109]) );
  NAND2X1 U15042 ( .A(n1203), .B(n6830), .Y(n11883) );
  NAND2X1 U15043 ( .A(n1194), .B(n6809), .Y(top_core_KE_sb1_n312) );
  NAND2X1 U15044 ( .A(n1163), .B(n6534), .Y(n12514) );
  NAND2X1 U15045 ( .A(n1154), .B(n6512), .Y(n12199) );
  NAND2X1 U15046 ( .A(n1149), .B(n6477), .Y(n13459) );
  NAND2X1 U15047 ( .A(n1189), .B(n6780), .Y(n12829) );
  NAND2X1 U15048 ( .A(n1158), .B(n6523), .Y(n13774) );
  NAND2X1 U15049 ( .A(n1198), .B(n6819), .Y(n13144) );
  INVX1 U15050 ( .A(n11879), .Y(n6922) );
  INVX1 U15051 ( .A(top_core_KE_sb1_n308), .Y(n6876) );
  INVX1 U15052 ( .A(n12510), .Y(n6629) );
  INVX1 U15053 ( .A(n12195), .Y(n6582) );
  OAI22X1 U15054 ( .A0(n2848), .A1(n17085), .B0(n17086), .B1(n17087), .Y(
        n17079) );
  AOI211X1 U15055 ( .A0(n5378), .A1(n2901), .B0(n17088), .C0(n17089), .Y(
        n17086) );
  OAI21XL U15056 ( .A0(n1309), .A1(n17090), .B0(n17091), .Y(n17089) );
  OAI22X1 U15057 ( .A0(n3449), .A1(n13935), .B0(n13936), .B1(n13937), .Y(
        n13929) );
  AOI211X1 U15058 ( .A0(n6149), .A1(n3506), .B0(n13938), .C0(n13939), .Y(
        n13936) );
  OAI21XL U15059 ( .A0(n1279), .A1(n13940), .B0(n13941), .Y(n13939) );
  OAI22X1 U15060 ( .A0(n2606), .A1(n18345), .B0(n18346), .B1(n18347), .Y(
        n18339) );
  AOI211X1 U15061 ( .A0(n5024), .A1(n2655), .B0(n18348), .C0(n18349), .Y(
        n18346) );
  OAI21XL U15062 ( .A0(n1321), .A1(n18350), .B0(n18351), .Y(n18349) );
  OAI22X1 U15063 ( .A0(n3208), .A1(n15195), .B0(n15196), .B1(n15197), .Y(
        n15189) );
  AOI211X1 U15064 ( .A0(n5850), .A1(n3261), .B0(n15198), .C0(n15199), .Y(
        n15196) );
  OAI21XL U15065 ( .A0(n1291), .A1(n15200), .B0(n15201), .Y(n15199) );
  OAI22X1 U15066 ( .A0(n3147), .A1(n15510), .B0(n15511), .B1(n15512), .Y(
        n15504) );
  AOI211X1 U15067 ( .A0(n5766), .A1(n3200), .B0(n15513), .C0(n15514), .Y(
        n15511) );
  OAI21XL U15068 ( .A0(n1294), .A1(n15515), .B0(n15516), .Y(n15514) );
  OAI22X1 U15069 ( .A0(n2545), .A1(n18660), .B0(n18661), .B1(n18662), .Y(
        n18654) );
  AOI211X1 U15070 ( .A0(n4908), .A1(n2594), .B0(n18663), .C0(n18664), .Y(
        n18661) );
  OAI21XL U15071 ( .A0(n1324), .A1(n18665), .B0(n18666), .Y(n18664) );
  OAI22X1 U15072 ( .A0(n2909), .A1(n16770), .B0(n16771), .B1(n16772), .Y(
        n16764) );
  AOI211X1 U15073 ( .A0(n5462), .A1(n2962), .B0(n16773), .C0(n16774), .Y(
        n16771) );
  OAI21XL U15074 ( .A0(n1306), .A1(n16775), .B0(n16776), .Y(n16774) );
  OAI22X1 U15075 ( .A0(n3269), .A1(n14880), .B0(n14881), .B1(n14882), .Y(
        n14874) );
  AOI211X1 U15076 ( .A0(n5926), .A1(n3315), .B0(n14883), .C0(n14884), .Y(
        n14881) );
  OAI21XL U15077 ( .A0(n1288), .A1(n14885), .B0(n14886), .Y(n14884) );
  OAI22X1 U15078 ( .A0(n2970), .A1(n16455), .B0(n16456), .B1(n16457), .Y(
        n16449) );
  AOI211X1 U15079 ( .A0(n5538), .A1(n3019), .B0(n16458), .C0(n16459), .Y(
        n16456) );
  OAI21XL U15080 ( .A0(n1303), .A1(n16460), .B0(n16461), .Y(n16459) );
  OAI22X1 U15081 ( .A0(n2667), .A1(n18030), .B0(n18031), .B1(n18032), .Y(
        n18024) );
  AOI211X1 U15082 ( .A0(n5108), .A1(n2723), .B0(n18033), .C0(n18034), .Y(
        n18031) );
  OAI21XL U15083 ( .A0(n1318), .A1(n18035), .B0(n18036), .Y(n18034) );
  OAI22X1 U15084 ( .A0(n3330), .A1(n14565), .B0(n14566), .B1(n14567), .Y(
        n14559) );
  AOI211X1 U15085 ( .A0(n6002), .A1(n3379), .B0(n14568), .C0(n14569), .Y(
        n14566) );
  OAI21XL U15086 ( .A0(n1285), .A1(n14570), .B0(n14571), .Y(n14569) );
  OAI22X1 U15087 ( .A0(n3028), .A1(n16140), .B0(n16141), .B1(n16142), .Y(
        n16134) );
  AOI211X1 U15088 ( .A0(n5614), .A1(n3077), .B0(n16143), .C0(n16144), .Y(
        n16141) );
  OAI21XL U15089 ( .A0(n1300), .A1(n16145), .B0(n16146), .Y(n16144) );
  OAI22X1 U15090 ( .A0(n2727), .A1(n17715), .B0(n17716), .B1(n17717), .Y(
        n17709) );
  AOI211X1 U15091 ( .A0(n5216), .A1(n2778), .B0(n17718), .C0(n17719), .Y(
        n17716) );
  OAI21XL U15092 ( .A0(n1315), .A1(n17720), .B0(n17721), .Y(n17719) );
  OAI22X1 U15093 ( .A0(n3388), .A1(n14250), .B0(n14251), .B1(n14252), .Y(
        n14244) );
  AOI211X1 U15094 ( .A0(n6078), .A1(n3445), .B0(n14253), .C0(n14254), .Y(
        n14251) );
  OAI21XL U15095 ( .A0(n1282), .A1(n14255), .B0(n14256), .Y(n14254) );
  OAI22X1 U15096 ( .A0(n3089), .A1(n15825), .B0(n15826), .B1(n15827), .Y(
        n15819) );
  AOI211X1 U15097 ( .A0(n5690), .A1(n3138), .B0(n15828), .C0(n15829), .Y(
        n15826) );
  OAI21XL U15098 ( .A0(n1297), .A1(n15830), .B0(n15831), .Y(n15829) );
  OAI22X1 U15099 ( .A0(n2788), .A1(n17400), .B0(n17401), .B1(n17402), .Y(
        n17394) );
  AOI211X1 U15100 ( .A0(n5294), .A1(n2838), .B0(n17403), .C0(n17404), .Y(
        n17401) );
  OAI21XL U15101 ( .A0(n1312), .A1(n17405), .B0(n17406), .Y(n17404) );
  XOR2X1 U15102 ( .A(top_core_EC_mc_mix_in_4_96_), .B(
        top_core_EC_mc_mix_in_2_96_), .Y(top_core_EC_mc_mix_in_8[98]) );
  NAND2X1 U15103 ( .A(n1802), .B(n11712), .Y(n11676) );
  NAND2X1 U15104 ( .A(n1823), .B(top_core_KE_sb1_n138), .Y(
        top_core_KE_sb1_n101) );
  NAND2X1 U15105 ( .A(n1760), .B(n12343), .Y(n12307) );
  NAND2X1 U15106 ( .A(n1680), .B(n13289), .Y(n13253) );
  NAND2X1 U15107 ( .A(n1781), .B(n12028), .Y(n11992) );
  NAND2X1 U15108 ( .A(n1709), .B(n12974), .Y(n12938) );
  NAND2X1 U15109 ( .A(n1651), .B(n13604), .Y(n13568) );
  NAND2X1 U15110 ( .A(n1738), .B(n12659), .Y(n12623) );
  NAND2X1 U15111 ( .A(n6552), .B(n1687), .Y(n13301) );
  NAND2X1 U15112 ( .A(n6847), .B(n1745), .Y(n12671) );
  NAND2X1 U15113 ( .A(n6893), .B(n1716), .Y(n12986) );
  NAND2X1 U15114 ( .A(n6914), .B(n1222), .Y(n11725) );
  NAND2X1 U15115 ( .A(n6868), .B(n1216), .Y(top_core_KE_sb1_n152) );
  NAND2X1 U15116 ( .A(n6621), .B(n1181), .Y(n12356) );
  NAND2X1 U15117 ( .A(n6574), .B(n1176), .Y(n12041) );
  NAND2X1 U15118 ( .A(n6917), .B(n1809), .Y(n11724) );
  NAND2X1 U15119 ( .A(n6871), .B(n1830), .Y(top_core_KE_sb1_n151) );
  NAND2X1 U15120 ( .A(n6624), .B(n1767), .Y(n12355) );
  NAND2X1 U15121 ( .A(n6577), .B(n1788), .Y(n12040) );
  NAND2X1 U15122 ( .A(n6600), .B(n1658), .Y(n13616) );
  CLKINVX3 U15123 ( .A(n12290), .Y(n6616) );
  AOI22XL U15124 ( .A0(n11712), .A1(n1259), .B0(n11827), .B1(n681), .Y(n11911)
         );
  AOI22XL U15125 ( .A0(top_core_KE_sb1_n138), .A1(n1331), .B0(
        top_core_KE_sb1_n256), .B1(n682), .Y(top_core_KE_sb1_n340) );
  AOI22XL U15126 ( .A0(n12343), .A1(n1266), .B0(n12458), .B1(n683), .Y(n12542)
         );
  AOI22XL U15127 ( .A0(n12028), .A1(n1262), .B0(n12143), .B1(n684), .Y(n12227)
         );
  AOI22XL U15128 ( .A0(n12659), .A1(n1269), .B0(n12773), .B1(n688), .Y(n12857)
         );
  AOI22XL U15129 ( .A0(n13604), .A1(n1278), .B0(n13718), .B1(n685), .Y(n13802)
         );
  AOI22XL U15130 ( .A0(n12974), .A1(n1272), .B0(n13088), .B1(n687), .Y(n13172)
         );
  AOI22X1 U15131 ( .A0(n17153), .A1(n337), .B0(n5390), .B1(n2877), .Y(n17226)
         );
  AOI22X1 U15132 ( .A0(n14003), .A1(n338), .B0(n6172), .B1(n3474), .Y(n14076)
         );
  AOI22X1 U15133 ( .A0(n15263), .A1(n340), .B0(n5862), .B1(n3237), .Y(n15336)
         );
  AOI22X1 U15134 ( .A0(n18413), .A1(n339), .B0(n5036), .B1(n2635), .Y(n18486)
         );
  AOI22X1 U15135 ( .A0(n15578), .A1(n341), .B0(n5778), .B1(n3176), .Y(n15651)
         );
  AOI22X1 U15136 ( .A0(n16838), .A1(n342), .B0(n5474), .B1(n2934), .Y(n16911)
         );
  AOI22X1 U15137 ( .A0(n18728), .A1(n343), .B0(n4920), .B1(n2574), .Y(n18801)
         );
  AOI22X1 U15138 ( .A0(n14948), .A1(n344), .B0(n5938), .B1(n3297), .Y(n15021)
         );
  AOI22X1 U15139 ( .A0(n16523), .A1(n345), .B0(n5550), .B1(n2995), .Y(n16596)
         );
  AOI22X1 U15140 ( .A0(n18098), .A1(n346), .B0(n5120), .B1(n2692), .Y(n18171)
         );
  AOI22X1 U15141 ( .A0(n14633), .A1(n347), .B0(n6014), .B1(n3359), .Y(n14706)
         );
  AOI22X1 U15142 ( .A0(n16208), .A1(n348), .B0(n5626), .B1(n3057), .Y(n16281)
         );
  AOI22X1 U15143 ( .A0(n17783), .A1(n349), .B0(n5228), .B1(n2756), .Y(n17856)
         );
  AOI22X1 U15144 ( .A0(n14318), .A1(n350), .B0(n6090), .B1(n3413), .Y(n14391)
         );
  AOI22X1 U15145 ( .A0(n15893), .A1(n351), .B0(n5702), .B1(n3118), .Y(n15966)
         );
  AOI22X1 U15146 ( .A0(n17468), .A1(n352), .B0(n5306), .B1(n2816), .Y(n17541)
         );
  XNOR2X1 U15147 ( .A(top_core_EC_mc_mix_in_8[63]), .B(top_core_EC_mc_n400), 
        .Y(top_core_EC_mc_n324) );
  XNOR2X1 U15148 ( .A(top_core_EC_mc_mix_in_8[95]), .B(top_core_EC_mc_n141), 
        .Y(top_core_EC_mc_n65) );
  XNOR2X1 U15149 ( .A(top_core_EC_mc_mix_in_8[127]), .B(top_core_EC_mc_n800), 
        .Y(top_core_EC_mc_n730) );
  XNOR2X1 U15150 ( .A(top_core_EC_mc_mix_in_2_90_), .B(top_core_EC_mc_n165), 
        .Y(top_core_EC_mc_n89) );
  XNOR2X1 U15151 ( .A(top_core_EC_mc_mix_in_2_122_), .B(top_core_EC_mc_n26), 
        .Y(top_core_EC_mc_n753) );
  AOI22X1 U15152 ( .A0(n5319), .A1(n10146), .B0(n5318), .B1(n10147), .Y(n10145) );
  INVX1 U15153 ( .A(n10092), .Y(n5319) );
  INVX1 U15154 ( .A(n10090), .Y(n5318) );
  AOI22X1 U15155 ( .A0(n6104), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n332), 
        .B0(n6103), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n333), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n331) );
  INVX1 U15156 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n278), .Y(n6104) );
  INVX1 U15157 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n276), .Y(n6103) );
  AOI22X1 U15158 ( .A0(n5791), .A1(n8394), .B0(n5790), .B1(n8395), .Y(n8393)
         );
  INVX1 U15159 ( .A(n8340), .Y(n5791) );
  INVX1 U15160 ( .A(n8338), .Y(n5790) );
  AOI22X1 U15161 ( .A0(n4965), .A1(n11314), .B0(n4964), .B1(n11315), .Y(n11313) );
  INVX1 U15162 ( .A(n11260), .Y(n4965) );
  INVX1 U15163 ( .A(n11258), .Y(n4964) );
  AOI22X1 U15164 ( .A0(n5049), .A1(n11022), .B0(n5048), .B1(n11023), .Y(n11021) );
  INVX1 U15165 ( .A(n10968), .Y(n5049) );
  INVX1 U15166 ( .A(n10966), .Y(n5048) );
  AOI22X1 U15167 ( .A0(n6019), .A1(n7518), .B0(n6018), .B1(n7519), .Y(n7517)
         );
  INVX1 U15168 ( .A(n7464), .Y(n6019) );
  INVX1 U15169 ( .A(n7462), .Y(n6018) );
  AOI22X1 U15170 ( .A0(n5555), .A1(n9270), .B0(n5554), .B1(n9271), .Y(n9269)
         );
  INVX1 U15171 ( .A(n9216), .Y(n5555) );
  INVX1 U15172 ( .A(n9214), .Y(n5554) );
  AOI22X1 U15173 ( .A0(n5235), .A1(n10438), .B0(n5234), .B1(n10439), .Y(n10437) );
  INVX1 U15174 ( .A(n10384), .Y(n5235) );
  INVX1 U15175 ( .A(n10382), .Y(n5234) );
  AOI22X1 U15176 ( .A0(n5479), .A1(n9562), .B0(n5478), .B1(n9563), .Y(n9561)
         );
  INVX1 U15177 ( .A(n9508), .Y(n5479) );
  INVX1 U15178 ( .A(n9506), .Y(n5478) );
  AOI22X1 U15179 ( .A0(n5707), .A1(n8686), .B0(n5706), .B1(n8687), .Y(n8685)
         );
  INVX1 U15180 ( .A(n8632), .Y(n5707) );
  INVX1 U15181 ( .A(n8630), .Y(n5706) );
  AOI22X1 U15182 ( .A0(n5943), .A1(n7810), .B0(n5942), .B1(n7811), .Y(n7809)
         );
  INVX1 U15183 ( .A(n7756), .Y(n5943) );
  INVX1 U15184 ( .A(n7754), .Y(n5942) );
  AOI22X1 U15185 ( .A0(n4844), .A1(n11606), .B0(n4843), .B1(n11607), .Y(n11605) );
  INVX1 U15186 ( .A(n11552), .Y(n4844) );
  INVX1 U15187 ( .A(n11550), .Y(n4843) );
  AOI22X1 U15188 ( .A0(n5157), .A1(n10730), .B0(n5156), .B1(n10731), .Y(n10729) );
  INVX1 U15189 ( .A(n10676), .Y(n5157) );
  INVX1 U15190 ( .A(n10674), .Y(n5156) );
  AOI22X1 U15191 ( .A0(n5398), .A1(n9854), .B0(n5397), .B1(n9855), .Y(n9853)
         );
  INVX1 U15192 ( .A(n9800), .Y(n5398) );
  INVX1 U15193 ( .A(n9798), .Y(n5397) );
  AOI22X1 U15194 ( .A0(n5631), .A1(n8978), .B0(n5630), .B1(n8979), .Y(n8977)
         );
  INVX1 U15195 ( .A(n8924), .Y(n5631) );
  INVX1 U15196 ( .A(n8922), .Y(n5630) );
  AOI22X1 U15197 ( .A0(n5867), .A1(n8102), .B0(n5866), .B1(n8103), .Y(n8101)
         );
  INVX1 U15198 ( .A(n8048), .Y(n5867) );
  INVX1 U15199 ( .A(n8046), .Y(n5866) );
  XNOR2X1 U15200 ( .A(n1539), .B(top_core_EC_mc_n449), .Y(top_core_EC_mc_n373)
         );
  XNOR2X1 U15201 ( .A(n1541), .B(top_core_EC_mc_n392), .Y(top_core_EC_mc_n316)
         );
  XNOR2X1 U15202 ( .A(n1540), .B(top_core_EC_mc_n384), .Y(top_core_EC_mc_n308)
         );
  XNOR2X1 U15203 ( .A(n1533), .B(top_core_EC_mc_n181), .Y(top_core_EC_mc_n114)
         );
  XNOR2X1 U15204 ( .A(n1535), .B(top_core_EC_mc_n133), .Y(top_core_EC_mc_n57)
         );
  XNOR2X1 U15205 ( .A(n1534), .B(top_core_EC_mc_n125), .Y(top_core_EC_mc_n49)
         );
  XNOR2X1 U15206 ( .A(n1551), .B(top_core_EC_mc_n44), .Y(top_core_EC_mc_n767)
         );
  XNOR2X1 U15207 ( .A(n1553), .B(top_core_EC_mc_n792), .Y(top_core_EC_mc_n722)
         );
  XNOR2X1 U15208 ( .A(n1552), .B(top_core_EC_mc_n784), .Y(top_core_EC_mc_n714)
         );
  XOR2X1 U15209 ( .A(n1540), .B(n1539), .Y(top_core_EC_mc_mix_in_8[58]) );
  XOR2X1 U15210 ( .A(n1540), .B(top_core_EC_mc_mix_in_2_59_), .Y(
        top_core_EC_mc_mix_in_8[61]) );
  XOR2X1 U15211 ( .A(n1534), .B(n1533), .Y(top_core_EC_mc_mix_in_8[90]) );
  XOR2X1 U15212 ( .A(n1534), .B(top_core_EC_mc_mix_in_2_91_), .Y(
        top_core_EC_mc_mix_in_8[93]) );
  XOR2X1 U15213 ( .A(n1552), .B(top_core_EC_mc_mix_in_2_123_), .Y(
        top_core_EC_mc_mix_in_8[125]) );
  NAND2XL U15214 ( .A(n76), .B(n13697), .Y(n13533) );
  CLKINVX3 U15215 ( .A(n12305), .Y(n6530) );
  OAI21XL U15216 ( .A0(n9951), .A1(n9952), .B0(n2856), .Y(n9939) );
  OAI221XL U15217 ( .A0(n1245), .A1(n9918), .B0(n2882), .B1(n9943), .C0(n9953), 
        .Y(n9952) );
  AOI21X1 U15218 ( .A0(n353), .A1(n9954), .B0(n5364), .Y(n9953) );
  OAI21XL U15219 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n136), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n137), .B0(n3461), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n124) );
  OAI221XL U15220 ( .A0(n1327), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n102), 
        .B0(n3483), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n128), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n138), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n137) );
  AOI21X1 U15221 ( .A0(n354), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n139), 
        .B0(n6154), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n138) );
  OAI21XL U15222 ( .A0(n11119), .A1(n11120), .B0(n2620), .Y(n11107) );
  OAI221XL U15223 ( .A0(n1253), .A1(n11086), .B0(n2640), .B1(n11111), .C0(
        n11121), .Y(n11120) );
  AOI21X1 U15224 ( .A0(n356), .A1(n11122), .B0(n5010), .Y(n11121) );
  OAI21XL U15225 ( .A0(n8199), .A1(n8200), .B0(n3216), .Y(n8187) );
  OAI221XL U15226 ( .A0(n1233), .A1(n8166), .B0(n3242), .B1(n8191), .C0(n8201), 
        .Y(n8200) );
  AOI21X1 U15227 ( .A0(n355), .A1(n8202), .B0(n5836), .Y(n8201) );
  OAI21XL U15228 ( .A0(n10827), .A1(n10828), .B0(n2675), .Y(n10815) );
  OAI221XL U15229 ( .A0(n1251), .A1(n10794), .B0(n2701), .B1(n10819), .C0(
        n10829), .Y(n10828) );
  AOI21X1 U15230 ( .A0(n357), .A1(n10830), .B0(n5094), .Y(n10829) );
  OAI21XL U15231 ( .A0(n9075), .A1(n9076), .B0(n3042), .Y(n9063) );
  OAI221XL U15232 ( .A0(n1239), .A1(n9042), .B0(n3062), .B1(n9067), .C0(n9077), 
        .Y(n9076) );
  AOI21X1 U15233 ( .A0(n359), .A1(n9078), .B0(n5600), .Y(n9077) );
  OAI21XL U15234 ( .A0(n7323), .A1(n7324), .B0(n3402), .Y(n7311) );
  OAI221XL U15235 ( .A0(n1227), .A1(n7290), .B0(n3422), .B1(n7315), .C0(n7325), 
        .Y(n7324) );
  AOI21X1 U15236 ( .A0(n358), .A1(n7326), .B0(n6064), .Y(n7325) );
  OAI21XL U15237 ( .A0(n10243), .A1(n10244), .B0(n2802), .Y(n10231) );
  OAI221XL U15238 ( .A0(n1247), .A1(n10210), .B0(n2822), .B1(n10235), .C0(
        n10245), .Y(n10244) );
  AOI21X1 U15239 ( .A0(n360), .A1(n10246), .B0(n5280), .Y(n10245) );
  OAI21XL U15240 ( .A0(n9367), .A1(n9368), .B0(n2984), .Y(n9355) );
  OAI221XL U15241 ( .A0(n1241), .A1(n9334), .B0(n3004), .B1(n9359), .C0(n9369), 
        .Y(n9368) );
  AOI21X1 U15242 ( .A0(n361), .A1(n9370), .B0(n5524), .Y(n9369) );
  OAI21XL U15243 ( .A0(n8491), .A1(n8492), .B0(n3161), .Y(n8479) );
  OAI221XL U15244 ( .A0(n1235), .A1(n8458), .B0(n3181), .B1(n8483), .C0(n8493), 
        .Y(n8492) );
  AOI21X1 U15245 ( .A0(n362), .A1(n8494), .B0(n5752), .Y(n8493) );
  OAI21XL U15246 ( .A0(n7615), .A1(n7616), .B0(n3344), .Y(n7603) );
  OAI221XL U15247 ( .A0(n1229), .A1(n7582), .B0(n3364), .B1(n7607), .C0(n7617), 
        .Y(n7616) );
  AOI21X1 U15248 ( .A0(n363), .A1(n7618), .B0(n5988), .Y(n7617) );
  OAI21XL U15249 ( .A0(n11411), .A1(n11412), .B0(n2558), .Y(n11399) );
  OAI221XL U15250 ( .A0(n1255), .A1(n11378), .B0(n2579), .B1(n11403), .C0(
        n11413), .Y(n11412) );
  AOI21X1 U15251 ( .A0(n364), .A1(n11414), .B0(n4894), .Y(n11413) );
  OAI21XL U15252 ( .A0(n10535), .A1(n10536), .B0(n2735), .Y(n10523) );
  OAI221XL U15253 ( .A0(n1249), .A1(n10502), .B0(n2761), .B1(n10527), .C0(
        n10537), .Y(n10536) );
  AOI21X1 U15254 ( .A0(n365), .A1(n10538), .B0(n5202), .Y(n10537) );
  OAI21XL U15255 ( .A0(n9659), .A1(n9660), .B0(n2923), .Y(n9647) );
  OAI221XL U15256 ( .A0(n1243), .A1(n9626), .B0(n2943), .B1(n9651), .C0(n9661), 
        .Y(n9660) );
  AOI21X1 U15257 ( .A0(n366), .A1(n9662), .B0(n5448), .Y(n9661) );
  OAI21XL U15258 ( .A0(n8783), .A1(n8784), .B0(n3097), .Y(n8771) );
  OAI221XL U15259 ( .A0(n1237), .A1(n8750), .B0(n3123), .B1(n8775), .C0(n8785), 
        .Y(n8784) );
  AOI21X1 U15260 ( .A0(n367), .A1(n8786), .B0(n5676), .Y(n8785) );
  OAI21XL U15261 ( .A0(n7907), .A1(n7908), .B0(n3283), .Y(n7895) );
  OAI221XL U15262 ( .A0(n1231), .A1(n7874), .B0(n3303), .B1(n7899), .C0(n7909), 
        .Y(n7908) );
  AOI21X1 U15263 ( .A0(n368), .A1(n7910), .B0(n5912), .Y(n7909) );
  AOI21X1 U15264 ( .A0(n17099), .A1(n17006), .B0(n17035), .Y(n17097) );
  AOI21X1 U15265 ( .A0(n13949), .A1(n13856), .B0(n13885), .Y(n13947) );
  AOI21X1 U15266 ( .A0(n18359), .A1(n18266), .B0(n18295), .Y(n18357) );
  AOI21X1 U15267 ( .A0(n15209), .A1(n15116), .B0(n15145), .Y(n15207) );
  AOI21X1 U15268 ( .A0(n15524), .A1(n15431), .B0(n15460), .Y(n15522) );
  AOI21X1 U15269 ( .A0(n18674), .A1(n18581), .B0(n18610), .Y(n18672) );
  AOI21X1 U15270 ( .A0(n16784), .A1(n16691), .B0(n16720), .Y(n16782) );
  AOI21X1 U15271 ( .A0(n14894), .A1(n14801), .B0(n14830), .Y(n14892) );
  AOI21X1 U15272 ( .A0(n16469), .A1(n16376), .B0(n16405), .Y(n16467) );
  AOI21X1 U15273 ( .A0(n18044), .A1(n17951), .B0(n17980), .Y(n18042) );
  AOI21X1 U15274 ( .A0(n14579), .A1(n14486), .B0(n14515), .Y(n14577) );
  AOI21X1 U15275 ( .A0(n16154), .A1(n16061), .B0(n16090), .Y(n16152) );
  AOI21X1 U15276 ( .A0(n17729), .A1(n17636), .B0(n17665), .Y(n17727) );
  AOI21X1 U15277 ( .A0(n14264), .A1(n14171), .B0(n14200), .Y(n14262) );
  AOI21X1 U15278 ( .A0(n15839), .A1(n15746), .B0(n15775), .Y(n15837) );
  AOI21X1 U15279 ( .A0(n17414), .A1(n17321), .B0(n17350), .Y(n17412) );
  AOI21X1 U15280 ( .A0(n13869), .A1(n3493), .B0(n13870), .Y(n13865) );
  AOI21X1 U15281 ( .A0(n17019), .A1(n2892), .B0(n17020), .Y(n17015) );
  AOI21X1 U15282 ( .A0(n18279), .A1(top_core_EC_ss_in[112]), .B0(n18280), .Y(
        n18275) );
  AOI21X1 U15283 ( .A0(n15129), .A1(n3252), .B0(n15130), .Y(n15125) );
  AOI21X1 U15284 ( .A0(n15444), .A1(n3191), .B0(n15445), .Y(n15440) );
  AOI21X1 U15285 ( .A0(n18594), .A1(n2589), .B0(n18595), .Y(n18590) );
  AOI21X1 U15286 ( .A0(n16704), .A1(n2953), .B0(n16705), .Y(n16700) );
  AOI21X1 U15287 ( .A0(n14814), .A1(n3313), .B0(n14815), .Y(n14810) );
  AOI21X1 U15288 ( .A0(n16389), .A1(n3014), .B0(n16390), .Y(n16385) );
  AOI21X1 U15289 ( .A0(n17964), .A1(n2710), .B0(n17965), .Y(n17960) );
  AOI21X1 U15290 ( .A0(n14499), .A1(n3374), .B0(n14500), .Y(n14495) );
  AOI21X1 U15291 ( .A0(n16074), .A1(top_core_EC_ss_in[56]), .B0(n16075), .Y(
        n16070) );
  AOI21X1 U15292 ( .A0(n17649), .A1(n2771), .B0(n17650), .Y(n17645) );
  AOI21X1 U15293 ( .A0(n14184), .A1(n3432), .B0(n14185), .Y(n14180) );
  AOI21X1 U15294 ( .A0(n15759), .A1(n3133), .B0(n15760), .Y(n15755) );
  AOI21X1 U15295 ( .A0(n17334), .A1(n2832), .B0(n17335), .Y(n17330) );
  AOI21X1 U15296 ( .A0(n5330), .A1(n17122), .B0(n5328), .Y(n17115) );
  OAI21XL U15297 ( .A0(n481), .A1(n1000), .B0(n1309), .Y(n17122) );
  AOI21X1 U15298 ( .A0(n6114), .A1(n13972), .B0(n6112), .Y(n13965) );
  OAI21XL U15299 ( .A0(n482), .A1(n1140), .B0(n1279), .Y(n13972) );
  AOI21X1 U15300 ( .A0(n4976), .A1(n18382), .B0(n4974), .Y(n18375) );
  OAI21XL U15301 ( .A0(n483), .A1(n944), .B0(n1321), .Y(n18382) );
  AOI21X1 U15302 ( .A0(n5802), .A1(n15232), .B0(n5800), .Y(n15225) );
  OAI21XL U15303 ( .A0(n484), .A1(n1084), .B0(n1291), .Y(n15232) );
  AOI21X1 U15304 ( .A0(n5718), .A1(n15547), .B0(n5716), .Y(n15540) );
  OAI21XL U15305 ( .A0(n490), .A1(n1070), .B0(n1294), .Y(n15547) );
  AOI21X1 U15306 ( .A0(n4860), .A1(n18697), .B0(n4858), .Y(n18690) );
  OAI21XL U15307 ( .A0(n492), .A1(n930), .B0(n1324), .Y(n18697) );
  AOI21X1 U15308 ( .A0(n5414), .A1(n16807), .B0(n5412), .Y(n16800) );
  OAI21XL U15309 ( .A0(n494), .A1(n1014), .B0(n1306), .Y(n16807) );
  AOI21X1 U15310 ( .A0(n5878), .A1(n14917), .B0(n5876), .Y(n14910) );
  OAI21XL U15311 ( .A0(n496), .A1(n1098), .B0(n1288), .Y(n14917) );
  AOI21X1 U15312 ( .A0(n5490), .A1(n16492), .B0(n5488), .Y(n16485) );
  OAI21XL U15313 ( .A0(n489), .A1(n1028), .B0(n1303), .Y(n16492) );
  AOI21X1 U15314 ( .A0(n5060), .A1(n18067), .B0(n5058), .Y(n18060) );
  OAI21XL U15315 ( .A0(n485), .A1(n958), .B0(n1318), .Y(n18067) );
  AOI21X1 U15316 ( .A0(n5954), .A1(n14602), .B0(n5952), .Y(n14595) );
  OAI21XL U15317 ( .A0(n491), .A1(n1112), .B0(n1285), .Y(n14602) );
  AOI21X1 U15318 ( .A0(n5566), .A1(n16177), .B0(n5564), .Y(n16170) );
  OAI21XL U15319 ( .A0(n486), .A1(n1042), .B0(n1300), .Y(n16177) );
  AOI21X1 U15320 ( .A0(n5168), .A1(n17752), .B0(n5166), .Y(n17745) );
  OAI21XL U15321 ( .A0(n493), .A1(n972), .B0(n1315), .Y(n17752) );
  AOI21X1 U15322 ( .A0(n6030), .A1(n14287), .B0(n6028), .Y(n14280) );
  OAI21XL U15323 ( .A0(n487), .A1(n1126), .B0(n1282), .Y(n14287) );
  AOI21X1 U15324 ( .A0(n5642), .A1(n15862), .B0(n5640), .Y(n15855) );
  OAI21XL U15325 ( .A0(n495), .A1(n1056), .B0(n1297), .Y(n15862) );
  AOI21X1 U15326 ( .A0(n5246), .A1(n17437), .B0(n5244), .Y(n17430) );
  OAI21XL U15327 ( .A0(n488), .A1(n986), .B0(n1312), .Y(n17437) );
  OAI21XL U15328 ( .A0(n1651), .A1(n76), .B0(n13561), .Y(n13635) );
  AOI22XL U15329 ( .A0(n6904), .A1(n1222), .B0(n6914), .B1(n1259), .Y(n11897)
         );
  AOI22XL U15330 ( .A0(n6858), .A1(n1216), .B0(n6868), .B1(n1331), .Y(
        top_core_KE_sb1_n326) );
  AOI22XL U15331 ( .A0(n6611), .A1(n1181), .B0(n6621), .B1(n1266), .Y(n12528)
         );
  AOI22XL U15332 ( .A0(n6564), .A1(n1176), .B0(n6574), .B1(n1262), .Y(n12213)
         );
  AOI22X1 U15333 ( .A0(n10107), .A1(n2851), .B0(n2855), .B1(n10108), .Y(n10091) );
  OAI221XL U15334 ( .A0(n481), .A1(n9943), .B0(n1001), .B1(n9919), .C0(n10111), 
        .Y(n10107) );
  AOI222X1 U15335 ( .A0(n5366), .A1(top_core_EC_ss_in[80]), .B0(n465), .B1(
        n10081), .C0(n1615), .C1(n5350), .Y(n10110) );
  AOI22X1 U15336 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n293), .A1(n3452), 
        .B0(n3456), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n294), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n277) );
  OAI221XL U15337 ( .A0(n482), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n128), 
        .B0(n1143), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n104), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n297), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n293) );
  AOI222X1 U15338 ( .A0(n6156), .A1(top_core_EC_ss_in[0]), .B0(n466), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n267), .C0(n1625), .C1(n6146), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n296) );
  AOI22X1 U15339 ( .A0(n8355), .A1(n3211), .B0(n3215), .B1(n8356), .Y(n8339)
         );
  OAI221XL U15340 ( .A0(n484), .A1(n8191), .B0(n1085), .B1(n8167), .C0(n8359), 
        .Y(n8355) );
  AOI222X1 U15341 ( .A0(n5838), .A1(top_core_EC_ss_in[32]), .B0(n468), .B1(
        n8329), .C0(n1621), .C1(n5822), .Y(n8358) );
  AOI22X1 U15342 ( .A0(n11275), .A1(n2609), .B0(n2613), .B1(n11276), .Y(n11259) );
  OAI221XL U15343 ( .A0(n483), .A1(n11111), .B0(n945), .B1(n11087), .C0(n11279), .Y(n11275) );
  AOI222X1 U15344 ( .A0(n5012), .A1(n2651), .B0(n467), .B1(n11249), .C0(n1611), 
        .C1(n4996), .Y(n11278) );
  AOI22X1 U15345 ( .A0(n10983), .A1(n2670), .B0(n2674), .B1(n10984), .Y(n10967) );
  OAI221XL U15346 ( .A0(n485), .A1(n10819), .B0(n959), .B1(n10795), .C0(n10987), .Y(n10983) );
  AOI222X1 U15347 ( .A0(n5096), .A1(top_core_EC_ss_in[104]), .B0(n474), .B1(
        n10957), .C0(n1612), .C1(n5080), .Y(n10986) );
  AOI22X1 U15348 ( .A0(n7479), .A1(n3391), .B0(n3395), .B1(n7480), .Y(n7463)
         );
  OAI221XL U15349 ( .A0(n487), .A1(n7315), .B0(n1127), .B1(n7291), .C0(n7483), 
        .Y(n7479) );
  AOI222X1 U15350 ( .A0(n6066), .A1(top_core_EC_ss_in[8]), .B0(n478), .B1(
        n7453), .C0(n1624), .C1(n6050), .Y(n7482) );
  AOI22X1 U15351 ( .A0(n9231), .A1(n3031), .B0(n3035), .B1(n9232), .Y(n9215)
         );
  OAI221XL U15352 ( .A0(n486), .A1(n9067), .B0(n1043), .B1(n9043), .C0(n9235), 
        .Y(n9231) );
  AOI222X1 U15353 ( .A0(n5602), .A1(n3073), .B0(n476), .B1(n9205), .C0(n1618), 
        .C1(n5586), .Y(n9234) );
  AOI22X1 U15354 ( .A0(n10399), .A1(n2791), .B0(n2795), .B1(n10400), .Y(n10383) );
  OAI221XL U15355 ( .A0(n488), .A1(n10235), .B0(n987), .B1(n10211), .C0(n10403), .Y(n10399) );
  AOI222X1 U15356 ( .A0(n5282), .A1(n2834), .B0(n480), .B1(n10373), .C0(n1614), 
        .C1(n5266), .Y(n10402) );
  AOI22X1 U15357 ( .A0(n9523), .A1(n2973), .B0(n2977), .B1(n9524), .Y(n9507)
         );
  OAI221XL U15358 ( .A0(n489), .A1(n9359), .B0(n1029), .B1(n9335), .C0(n9527), 
        .Y(n9523) );
  AOI222X1 U15359 ( .A0(n5526), .A1(n3016), .B0(n473), .B1(n9497), .C0(n1617), 
        .C1(n5510), .Y(n9526) );
  AOI22X1 U15360 ( .A0(n8647), .A1(n3150), .B0(n3154), .B1(n8648), .Y(n8631)
         );
  OAI221XL U15361 ( .A0(n490), .A1(n8483), .B0(n1071), .B1(n8459), .C0(n8651), 
        .Y(n8647) );
  AOI222X1 U15362 ( .A0(n5754), .A1(top_core_EC_ss_in[40]), .B0(n469), .B1(
        n8621), .C0(n1620), .C1(n5738), .Y(n8650) );
  AOI22X1 U15363 ( .A0(n7771), .A1(n3333), .B0(n3337), .B1(n7772), .Y(n7755)
         );
  OAI221XL U15364 ( .A0(n491), .A1(n7607), .B0(n1113), .B1(n7583), .C0(n7775), 
        .Y(n7771) );
  AOI222X1 U15365 ( .A0(n5990), .A1(n3376), .B0(n475), .B1(n7745), .C0(n1623), 
        .C1(n5974), .Y(n7774) );
  AOI22X1 U15366 ( .A0(n11567), .A1(n2548), .B0(n2552), .B1(n11568), .Y(n11551) );
  OAI221XL U15367 ( .A0(n492), .A1(n11403), .B0(n931), .B1(n11379), .C0(n11571), .Y(n11567) );
  AOI222X1 U15368 ( .A0(n4896), .A1(n2590), .B0(n471), .B1(n11541), .C0(n1610), 
        .C1(n4880), .Y(n11570) );
  AOI22X1 U15369 ( .A0(n10691), .A1(n2730), .B0(n2734), .B1(n10692), .Y(n10675) );
  OAI221XL U15370 ( .A0(n493), .A1(n10527), .B0(n973), .B1(n10503), .C0(n10695), .Y(n10691) );
  AOI222X1 U15371 ( .A0(n5204), .A1(n2773), .B0(n477), .B1(n10665), .C0(n1613), 
        .C1(n5188), .Y(n10694) );
  AOI22X1 U15372 ( .A0(n9815), .A1(n2912), .B0(n2916), .B1(n9816), .Y(n9799)
         );
  OAI221XL U15373 ( .A0(n494), .A1(n9651), .B0(n1015), .B1(n9627), .C0(n9819), 
        .Y(n9815) );
  AOI222X1 U15374 ( .A0(n5450), .A1(top_core_EC_ss_in[72]), .B0(n470), .B1(
        n9789), .C0(n1616), .C1(n5434), .Y(n9818) );
  AOI22X1 U15375 ( .A0(n8939), .A1(n3092), .B0(n3096), .B1(n8940), .Y(n8923)
         );
  OAI221XL U15376 ( .A0(n495), .A1(n8775), .B0(n1057), .B1(n8751), .C0(n8943), 
        .Y(n8939) );
  AOI222X1 U15377 ( .A0(n5678), .A1(n3135), .B0(n479), .B1(n8913), .C0(n1619), 
        .C1(n5662), .Y(n8942) );
  AOI22X1 U15378 ( .A0(n8063), .A1(n3272), .B0(n3276), .B1(n8064), .Y(n8047)
         );
  OAI221XL U15379 ( .A0(n496), .A1(n7899), .B0(n1099), .B1(n7875), .C0(n8067), 
        .Y(n8063) );
  AOI222X1 U15380 ( .A0(n5914), .A1(top_core_EC_ss_in[24]), .B0(n472), .B1(
        n8037), .C0(n1622), .C1(n5898), .Y(n8066) );
  AOI21XL U15381 ( .A0(n13286), .A1(n13346), .B0(n6637), .Y(n13506) );
  INVX1 U15382 ( .A(n13444), .Y(n6637) );
  AOI21XL U15383 ( .A0(n12656), .A1(n12716), .B0(n6929), .Y(n12876) );
  INVX1 U15384 ( .A(n12814), .Y(n6929) );
  AOI21XL U15385 ( .A0(n13601), .A1(n13661), .B0(n6654), .Y(n13821) );
  INVX1 U15386 ( .A(n13759), .Y(n6654) );
  AOI21XL U15387 ( .A0(n12971), .A1(n13031), .B0(n6944), .Y(n13191) );
  INVX1 U15388 ( .A(n13129), .Y(n6944) );
  AOI21XL U15389 ( .A0(n1203), .A1(n11691), .B0(n11764), .Y(n11763) );
  AOI21XL U15390 ( .A0(n1194), .A1(top_core_KE_sb1_n116), .B0(
        top_core_KE_sb1_n192), .Y(top_core_KE_sb1_n191) );
  AOI21XL U15391 ( .A0(n1163), .A1(n12322), .B0(n12395), .Y(n12394) );
  AOI21XL U15392 ( .A0(n1149), .A1(n13268), .B0(n13341), .Y(n13340) );
  AOI21XL U15393 ( .A0(n1154), .A1(n12007), .B0(n12080), .Y(n12079) );
  AOI21XL U15394 ( .A0(n1189), .A1(n12638), .B0(n12711), .Y(n12710) );
  AOI21XL U15395 ( .A0(n1158), .A1(n13583), .B0(n13656), .Y(n13655) );
  AOI21XL U15396 ( .A0(n1198), .A1(n12953), .B0(n13026), .Y(n13025) );
  AOI21X1 U15397 ( .A0(n11704), .A1(n1815), .B0(n1205), .Y(n11762) );
  AOI21X1 U15398 ( .A0(top_core_KE_sb1_n129), .A1(n1836), .B0(n1196), .Y(
        top_core_KE_sb1_n190) );
  AOI21X1 U15399 ( .A0(n12335), .A1(n1772), .B0(n1165), .Y(n12393) );
  AOI21X1 U15400 ( .A0(n13281), .A1(n1689), .B0(n1152), .Y(n13339) );
  AOI21X1 U15401 ( .A0(n12020), .A1(n1794), .B0(n1156), .Y(n12078) );
  AOI21X1 U15402 ( .A0(n12651), .A1(n1747), .B0(n1192), .Y(n12709) );
  AOI21X1 U15403 ( .A0(n13596), .A1(n1661), .B0(n1161), .Y(n13654) );
  AOI21X1 U15404 ( .A0(n12966), .A1(n1718), .B0(n1201), .Y(n13024) );
  AOI2BB2X1 U15405 ( .B0(n6775), .B1(n12744), .A0N(n54), .A1N(n12609), .Y(
        n12856) );
  AOI2BB2X1 U15406 ( .B0(n6815), .B1(n13059), .A0N(n56), .A1N(n12924), .Y(
        n13171) );
  AOI22XL U15407 ( .A0(n753), .A1(n1811), .B0(n1203), .B1(n11705), .Y(n11899)
         );
  AOI22XL U15408 ( .A0(n754), .A1(n1832), .B0(n1194), .B1(top_core_KE_sb1_n130), .Y(top_core_KE_sb1_n328) );
  AOI22XL U15409 ( .A0(n752), .A1(n1769), .B0(n1163), .B1(n12336), .Y(n12530)
         );
  AOI22XL U15410 ( .A0(n748), .A1(n1691), .B0(n1149), .B1(n13282), .Y(n13475)
         );
  AOI22XL U15411 ( .A0(n755), .A1(n1790), .B0(n1154), .B1(n12021), .Y(n12215)
         );
  AOI22XL U15412 ( .A0(n749), .A1(n1749), .B0(n1189), .B1(n12652), .Y(n12845)
         );
  AOI22XL U15413 ( .A0(n751), .A1(n1661), .B0(n1158), .B1(n13597), .Y(n13790)
         );
  AOI22XL U15414 ( .A0(n750), .A1(n1720), .B0(n1198), .B1(n12967), .Y(n13160)
         );
  AOI2BB2X1 U15415 ( .B0(n1724), .B1(n12860), .A0N(n12622), .A1N(n694), .Y(
        n12858) );
  OAI22XL U15416 ( .A0(n1214), .A1(n181), .B0(n1747), .B1(n4), .Y(n12860) );
  AOI2BB2X1 U15417 ( .B0(n1695), .B1(n13175), .A0N(n12937), .A1N(n696), .Y(
        n13173) );
  OAI22XL U15418 ( .A0(n1220), .A1(n182), .B0(n1718), .B1(n5), .Y(n13175) );
  AOI21X1 U15419 ( .A0(n5320), .A1(n17178), .B0(n17179), .Y(n17177) );
  INVX1 U15420 ( .A(n16987), .Y(n5320) );
  NAND4BXL U15421 ( .AN(n17189), .B(n17041), .C(n17190), .D(n17191), .Y(n17178) );
  AOI31X1 U15422 ( .A0(n17180), .A1(n17181), .A2(n17182), .B0(n16989), .Y(
        n17179) );
  AOI21X1 U15423 ( .A0(n6101), .A1(n14028), .B0(n14029), .Y(n14027) );
  INVX1 U15424 ( .A(n13837), .Y(n6101) );
  NAND4BXL U15425 ( .AN(n14039), .B(n13891), .C(n14040), .D(n14041), .Y(n14028) );
  AOI31X1 U15426 ( .A0(n14030), .A1(n14031), .A2(n14032), .B0(n13839), .Y(
        n14029) );
  AOI21X1 U15427 ( .A0(n4966), .A1(n18438), .B0(n18439), .Y(n18437) );
  INVX1 U15428 ( .A(n18247), .Y(n4966) );
  NAND4BXL U15429 ( .AN(n18449), .B(n18301), .C(n18450), .D(n18451), .Y(n18438) );
  AOI31X1 U15430 ( .A0(n18440), .A1(n18441), .A2(n18442), .B0(n18249), .Y(
        n18439) );
  AOI21X1 U15431 ( .A0(n5792), .A1(n15288), .B0(n15289), .Y(n15287) );
  INVX1 U15432 ( .A(n15097), .Y(n5792) );
  NAND4BXL U15433 ( .AN(n15299), .B(n15151), .C(n15300), .D(n15301), .Y(n15288) );
  AOI31X1 U15434 ( .A0(n15290), .A1(n15291), .A2(n15292), .B0(n15099), .Y(
        n15289) );
  AOI21X1 U15435 ( .A0(n5708), .A1(n15603), .B0(n15604), .Y(n15602) );
  INVX1 U15436 ( .A(n15412), .Y(n5708) );
  NAND4BXL U15437 ( .AN(n15614), .B(n15466), .C(n15615), .D(n15616), .Y(n15603) );
  AOI31X1 U15438 ( .A0(n15605), .A1(n15606), .A2(n15607), .B0(n15414), .Y(
        n15604) );
  AOI21X1 U15439 ( .A0(n5403), .A1(n16863), .B0(n16864), .Y(n16862) );
  INVX1 U15440 ( .A(n16672), .Y(n5403) );
  NAND4BXL U15441 ( .AN(n16874), .B(n16726), .C(n16875), .D(n16876), .Y(n16863) );
  AOI31X1 U15442 ( .A0(n16865), .A1(n16866), .A2(n16867), .B0(n16674), .Y(
        n16864) );
  AOI21X1 U15443 ( .A0(n4849), .A1(n18753), .B0(n18754), .Y(n18752) );
  INVX1 U15444 ( .A(n18562), .Y(n4849) );
  NAND4BXL U15445 ( .AN(n18764), .B(n18616), .C(n18765), .D(n18766), .Y(n18753) );
  AOI31X1 U15446 ( .A0(n18755), .A1(n18756), .A2(n18757), .B0(n18564), .Y(
        n18754) );
  AOI21X1 U15447 ( .A0(n5868), .A1(n14973), .B0(n14974), .Y(n14972) );
  INVX1 U15448 ( .A(n14782), .Y(n5868) );
  NAND4BXL U15449 ( .AN(n14984), .B(n14836), .C(n14985), .D(n14986), .Y(n14973) );
  AOI31X1 U15450 ( .A0(n14975), .A1(n14976), .A2(n14977), .B0(n14784), .Y(
        n14974) );
  AOI21X1 U15451 ( .A0(n5480), .A1(n16548), .B0(n16549), .Y(n16547) );
  INVX1 U15452 ( .A(n16357), .Y(n5480) );
  NAND4BXL U15453 ( .AN(n16559), .B(n16411), .C(n16560), .D(n16561), .Y(n16548) );
  AOI31X1 U15454 ( .A0(n16550), .A1(n16551), .A2(n16552), .B0(n16359), .Y(
        n16549) );
  AOI21X1 U15455 ( .A0(n5050), .A1(n18123), .B0(n18124), .Y(n18122) );
  INVX1 U15456 ( .A(n17932), .Y(n5050) );
  NAND4BXL U15457 ( .AN(n18134), .B(n17986), .C(n18135), .D(n18136), .Y(n18123) );
  AOI31X1 U15458 ( .A0(n18125), .A1(n18126), .A2(n18127), .B0(n17934), .Y(
        n18124) );
  AOI21X1 U15459 ( .A0(n5944), .A1(n14658), .B0(n14659), .Y(n14657) );
  INVX1 U15460 ( .A(n14467), .Y(n5944) );
  NAND4BXL U15461 ( .AN(n14669), .B(n14521), .C(n14670), .D(n14671), .Y(n14658) );
  AOI31X1 U15462 ( .A0(n14660), .A1(n14661), .A2(n14662), .B0(n14469), .Y(
        n14659) );
  AOI21X1 U15463 ( .A0(n5556), .A1(n16233), .B0(n16234), .Y(n16232) );
  INVX1 U15464 ( .A(n16042), .Y(n5556) );
  NAND4BXL U15465 ( .AN(n16244), .B(n16096), .C(n16245), .D(n16246), .Y(n16233) );
  AOI31X1 U15466 ( .A0(n16235), .A1(n16236), .A2(n16237), .B0(n16044), .Y(
        n16234) );
  AOI21X1 U15467 ( .A0(n5158), .A1(n17808), .B0(n17809), .Y(n17807) );
  INVX1 U15468 ( .A(n17617), .Y(n5158) );
  NAND4BXL U15469 ( .AN(n17819), .B(n17671), .C(n17820), .D(n17821), .Y(n17808) );
  AOI31X1 U15470 ( .A0(n17810), .A1(n17811), .A2(n17812), .B0(n17619), .Y(
        n17809) );
  AOI21X1 U15471 ( .A0(n6020), .A1(n14343), .B0(n14344), .Y(n14342) );
  INVX1 U15472 ( .A(n14152), .Y(n6020) );
  NAND4BXL U15473 ( .AN(n14354), .B(n14206), .C(n14355), .D(n14356), .Y(n14343) );
  AOI31X1 U15474 ( .A0(n14345), .A1(n14346), .A2(n14347), .B0(n14154), .Y(
        n14344) );
  AOI21X1 U15475 ( .A0(n5632), .A1(n15918), .B0(n15919), .Y(n15917) );
  INVX1 U15476 ( .A(n15727), .Y(n5632) );
  NAND4BXL U15477 ( .AN(n15929), .B(n15781), .C(n15930), .D(n15931), .Y(n15918) );
  AOI31X1 U15478 ( .A0(n15920), .A1(n15921), .A2(n15922), .B0(n15729), .Y(
        n15919) );
  AOI21X1 U15479 ( .A0(n5236), .A1(n17493), .B0(n17494), .Y(n17492) );
  INVX1 U15480 ( .A(n17302), .Y(n5236) );
  NAND4BXL U15481 ( .AN(n17504), .B(n17356), .C(n17505), .D(n17506), .Y(n17493) );
  AOI31X1 U15482 ( .A0(n17495), .A1(n17496), .A2(n17497), .B0(n17304), .Y(
        n17494) );
  INVX1 U15483 ( .A(n11849), .Y(n6948) );
  INVX1 U15484 ( .A(top_core_KE_sb1_n278), .Y(n6933) );
  INVX1 U15485 ( .A(n12480), .Y(n6658) );
  INVX1 U15486 ( .A(n13425), .Y(n6633) );
  INVX1 U15487 ( .A(n12165), .Y(n6642) );
  INVX1 U15488 ( .A(n13110), .Y(n6940) );
  INVX1 U15489 ( .A(n13740), .Y(n6650) );
  INVX1 U15490 ( .A(n12795), .Y(n6925) );
  CLKINVX3 U15491 ( .A(n3987), .Y(n3983) );
  NAND2X1 U15492 ( .A(top_core_KE_n2703), .B(top_core_KE_n2701), .Y(
        top_core_KE_n895) );
  CLKINVX3 U15493 ( .A(n1679), .Y(n1673) );
  CLKINVX3 U15494 ( .A(n1736), .Y(n1731) );
  CLKINVX3 U15495 ( .A(n1707), .Y(n1702) );
  OAI21XL U15496 ( .A0(n667), .A1(n12337), .B0(n12403), .Y(n12402) );
  CLKINVX3 U15497 ( .A(n3975), .Y(n3963) );
  CLKINVX3 U15498 ( .A(n3973), .Y(n3964) );
  CLKINVX3 U15499 ( .A(n3974), .Y(n3972) );
  CLKINVX3 U15500 ( .A(n1669), .Y(n1666) );
  CLKINVX3 U15501 ( .A(n1698), .Y(n1695) );
  CLKINVX3 U15502 ( .A(n1727), .Y(n1724) );
  CLKINVX3 U15503 ( .A(n3985), .Y(n3976) );
  OAI2BB2X1 U15504 ( .B0(n1179), .B1(n13697), .A0N(n1277), .A1N(n13702), .Y(
        n13707) );
  OAI2BB2X1 U15505 ( .B0(n1174), .B1(n13382), .A0N(n1274), .A1N(n13387), .Y(
        n13392) );
  OAI2BB2X1 U15506 ( .B0(n1214), .B1(n12752), .A0N(n1268), .A1N(n12757), .Y(
        n12762) );
  OAI2BB2X1 U15507 ( .B0(n1220), .B1(n13067), .A0N(n1271), .A1N(n13072), .Y(
        n13077) );
  CLKINVX3 U15508 ( .A(n12437), .Y(n6626) );
  NAND4X1 U15509 ( .A(n13234), .B(n13283), .C(n13284), .D(n13285), .Y(n13273)
         );
  AOI22XL U15510 ( .A0(n13286), .A1(n52), .B0(n6544), .B1(n677), .Y(n13284) );
  NAND4X1 U15511 ( .A(n12604), .B(n12653), .C(n12654), .D(n12655), .Y(n12643)
         );
  AOI22XL U15512 ( .A0(n12656), .A1(n54), .B0(n6839), .B1(n678), .Y(n12654) );
  NAND4X1 U15513 ( .A(n12919), .B(n12968), .C(n12969), .D(n12970), .Y(n12958)
         );
  AOI22XL U15514 ( .A0(n12971), .A1(n56), .B0(n6885), .B1(n680), .Y(n12969) );
  NAND4X1 U15515 ( .A(n13549), .B(n13598), .C(n13599), .D(n13600), .Y(n13588)
         );
  AOI22XL U15516 ( .A0(n13601), .A1(n55), .B0(n6592), .B1(n679), .Y(n13599) );
  NAND4BXL U15517 ( .AN(n11817), .B(n11648), .C(n11799), .D(n11808), .Y(n11815) );
  NAND4BXL U15518 ( .AN(top_core_KE_sb1_n245), .B(top_core_KE_sb1_n73), .C(
        top_core_KE_sb1_n227), .D(top_core_KE_sb1_n236), .Y(
        top_core_KE_sb1_n243) );
  NAND4BXL U15519 ( .AN(n12448), .B(n12280), .C(n12430), .D(n12439), .Y(n12446) );
  NAND4BXL U15520 ( .AN(n12133), .B(n11964), .C(n12115), .D(n12124), .Y(n12131) );
  CLKINVX3 U15521 ( .A(top_core_KE_n900), .Y(n1632) );
  CLKINVX3 U15522 ( .A(top_core_io_inter_ok), .Y(n1582) );
  INVX1 U15523 ( .A(n11700), .Y(n6731) );
  INVX1 U15524 ( .A(top_core_KE_sb1_n125), .Y(n6794) );
  INVX1 U15525 ( .A(n12016), .Y(n6495) );
  INVX1 U15526 ( .A(n13277), .Y(n6462) );
  INVX1 U15527 ( .A(n12647), .Y(n6763) );
  INVX1 U15528 ( .A(n13592), .Y(n6419) );
  INVX1 U15529 ( .A(n12962), .Y(n6706) );
  INVX1 U15530 ( .A(n12331), .Y(n6439) );
  CLKINVX3 U15531 ( .A(top_core_io_inter_ok), .Y(n1583) );
  AOI21X1 U15532 ( .A0(n13721), .A1(n13722), .B0(n1635), .Y(n13719) );
  AOI211X1 U15533 ( .A0(n6592), .A1(n1652), .B0(n13633), .C0(n13723), .Y(
        n13722) );
  AOI21X1 U15534 ( .A0(n13608), .A1(n13598), .B0(n583), .Y(n13723) );
  CLKINVX3 U15535 ( .A(n1656), .Y(n1652) );
  AND2X2 U15536 ( .A(n1809), .B(n1807), .Y(n625) );
  AND2X2 U15537 ( .A(n1830), .B(n1828), .Y(n626) );
  AND2X2 U15538 ( .A(n1767), .B(n1764), .Y(n627) );
  AND2X2 U15539 ( .A(n1788), .B(n1786), .Y(n628) );
  AND2X2 U15540 ( .A(n1687), .B(n1684), .Y(n629) );
  AND2X2 U15541 ( .A(n1745), .B(n1742), .Y(n630) );
  AND2X2 U15542 ( .A(n1658), .B(n1655), .Y(n631) );
  AND2X2 U15543 ( .A(n1716), .B(n1713), .Y(n632) );
  CLKINVX3 U15544 ( .A(n3573), .Y(n3569) );
  INVX1 U15545 ( .A(top_core_EC_n948), .Y(n3573) );
  CLKINVX3 U15546 ( .A(n3573), .Y(n3572) );
  CLKINVX3 U15547 ( .A(n3708), .Y(n3696) );
  CLKINVX3 U15548 ( .A(n3706), .Y(n3697) );
  CLKINVX3 U15549 ( .A(n3705), .Y(n3698) );
  CLKINVX3 U15550 ( .A(n3708), .Y(n3699) );
  CLKINVX3 U15551 ( .A(n3707), .Y(n3700) );
  CLKINVX3 U15552 ( .A(n3706), .Y(n3701) );
  CLKINVX3 U15553 ( .A(n3706), .Y(n3702) );
  CLKINVX3 U15554 ( .A(n3705), .Y(n3703) );
  CLKINVX3 U15555 ( .A(n3708), .Y(n3689) );
  CLKINVX3 U15556 ( .A(n3708), .Y(n3690) );
  CLKINVX3 U15557 ( .A(n3707), .Y(n3691) );
  CLKINVX3 U15558 ( .A(n3707), .Y(n3692) );
  CLKINVX3 U15559 ( .A(n3705), .Y(n3693) );
  CLKINVX3 U15560 ( .A(n3708), .Y(n3694) );
  AOI21XL U15561 ( .A0(n11769), .A1(n11705), .B0(n673), .Y(n11944) );
  AOI21XL U15562 ( .A0(top_core_KE_sb1_n197), .A1(top_core_KE_sb1_n130), .B0(
        n674), .Y(top_core_KE_sb1_n374) );
  AOI21XL U15563 ( .A0(n12400), .A1(n12336), .B0(n675), .Y(n12575) );
  AOI21XL U15564 ( .A0(n13346), .A1(n1275), .B0(n677), .Y(n13520) );
  AOI21XL U15565 ( .A0(n12085), .A1(n12021), .B0(n676), .Y(n12260) );
  AOI21XL U15566 ( .A0(n12716), .A1(n12652), .B0(n678), .Y(n12890) );
  AOI21XL U15567 ( .A0(n13661), .A1(n13597), .B0(n679), .Y(n13835) );
  AOI21XL U15568 ( .A0(n13031), .A1(n12967), .B0(n680), .Y(n13205) );
  NAND4BXL U15569 ( .AN(n11833), .B(n11685), .C(n11834), .D(n11835), .Y(n11822) );
  AOI22X1 U15570 ( .A0(n11839), .A1(n625), .B0(n11654), .B1(n1203), .Y(n11834)
         );
  AOI21X1 U15571 ( .A0(n11837), .A1(n11838), .B0(n1795), .Y(n11836) );
  NAND4BXL U15572 ( .AN(top_core_KE_sb1_n262), .B(top_core_KE_sb1_n110), .C(
        top_core_KE_sb1_n263), .D(top_core_KE_sb1_n264), .Y(
        top_core_KE_sb1_n251) );
  AOI22X1 U15573 ( .A0(top_core_KE_sb1_n268), .A1(n626), .B0(
        top_core_KE_sb1_n79), .B1(n1194), .Y(top_core_KE_sb1_n263) );
  AOI21X1 U15574 ( .A0(top_core_KE_sb1_n266), .A1(top_core_KE_sb1_n267), .B0(
        n1816), .Y(top_core_KE_sb1_n265) );
  NAND4BXL U15575 ( .AN(n12464), .B(n12316), .C(n12465), .D(n12466), .Y(n12453) );
  AOI22X1 U15576 ( .A0(n12470), .A1(n627), .B0(n12286), .B1(n1163), .Y(n12465)
         );
  AOI21X1 U15577 ( .A0(n12468), .A1(n12469), .B0(n1752), .Y(n12467) );
  NAND4BXL U15578 ( .AN(n13409), .B(n13262), .C(n13410), .D(n13411), .Y(n13398) );
  AOI22X1 U15579 ( .A0(n13415), .A1(n629), .B0(n13231), .B1(n1149), .Y(n13410)
         );
  AOI21X1 U15580 ( .A0(n13413), .A1(n13414), .B0(n1672), .Y(n13412) );
  NAND4BXL U15581 ( .AN(n12149), .B(n12001), .C(n12150), .D(n12151), .Y(n12138) );
  AOI22X1 U15582 ( .A0(n12155), .A1(n628), .B0(n11970), .B1(n1154), .Y(n12150)
         );
  AOI21X1 U15583 ( .A0(n12153), .A1(n12154), .B0(n1774), .Y(n12152) );
  NAND4BXL U15584 ( .AN(n12779), .B(n12632), .C(n12780), .D(n12781), .Y(n12768) );
  AOI22X1 U15585 ( .A0(n12785), .A1(n630), .B0(n12601), .B1(n1189), .Y(n12780)
         );
  AOI21X1 U15586 ( .A0(n12783), .A1(n12784), .B0(n1729), .Y(n12782) );
  NAND4BXL U15587 ( .AN(n13724), .B(n13577), .C(n13725), .D(n13726), .Y(n13713) );
  AOI22X1 U15588 ( .A0(n13730), .A1(n631), .B0(n13546), .B1(n1158), .Y(n13725)
         );
  AOI21X1 U15589 ( .A0(n13728), .A1(n13729), .B0(n1635), .Y(n13727) );
  NAND4BXL U15590 ( .AN(n13094), .B(n12947), .C(n13095), .D(n13096), .Y(n13083) );
  AOI22X1 U15591 ( .A0(n13100), .A1(n632), .B0(n12916), .B1(n1198), .Y(n13095)
         );
  AOI21X1 U15592 ( .A0(n13098), .A1(n13099), .B0(n1700), .Y(n13097) );
  CLKINVX3 U15593 ( .A(n12483), .Y(n6611) );
  CLKINVX3 U15594 ( .A(n896), .Y(n3527) );
  CLKINVX3 U15595 ( .A(n896), .Y(n3528) );
  CLKINVX3 U15596 ( .A(n896), .Y(n3529) );
  CLKINVX3 U15597 ( .A(n896), .Y(n3530) );
  CLKINVX3 U15598 ( .A(n896), .Y(n3531) );
  CLKINVX3 U15599 ( .A(n896), .Y(n3532) );
  CLKINVX3 U15600 ( .A(n896), .Y(n3533) );
  CLKINVX3 U15601 ( .A(n1634), .Y(n1627) );
  CLKINVX3 U15602 ( .A(n1634), .Y(n1628) );
  CLKINVX3 U15603 ( .A(top_core_KE_n900), .Y(n1629) );
  CLKINVX3 U15604 ( .A(n1634), .Y(n1631) );
  CLKINVX3 U15605 ( .A(n1634), .Y(n1630) );
  CLKINVX3 U15606 ( .A(top_core_KE_n900), .Y(n1626) );
  CLKINVX3 U15607 ( .A(n3577), .Y(n3574) );
  CLKINVX3 U15608 ( .A(n3577), .Y(n3575) );
  CLKINVX3 U15609 ( .A(n1719), .Y(n1717) );
  CLKINVX3 U15610 ( .A(n1748), .Y(n1746) );
  CLKINVX3 U15611 ( .A(n1690), .Y(n1688) );
  AOI21X1 U15612 ( .A0(n13406), .A1(n13407), .B0(n1665), .Y(n13404) );
  AOI211X1 U15613 ( .A0(n6544), .A1(n1681), .B0(n13318), .C0(n13408), .Y(
        n13407) );
  AOI21X1 U15614 ( .A0(n13293), .A1(n13283), .B0(n580), .Y(n13408) );
  AOI21X1 U15615 ( .A0(n12776), .A1(n12777), .B0(n1723), .Y(n12774) );
  AOI211X1 U15616 ( .A0(n6839), .A1(n1739), .B0(n12688), .C0(n12778), .Y(
        n12777) );
  AOI21X1 U15617 ( .A0(n12663), .A1(n12653), .B0(n584), .Y(n12778) );
  AOI21X1 U15618 ( .A0(n13091), .A1(n13092), .B0(n1694), .Y(n13089) );
  AOI211X1 U15619 ( .A0(n6885), .A1(n1710), .B0(n13003), .C0(n13093), .Y(
        n13092) );
  AOI21X1 U15620 ( .A0(n12978), .A1(n12968), .B0(n582), .Y(n13093) );
  CLKINVX3 U15621 ( .A(n3581), .Y(n3578) );
  CLKINVX3 U15622 ( .A(n3581), .Y(n3579) );
  CLKINVX3 U15623 ( .A(n3581), .Y(n3580) );
  CLKINVX3 U15624 ( .A(n1634), .Y(n1633) );
  NAND4X1 U15625 ( .A(n11753), .B(n11773), .C(n11670), .D(n11757), .Y(n11770)
         );
  NAND4X1 U15626 ( .A(top_core_KE_sb1_n181), .B(top_core_KE_sb1_n201), .C(
        top_core_KE_sb1_n95), .D(top_core_KE_sb1_n185), .Y(
        top_core_KE_sb1_n198) );
  NAND4X1 U15627 ( .A(n12384), .B(n12404), .C(n12301), .D(n12388), .Y(n12401)
         );
  NAND4X1 U15628 ( .A(n13330), .B(n13350), .C(n13247), .D(n13334), .Y(n13347)
         );
  NAND4X1 U15629 ( .A(n12069), .B(n12089), .C(n11986), .D(n12073), .Y(n12086)
         );
  NAND4X1 U15630 ( .A(n12700), .B(n12720), .C(n12617), .D(n12704), .Y(n12717)
         );
  NAND4X1 U15631 ( .A(n13645), .B(n13665), .C(n13562), .D(n13649), .Y(n13662)
         );
  NAND4X1 U15632 ( .A(n13015), .B(n13035), .C(n12932), .D(n13019), .Y(n13032)
         );
  INVX1 U15633 ( .A(top_core_KE_n2695), .Y(n7011) );
  CLKINVX3 U15634 ( .A(n1762), .Y(n1761) );
  CLKINVX3 U15635 ( .A(n1700), .Y(n1696) );
  CLKINVX3 U15636 ( .A(n1729), .Y(n1725) );
  CLKINVX3 U15637 ( .A(n1671), .Y(n1667) );
  CLKINVX3 U15638 ( .A(n3707), .Y(n3695) );
  NAND4BXL U15639 ( .AN(n11642), .B(n11799), .C(n11908), .D(n11909), .Y(n11904) );
  AOI222X1 U15640 ( .A0(n673), .A1(n745), .B0(n6920), .B1(n1222), .C0(n1202), 
        .C1(n665), .Y(n11909) );
  AOI2BB2X1 U15641 ( .B0(n6919), .B1(n1809), .A0N(n11867), .A1N(n673), .Y(
        n11908) );
  NAND4BXL U15642 ( .AN(top_core_KE_sb1_n67), .B(top_core_KE_sb1_n227), .C(
        top_core_KE_sb1_n337), .D(top_core_KE_sb1_n338), .Y(
        top_core_KE_sb1_n333) );
  AOI222X1 U15643 ( .A0(n674), .A1(n746), .B0(n6874), .B1(n1216), .C0(n1193), 
        .C1(n666), .Y(top_core_KE_sb1_n338) );
  AOI2BB2X1 U15644 ( .B0(n6873), .B1(n1830), .A0N(top_core_KE_sb1_n296), .A1N(
        n674), .Y(top_core_KE_sb1_n337) );
  NAND4BXL U15645 ( .AN(n12274), .B(n12430), .C(n12539), .D(n12540), .Y(n12535) );
  AOI222X1 U15646 ( .A0(n675), .A1(n744), .B0(n6627), .B1(n1181), .C0(n1162), 
        .C1(n667), .Y(n12540) );
  AOI2BB2X1 U15647 ( .B0(n6626), .B1(n1767), .A0N(n12498), .A1N(n675), .Y(
        n12539) );
  NAND4BXL U15648 ( .AN(n11958), .B(n12115), .C(n12224), .D(n12225), .Y(n12220) );
  AOI222X1 U15649 ( .A0(n676), .A1(n747), .B0(n6580), .B1(n1176), .C0(n1153), 
        .C1(n668), .Y(n12225) );
  AOI2BB2X1 U15650 ( .B0(n6579), .B1(n1788), .A0N(n12183), .A1N(n676), .Y(
        n12224) );
  NAND4X1 U15651 ( .A(n13486), .B(n13487), .C(n13488), .D(n13489), .Y(n13479)
         );
  AOI2BB2X1 U15652 ( .B0(n1666), .B1(n13490), .A0N(n13252), .A1N(n692), .Y(
        n13488) );
  AOI2BB2X1 U15653 ( .B0(n6472), .B1(n13374), .A0N(n52), .A1N(n13239), .Y(
        n13486) );
  AOI22XL U15654 ( .A0(n13289), .A1(n13282), .B0(n13403), .B1(n686), .Y(n13487) );
  NAND4BXL U15655 ( .AN(n13241), .B(n13257), .C(n6558), .D(n13328), .Y(n13325)
         );
  AOI211X1 U15656 ( .A0(n6539), .A1(n602), .B0(n6635), .C0(n13329), .Y(n13328)
         );
  INVX1 U15657 ( .A(n13330), .Y(n6635) );
  AOI21XL U15658 ( .A0(n73), .A1(n13283), .B0(n1275), .Y(n13329) );
  NAND4BXL U15659 ( .AN(n12611), .B(n12627), .C(n6853), .D(n12698), .Y(n12695)
         );
  AOI211X1 U15660 ( .A0(n6834), .A1(n603), .B0(n6927), .C0(n12699), .Y(n12698)
         );
  INVX1 U15661 ( .A(n12700), .Y(n6927) );
  AOI21XL U15662 ( .A0(n74), .A1(n12653), .B0(n1269), .Y(n12699) );
  NAND4BXL U15663 ( .AN(n13556), .B(n13572), .C(n6606), .D(n13643), .Y(n13640)
         );
  AOI211X1 U15664 ( .A0(n6587), .A1(n609), .B0(n6652), .C0(n13644), .Y(n13643)
         );
  INVX1 U15665 ( .A(n13645), .Y(n6652) );
  AOI21XL U15666 ( .A0(n76), .A1(n13598), .B0(n1278), .Y(n13644) );
  NAND4BXL U15667 ( .AN(n12926), .B(n12942), .C(n6899), .D(n13013), .Y(n13010)
         );
  AOI211X1 U15668 ( .A0(n6880), .A1(n604), .B0(n6942), .C0(n13014), .Y(n13013)
         );
  INVX1 U15669 ( .A(n13015), .Y(n6942) );
  AOI21XL U15670 ( .A0(n75), .A1(n12968), .B0(n1272), .Y(n13014) );
  CLKINVX3 U15671 ( .A(n1662), .Y(n1659) );
  CLKINVX3 U15672 ( .A(n1807), .Y(n1803) );
  CLKINVX3 U15673 ( .A(n1828), .Y(n1824) );
  CLKINVX3 U15674 ( .A(n1786), .Y(n1782) );
  BUFX3 U15675 ( .A(n6589), .Y(n1157) );
  INVXL U15676 ( .A(n76), .Y(n6589) );
  BUFX3 U15677 ( .A(n723), .Y(n1134) );
  BUFX3 U15678 ( .A(n722), .Y(n995) );
  BUFX3 U15679 ( .A(n724), .Y(n939) );
  BUFX3 U15680 ( .A(n725), .Y(n1079) );
  BUFX3 U15681 ( .A(n726), .Y(n1065) );
  BUFX3 U15682 ( .A(n727), .Y(n1009) );
  BUFX3 U15683 ( .A(n728), .Y(n925) );
  BUFX3 U15684 ( .A(n729), .Y(n1093) );
  BUFX3 U15685 ( .A(n730), .Y(n1023) );
  BUFX3 U15686 ( .A(n731), .Y(n953) );
  BUFX3 U15687 ( .A(n732), .Y(n1107) );
  BUFX3 U15688 ( .A(n733), .Y(n1037) );
  BUFX3 U15689 ( .A(n734), .Y(n967) );
  BUFX3 U15690 ( .A(n735), .Y(n1121) );
  BUFX3 U15691 ( .A(n736), .Y(n1051) );
  BUFX3 U15692 ( .A(n737), .Y(n981) );
  CLKINVX3 U15693 ( .A(n765), .Y(n2145) );
  CLKINVX3 U15694 ( .A(n766), .Y(n3508) );
  CLKINVX3 U15695 ( .A(n764), .Y(n2236) );
  CLKINVX3 U15696 ( .A(n3568), .Y(n3565) );
  CLKINVX3 U15697 ( .A(n3568), .Y(n3566) );
  CLKINVX3 U15698 ( .A(n3568), .Y(n3567) );
  CLKINVX3 U15699 ( .A(n3548), .Y(n3544) );
  CLKINVX3 U15700 ( .A(n3548), .Y(n3545) );
  CLKINVX3 U15701 ( .A(n3548), .Y(n3546) );
  CLKINVX3 U15702 ( .A(n3548), .Y(n3547) );
  CLKINVX3 U15703 ( .A(n2252), .Y(n2248) );
  CLKINVX3 U15704 ( .A(n2252), .Y(n2250) );
  CLKINVX3 U15705 ( .A(n2252), .Y(n2245) );
  CLKINVX3 U15706 ( .A(n2253), .Y(n2251) );
  CLKINVX3 U15707 ( .A(n2252), .Y(n2249) );
  CLKINVX3 U15708 ( .A(n2252), .Y(n2246) );
  CLKINVX3 U15709 ( .A(n2253), .Y(n2247) );
  CLKINVX3 U15710 ( .A(n3525), .Y(n3516) );
  INVX1 U15711 ( .A(top_core_EC_n730), .Y(n3525) );
  BUFX3 U15712 ( .A(top_core_EC_mc_mix_in_4_24_), .Y(n1546) );
  OAI22X1 U15713 ( .A0(n2484), .A1(top_core_EC_ss_n206), .B0(n2369), .B1(n4832), .Y(top_core_EC_mc_mix_in_4_24_) );
  BUFX3 U15714 ( .A(top_core_EC_mc_mix_in_8[24]), .Y(n1547) );
  OAI22X1 U15715 ( .A0(n2482), .A1(top_core_EC_ss_n208), .B0(n2369), .B1(n4846), .Y(top_core_EC_mc_mix_in_8[24]) );
  XOR2X1 U15716 ( .A(top_core_EC_mc_mix_in_8[80]), .B(
        top_core_EC_mc_mix_in_4_80_), .Y(top_core_EC_mc_mix_in_8[81]) );
  XOR2X1 U15717 ( .A(top_core_EC_mc_mix_in_8[80]), .B(
        top_core_EC_mc_mix_in_4_82_), .Y(top_core_EC_mc_mix_in_8[83]) );
  XOR2X1 U15718 ( .A(top_core_EC_mc_mix_in_8[80]), .B(
        top_core_EC_mc_mix_in_4_83_), .Y(top_core_EC_mc_mix_in_8[84]) );
  XOR2X1 U15719 ( .A(top_core_EC_mc_mix_in_8[64]), .B(
        top_core_EC_mc_mix_in_4_64_), .Y(top_core_EC_mc_mix_in_8[65]) );
  XOR2X1 U15720 ( .A(top_core_EC_mc_mix_in_8[64]), .B(
        top_core_EC_mc_mix_in_4_66_), .Y(top_core_EC_mc_mix_in_8[67]) );
  XOR2X1 U15721 ( .A(top_core_EC_mc_mix_in_8[64]), .B(
        top_core_EC_mc_mix_in_4_67_), .Y(top_core_EC_mc_mix_in_8[68]) );
  XOR2X1 U15722 ( .A(top_core_EC_mc_mix_in_8[112]), .B(
        top_core_EC_mc_mix_in_4_115_), .Y(top_core_EC_mc_mix_in_8[116]) );
  XOR2X1 U15723 ( .A(top_core_EC_mc_mix_in_8[96]), .B(
        top_core_EC_mc_mix_in_4_99_), .Y(top_core_EC_mc_mix_in_8[100]) );
  BUFX3 U15724 ( .A(n6605), .Y(n1161) );
  INVXL U15725 ( .A(n183), .Y(n6605) );
  CLKINVX3 U15726 ( .A(n2188), .Y(n2183) );
  CLKINVX3 U15727 ( .A(n2189), .Y(n2184) );
  CLKINVX3 U15728 ( .A(n2189), .Y(n2185) );
  CLKINVX3 U15729 ( .A(n2188), .Y(n2186) );
  CLKINVX3 U15730 ( .A(n2189), .Y(n2187) );
  CLKINVX3 U15731 ( .A(n3577), .Y(n3576) );
  BUFX3 U15732 ( .A(top_core_EC_mc_mix_in_4_40_), .Y(n1543) );
  OAI22X1 U15733 ( .A0(n2433), .A1(top_core_EC_ss_n189), .B0(n2371), .B1(n5393), .Y(top_core_EC_mc_mix_in_4_40_) );
  BUFX3 U15734 ( .A(top_core_EC_mc_mix_in_8[40]), .Y(n1544) );
  OAI22X1 U15735 ( .A0(n2433), .A1(top_core_EC_ss_n190), .B0(n2370), .B1(n5400), .Y(top_core_EC_mc_mix_in_8[40]) );
  BUFX3 U15736 ( .A(top_core_EC_mc_mix_in_8[8]), .Y(n1550) );
  OAI22X1 U15737 ( .A0(n2410), .A1(top_core_EC_ss_n225), .B0(n2368), .B1(n5041), .Y(top_core_EC_mc_mix_in_8[8]) );
  BUFX3 U15738 ( .A(top_core_EC_mc_mix_in_4_8_), .Y(n1549) );
  OAI22X1 U15739 ( .A0(n2409), .A1(top_core_EC_ss_n224), .B0(n2368), .B1(n5040), .Y(top_core_EC_mc_mix_in_4_8_) );
  BUFX3 U15740 ( .A(top_core_EC_mc_mix_in_2_24_), .Y(n1545) );
  OAI22X1 U15741 ( .A0(n2401), .A1(top_core_EC_ss_n205), .B0(n2369), .B1(n4845), .Y(top_core_EC_mc_mix_in_2_24_) );
  CLKINVX3 U15742 ( .A(n2169), .Y(n2168) );
  CLKINVX3 U15743 ( .A(n2170), .Y(n2167) );
  CLKINVX3 U15744 ( .A(n2169), .Y(n2166) );
  CLKINVX3 U15745 ( .A(n2170), .Y(n2165) );
  CLKINVX3 U15746 ( .A(n2169), .Y(n2164) );
  CLKINVX3 U15747 ( .A(n2169), .Y(n2163) );
  CLKINVX3 U15748 ( .A(n2169), .Y(n2162) );
  CLKINVX3 U15749 ( .A(n2170), .Y(n2161) );
  INVX1 U15750 ( .A(n13949), .Y(n6172) );
  INVX1 U15751 ( .A(n17099), .Y(n5390) );
  INVX1 U15752 ( .A(n15209), .Y(n5862) );
  INVX1 U15753 ( .A(n18359), .Y(n5036) );
  INVX1 U15754 ( .A(n15524), .Y(n5778) );
  INVX1 U15755 ( .A(n16784), .Y(n5474) );
  INVX1 U15756 ( .A(n14894), .Y(n5938) );
  INVX1 U15757 ( .A(n16469), .Y(n5550) );
  INVX1 U15758 ( .A(n18044), .Y(n5120) );
  INVX1 U15759 ( .A(n14579), .Y(n6014) );
  INVX1 U15760 ( .A(n16154), .Y(n5626) );
  INVX1 U15761 ( .A(n17729), .Y(n5228) );
  INVX1 U15762 ( .A(n14264), .Y(n6090) );
  INVX1 U15763 ( .A(n15839), .Y(n5702) );
  INVX1 U15764 ( .A(n17414), .Y(n5306) );
  INVX1 U15765 ( .A(n18674), .Y(n4920) );
  XOR2X1 U15766 ( .A(n1556), .B(top_core_EC_mc_mix_in_4_106_), .Y(
        top_core_EC_mc_mix_in_8[107]) );
  CLKINVX3 U15767 ( .A(n1770), .Y(n1768) );
  XOR2X1 U15768 ( .A(n1553), .B(top_core_EC_mc_mix_in_4_122_), .Y(
        top_core_EC_mc_mix_in_8[123]) );
  CLKINVX3 U15769 ( .A(n2263), .Y(n2258) );
  CLKINVX3 U15770 ( .A(n2262), .Y(n2260) );
  CLKINVX3 U15771 ( .A(n2263), .Y(n2255) );
  CLKINVX3 U15772 ( .A(n2263), .Y(n2259) );
  CLKINVX3 U15773 ( .A(n2262), .Y(n2256) );
  CLKINVX3 U15774 ( .A(n2263), .Y(n2257) );
  XOR2X1 U15775 ( .A(n1553), .B(n1552), .Y(top_core_EC_mc_mix_in_8[121]) );
  XOR2X1 U15776 ( .A(n1556), .B(n1555), .Y(top_core_EC_mc_mix_in_8[105]) );
  CLKINVX3 U15777 ( .A(n2311), .Y(n2307) );
  CLKINVX3 U15778 ( .A(n2311), .Y(n2308) );
  CLKINVX3 U15779 ( .A(n2311), .Y(n2309) );
  CLKINVX3 U15780 ( .A(n2273), .Y(n2264) );
  INVX1 U15781 ( .A(top_core_KE_n1876), .Y(n2273) );
  CLKINVX3 U15782 ( .A(n2311), .Y(n2310) );
  CLKINVX3 U15783 ( .A(n2188), .Y(n2181) );
  CLKINVX3 U15784 ( .A(n2189), .Y(n2182) );
  CLKINVX3 U15785 ( .A(n2282), .Y(n2279) );
  CLKINVX3 U15786 ( .A(n2282), .Y(n2275) );
  CLKINVX3 U15787 ( .A(n2282), .Y(n2281) );
  CLKINVX3 U15788 ( .A(n2282), .Y(n2280) );
  CLKINVX3 U15789 ( .A(n2283), .Y(n2277) );
  CLKINVX3 U15790 ( .A(n2283), .Y(n2276) );
  CLKINVX3 U15791 ( .A(n2282), .Y(n2278) );
  OAI2BB1X1 U15792 ( .A0N(n17140), .A1N(n17141), .B0(n992), .Y(n17139) );
  AOI22X1 U15793 ( .A0(n17051), .A1(n17146), .B0(n2846), .B1(n17147), .Y(
        n17140) );
  AOI22X1 U15794 ( .A0(n481), .A1(n17068), .B0(n5321), .B1(n17142), .Y(n17141)
         );
  OAI221XL U15795 ( .A0(n1003), .A1(n17072), .B0(n386), .B1(n106), .C0(n17156), 
        .Y(n17146) );
  OAI2BB1X1 U15796 ( .A0N(n13990), .A1N(n13991), .B0(n1132), .Y(n13989) );
  AOI22X1 U15797 ( .A0(n13901), .A1(n13996), .B0(n3447), .B1(n13997), .Y(
        n13990) );
  AOI22X1 U15798 ( .A0(n482), .A1(n13918), .B0(n6105), .B1(n13992), .Y(n13991)
         );
  OAI221XL U15799 ( .A0(n1142), .A1(n13922), .B0(n385), .B1(n107), .C0(n14006), 
        .Y(n13996) );
  OAI2BB1X1 U15800 ( .A0N(n18400), .A1N(n18401), .B0(n936), .Y(n18399) );
  AOI22X1 U15801 ( .A0(n18311), .A1(n18406), .B0(n2604), .B1(n18407), .Y(
        n18400) );
  AOI22X1 U15802 ( .A0(n483), .A1(n18328), .B0(n4967), .B1(n18402), .Y(n18401)
         );
  OAI221XL U15803 ( .A0(n947), .A1(n18332), .B0(n387), .B1(n108), .C0(n18416), 
        .Y(n18406) );
  OAI2BB1X1 U15804 ( .A0N(n15250), .A1N(n15251), .B0(n1076), .Y(n15249) );
  AOI22X1 U15805 ( .A0(n15161), .A1(n15256), .B0(n3206), .B1(n15257), .Y(
        n15250) );
  AOI22X1 U15806 ( .A0(n484), .A1(n15178), .B0(n5793), .B1(n15252), .Y(n15251)
         );
  OAI221XL U15807 ( .A0(n1087), .A1(n15182), .B0(n388), .B1(n109), .C0(n15266), 
        .Y(n15256) );
  OAI2BB1X1 U15808 ( .A0N(n15565), .A1N(n15566), .B0(n1062), .Y(n15564) );
  AOI22X1 U15809 ( .A0(n15476), .A1(n15571), .B0(n3145), .B1(n15572), .Y(
        n15565) );
  AOI22X1 U15810 ( .A0(n490), .A1(n15493), .B0(n5709), .B1(n15567), .Y(n15566)
         );
  OAI221XL U15811 ( .A0(n1073), .A1(n15497), .B0(n389), .B1(n110), .C0(n15581), 
        .Y(n15571) );
  OAI2BB1X1 U15812 ( .A0N(n18715), .A1N(n18716), .B0(n922), .Y(n18714) );
  AOI22X1 U15813 ( .A0(n18626), .A1(n18721), .B0(n2543), .B1(n18722), .Y(
        n18715) );
  AOI22X1 U15814 ( .A0(n492), .A1(n18643), .B0(n4851), .B1(n18717), .Y(n18716)
         );
  OAI221XL U15815 ( .A0(n933), .A1(n18647), .B0(n390), .B1(n111), .C0(n18731), 
        .Y(n18721) );
  OAI2BB1X1 U15816 ( .A0N(n16825), .A1N(n16826), .B0(n1006), .Y(n16824) );
  AOI22X1 U15817 ( .A0(n16736), .A1(n16831), .B0(n2907), .B1(n16832), .Y(
        n16825) );
  AOI22X1 U15818 ( .A0(n494), .A1(n16753), .B0(n5405), .B1(n16827), .Y(n16826)
         );
  OAI221XL U15819 ( .A0(n1017), .A1(n16757), .B0(n391), .B1(n112), .C0(n16841), 
        .Y(n16831) );
  OAI2BB1X1 U15820 ( .A0N(n14935), .A1N(n14936), .B0(n1090), .Y(n14934) );
  AOI22X1 U15821 ( .A0(n14846), .A1(n14941), .B0(n3267), .B1(n14942), .Y(
        n14935) );
  AOI22X1 U15822 ( .A0(n496), .A1(n14863), .B0(n5869), .B1(n14937), .Y(n14936)
         );
  OAI221XL U15823 ( .A0(n1101), .A1(n14867), .B0(n392), .B1(n113), .C0(n14951), 
        .Y(n14941) );
  OAI2BB1X1 U15824 ( .A0N(n16510), .A1N(n16511), .B0(n1020), .Y(n16509) );
  AOI22X1 U15825 ( .A0(n16421), .A1(n16516), .B0(n2968), .B1(n16517), .Y(
        n16510) );
  AOI22X1 U15826 ( .A0(n489), .A1(n16438), .B0(n5481), .B1(n16512), .Y(n16511)
         );
  OAI221XL U15827 ( .A0(n1031), .A1(n16442), .B0(n393), .B1(n114), .C0(n16526), 
        .Y(n16516) );
  OAI2BB1X1 U15828 ( .A0N(n18085), .A1N(n18086), .B0(n950), .Y(n18084) );
  AOI22X1 U15829 ( .A0(n17996), .A1(n18091), .B0(n2665), .B1(n18092), .Y(
        n18085) );
  AOI22X1 U15830 ( .A0(n485), .A1(n18013), .B0(n5051), .B1(n18087), .Y(n18086)
         );
  OAI221XL U15831 ( .A0(n961), .A1(n18017), .B0(n394), .B1(n115), .C0(n18101), 
        .Y(n18091) );
  OAI2BB1X1 U15832 ( .A0N(n14620), .A1N(n14621), .B0(n1104), .Y(n14619) );
  AOI22X1 U15833 ( .A0(n14531), .A1(n14626), .B0(n3328), .B1(n14627), .Y(
        n14620) );
  AOI22X1 U15834 ( .A0(n491), .A1(n14548), .B0(n5945), .B1(n14622), .Y(n14621)
         );
  OAI221XL U15835 ( .A0(n1115), .A1(n14552), .B0(n395), .B1(n116), .C0(n14636), 
        .Y(n14626) );
  OAI2BB1X1 U15836 ( .A0N(n16195), .A1N(n16196), .B0(n1034), .Y(n16194) );
  AOI22X1 U15837 ( .A0(n16106), .A1(n16201), .B0(n3026), .B1(n16202), .Y(
        n16195) );
  AOI22X1 U15838 ( .A0(n486), .A1(n16123), .B0(n5557), .B1(n16197), .Y(n16196)
         );
  OAI221XL U15839 ( .A0(n1045), .A1(n16127), .B0(n396), .B1(n117), .C0(n16211), 
        .Y(n16201) );
  OAI2BB1X1 U15840 ( .A0N(n17770), .A1N(n17771), .B0(n964), .Y(n17769) );
  AOI22X1 U15841 ( .A0(n17681), .A1(n17776), .B0(n2725), .B1(n17777), .Y(
        n17770) );
  AOI22X1 U15842 ( .A0(n493), .A1(n17698), .B0(n5159), .B1(n17772), .Y(n17771)
         );
  OAI221XL U15843 ( .A0(n975), .A1(n17702), .B0(n397), .B1(n118), .C0(n17786), 
        .Y(n17776) );
  OAI2BB1X1 U15844 ( .A0N(n14305), .A1N(n14306), .B0(n1118), .Y(n14304) );
  AOI22X1 U15845 ( .A0(n14216), .A1(n14311), .B0(n3386), .B1(n14312), .Y(
        n14305) );
  AOI22X1 U15846 ( .A0(n487), .A1(n14233), .B0(n6021), .B1(n14307), .Y(n14306)
         );
  OAI221XL U15847 ( .A0(n1129), .A1(n14237), .B0(n398), .B1(n119), .C0(n14321), 
        .Y(n14311) );
  OAI2BB1X1 U15848 ( .A0N(n15880), .A1N(n15881), .B0(n1048), .Y(n15879) );
  AOI22X1 U15849 ( .A0(n15791), .A1(n15886), .B0(n3087), .B1(n15887), .Y(
        n15880) );
  AOI22X1 U15850 ( .A0(n495), .A1(n15808), .B0(n5633), .B1(n15882), .Y(n15881)
         );
  OAI221XL U15851 ( .A0(n1059), .A1(n15812), .B0(n399), .B1(n120), .C0(n15896), 
        .Y(n15886) );
  OAI2BB1X1 U15852 ( .A0N(n17455), .A1N(n17456), .B0(n978), .Y(n17454) );
  AOI22X1 U15853 ( .A0(n17366), .A1(n17461), .B0(n2786), .B1(n17462), .Y(
        n17455) );
  AOI22X1 U15854 ( .A0(n488), .A1(n17383), .B0(n5237), .B1(n17457), .Y(n17456)
         );
  OAI221XL U15855 ( .A0(n989), .A1(n17387), .B0(n400), .B1(n121), .C0(n17471), 
        .Y(n17461) );
  XOR2X1 U15856 ( .A(top_core_EC_mc_mix_in_8[96]), .B(
        top_core_EC_mc_mix_in_4_96_), .Y(top_core_EC_mc_mix_in_8[97]) );
  XOR2X1 U15857 ( .A(top_core_EC_mc_mix_in_8[96]), .B(
        top_core_EC_mc_mix_in_4_98_), .Y(top_core_EC_mc_mix_in_8[99]) );
  BUFX3 U15858 ( .A(top_core_EC_mc_mix_in_2_40_), .Y(n1542) );
  OAI22X1 U15859 ( .A0(n2433), .A1(top_core_EC_ss_n188), .B0(n2371), .B1(n5399), .Y(top_core_EC_mc_mix_in_2_40_) );
  XNOR2X1 U15860 ( .A(top_core_EC_mc_mix_in_8[95]), .B(top_core_EC_mc_n149), 
        .Y(top_core_EC_mc_n268) );
  XNOR2X1 U15861 ( .A(top_core_EC_mc_mix_in_8[127]), .B(top_core_EC_mc_n808), 
        .Y(top_core_EC_mc_n916) );
  XNOR2X1 U15862 ( .A(top_core_EC_mc_mix_in_8[79]), .B(top_core_EC_mc_n141), 
        .Y(top_core_EC_mc_n205) );
  XNOR2X1 U15863 ( .A(top_core_EC_mc_mix_in_8[111]), .B(top_core_EC_mc_n800), 
        .Y(top_core_EC_mc_n854) );
  BUFX3 U15864 ( .A(top_core_EC_mc_mix_in_2_8_), .Y(n1548) );
  OAI22X1 U15865 ( .A0(n2408), .A1(top_core_EC_ss_n223), .B0(n2368), .B1(n5039), .Y(top_core_EC_mc_mix_in_2_8_) );
  XNOR2X1 U15866 ( .A(top_core_EC_mc_mix_in_2_90_), .B(top_core_EC_mc_n173), 
        .Y(top_core_EC_mc_n292) );
  XNOR2X1 U15867 ( .A(top_core_EC_mc_mix_in_2_122_), .B(top_core_EC_mc_n35), 
        .Y(top_core_EC_mc_n31) );
  INVX1 U15868 ( .A(top_core_EC_mix_out_61_), .Y(n4936) );
  OAI22X1 U15869 ( .A0(top_core_EC_mc_n322), .A1(n2457), .B0(n2381), .B1(
        top_core_EC_mc_n323), .Y(top_core_EC_mix_out_61_) );
  XOR2X1 U15870 ( .A(top_core_EC_mc_n324), .B(top_core_EC_mc_n325), .Y(
        top_core_EC_mc_n323) );
  XNOR2X1 U15871 ( .A(top_core_EC_mc_mix_in_8[63]), .B(top_core_EC_mc_n326), 
        .Y(top_core_EC_mc_n322) );
  INVX1 U15872 ( .A(top_core_EC_mix_out_62_), .Y(n4933) );
  OAI22X1 U15873 ( .A0(top_core_EC_mc_n314), .A1(n2458), .B0(n2382), .B1(
        top_core_EC_mc_n315), .Y(top_core_EC_mix_out_62_) );
  XOR2X1 U15874 ( .A(top_core_EC_mc_n316), .B(top_core_EC_mc_n317), .Y(
        top_core_EC_mc_n315) );
  XNOR2X1 U15875 ( .A(n1541), .B(top_core_EC_mc_n318), .Y(top_core_EC_mc_n314)
         );
  INVX1 U15876 ( .A(top_core_EC_mix_out_63_), .Y(n4925) );
  OAI22X1 U15877 ( .A0(top_core_EC_mc_n306), .A1(n2459), .B0(n2382), .B1(
        top_core_EC_mc_n307), .Y(top_core_EC_mix_out_63_) );
  XOR2X1 U15878 ( .A(top_core_EC_mc_n308), .B(top_core_EC_mc_n309), .Y(
        top_core_EC_mc_n307) );
  XNOR2X1 U15879 ( .A(n1540), .B(top_core_EC_mc_n310), .Y(top_core_EC_mc_n306)
         );
  INVX1 U15880 ( .A(top_core_EC_mix_out_64_), .Y(n4806) );
  OAI22X1 U15881 ( .A0(top_core_EC_mc_n298), .A1(n2452), .B0(n2382), .B1(
        top_core_EC_mc_n299), .Y(top_core_EC_mix_out_64_) );
  XOR2X1 U15882 ( .A(top_core_EC_mc_n300), .B(top_core_EC_mc_n301), .Y(
        top_core_EC_mc_n299) );
  XNOR2X1 U15883 ( .A(top_core_EC_mix_in[88]), .B(top_core_EC_mc_n302), .Y(
        top_core_EC_mc_n298) );
  INVX1 U15884 ( .A(top_core_EC_mix_out_65_), .Y(n4804) );
  OAI22X1 U15885 ( .A0(top_core_EC_mc_n290), .A1(n2453), .B0(n2382), .B1(
        top_core_EC_mc_n291), .Y(top_core_EC_mix_out_65_) );
  XOR2X1 U15886 ( .A(top_core_EC_mc_n292), .B(top_core_EC_mc_n293), .Y(
        top_core_EC_mc_n291) );
  XNOR2X1 U15887 ( .A(top_core_EC_mc_mix_in_2_90_), .B(top_core_EC_mc_n294), 
        .Y(top_core_EC_mc_n290) );
  INVX1 U15888 ( .A(top_core_EC_mix_out_66_), .Y(n4798) );
  OAI22X1 U15889 ( .A0(top_core_EC_mc_n282), .A1(n2455), .B0(n2382), .B1(
        top_core_EC_mc_n283), .Y(top_core_EC_mix_out_66_) );
  XOR2X1 U15890 ( .A(top_core_EC_mc_n284), .B(top_core_EC_mc_n285), .Y(
        top_core_EC_mc_n283) );
  XNOR2X1 U15891 ( .A(top_core_EC_mix_in[90]), .B(top_core_EC_mc_n286), .Y(
        top_core_EC_mc_n282) );
  INVX1 U15892 ( .A(top_core_EC_mix_out_67_), .Y(n4793) );
  OAI22X1 U15893 ( .A0(top_core_EC_mc_n274), .A1(n2429), .B0(n2382), .B1(
        top_core_EC_mc_n275), .Y(top_core_EC_mix_out_67_) );
  XOR2X1 U15894 ( .A(top_core_EC_mc_n276), .B(top_core_EC_mc_n277), .Y(
        top_core_EC_mc_n275) );
  XNOR2X1 U15895 ( .A(top_core_EC_mix_in[91]), .B(top_core_EC_mc_n278), .Y(
        top_core_EC_mc_n274) );
  INVX1 U15896 ( .A(top_core_EC_mix_out_68_), .Y(n4803) );
  OAI22X1 U15897 ( .A0(top_core_EC_mc_n266), .A1(n2431), .B0(n2382), .B1(
        top_core_EC_mc_n267), .Y(top_core_EC_mix_out_68_) );
  XOR2X1 U15898 ( .A(top_core_EC_mc_n268), .B(top_core_EC_mc_n269), .Y(
        top_core_EC_mc_n267) );
  XNOR2X1 U15899 ( .A(top_core_EC_mc_mix_in_8[95]), .B(top_core_EC_mc_n270), 
        .Y(top_core_EC_mc_n266) );
  INVX1 U15900 ( .A(top_core_EC_mix_out_69_), .Y(n4787) );
  OAI22X1 U15901 ( .A0(top_core_EC_mc_n258), .A1(n2450), .B0(n2382), .B1(
        top_core_EC_mc_n259), .Y(top_core_EC_mix_out_69_) );
  XOR2X1 U15902 ( .A(top_core_EC_mc_n260), .B(top_core_EC_mc_n261), .Y(
        top_core_EC_mc_n259) );
  XNOR2X1 U15903 ( .A(n1535), .B(top_core_EC_mc_n262), .Y(top_core_EC_mc_n258)
         );
  INVX1 U15904 ( .A(top_core_EC_mix_out_70_), .Y(n4782) );
  OAI22X1 U15905 ( .A0(top_core_EC_mc_n241), .A1(n2530), .B0(n2382), .B1(
        top_core_EC_mc_n242), .Y(top_core_EC_mix_out_70_) );
  XOR2X1 U15906 ( .A(top_core_EC_mc_n243), .B(top_core_EC_mc_n244), .Y(
        top_core_EC_mc_n242) );
  XNOR2X1 U15907 ( .A(n1534), .B(top_core_EC_mc_n245), .Y(top_core_EC_mc_n241)
         );
  INVX1 U15908 ( .A(top_core_EC_mix_out_71_), .Y(n4775) );
  OAI22X1 U15909 ( .A0(top_core_EC_mc_n233), .A1(n2529), .B0(n2382), .B1(
        top_core_EC_mc_n234), .Y(top_core_EC_mix_out_71_) );
  XOR2X1 U15910 ( .A(top_core_EC_mc_n235), .B(top_core_EC_mc_n236), .Y(
        top_core_EC_mc_n234) );
  XNOR2X1 U15911 ( .A(n1533), .B(top_core_EC_mc_n237), .Y(top_core_EC_mc_n233)
         );
  INVX1 U15912 ( .A(top_core_EC_mix_out_72_), .Y(n4805) );
  OAI22X1 U15913 ( .A0(top_core_EC_mc_n228), .A1(n2525), .B0(n2382), .B1(
        top_core_EC_mc_n229), .Y(top_core_EC_mix_out_72_) );
  XOR2X1 U15914 ( .A(top_core_EC_mc_n230), .B(top_core_EC_mc_n231), .Y(
        top_core_EC_mc_n229) );
  XNOR2X1 U15915 ( .A(n1536), .B(top_core_EC_mc_n232), .Y(top_core_EC_mc_n228)
         );
  INVX1 U15916 ( .A(top_core_EC_mix_out_74_), .Y(n4795) );
  OAI22X1 U15917 ( .A0(top_core_EC_mc_n218), .A1(n2542), .B0(n2382), .B1(
        top_core_EC_mc_n219), .Y(top_core_EC_mix_out_74_) );
  XOR2X1 U15918 ( .A(top_core_EC_mc_n220), .B(top_core_EC_mc_n221), .Y(
        top_core_EC_mc_n219) );
  XNOR2X1 U15919 ( .A(top_core_EC_mc_mix_in_2_74_), .B(top_core_EC_mc_n222), 
        .Y(top_core_EC_mc_n218) );
  INVX1 U15920 ( .A(top_core_EC_mix_out_77_), .Y(n4780) );
  OAI22X1 U15921 ( .A0(top_core_EC_mc_n203), .A1(n2439), .B0(n2383), .B1(
        top_core_EC_mc_n204), .Y(top_core_EC_mix_out_77_) );
  XOR2X1 U15922 ( .A(top_core_EC_mc_n205), .B(top_core_EC_mc_n206), .Y(
        top_core_EC_mc_n204) );
  XNOR2X1 U15923 ( .A(top_core_EC_mc_mix_in_8[79]), .B(top_core_EC_mc_n207), 
        .Y(top_core_EC_mc_n203) );
  INVX1 U15924 ( .A(top_core_EC_mix_out_78_), .Y(n4783) );
  OAI22X1 U15925 ( .A0(top_core_EC_mc_n198), .A1(n2426), .B0(n2383), .B1(
        top_core_EC_mc_n199), .Y(top_core_EC_mix_out_78_) );
  XOR2X1 U15926 ( .A(top_core_EC_mc_n200), .B(top_core_EC_mc_n201), .Y(
        top_core_EC_mc_n199) );
  XNOR2X1 U15927 ( .A(n1538), .B(top_core_EC_mc_n202), .Y(top_core_EC_mc_n198)
         );
  INVX1 U15928 ( .A(top_core_EC_mix_out_79_), .Y(n4776) );
  OAI22X1 U15929 ( .A0(top_core_EC_mc_n193), .A1(n2433), .B0(n2383), .B1(
        top_core_EC_mc_n194), .Y(top_core_EC_mix_out_79_) );
  XOR2X1 U15930 ( .A(top_core_EC_mc_n195), .B(top_core_EC_mc_n196), .Y(
        top_core_EC_mc_n194) );
  XNOR2X1 U15931 ( .A(n1537), .B(top_core_EC_mc_n197), .Y(top_core_EC_mc_n193)
         );
  INVX1 U15932 ( .A(top_core_EC_mix_out_80_), .Y(n4800) );
  OAI22X1 U15933 ( .A0(top_core_EC_mc_n176), .A1(n2451), .B0(n2383), .B1(
        top_core_EC_mc_n177), .Y(top_core_EC_mix_out_80_) );
  XOR2X1 U15934 ( .A(top_core_EC_mc_n114), .B(top_core_EC_mc_n178), .Y(
        top_core_EC_mc_n177) );
  XNOR2X1 U15935 ( .A(n1533), .B(top_core_EC_mc_n179), .Y(top_core_EC_mc_n176)
         );
  INVX1 U15936 ( .A(top_core_EC_mix_out_82_), .Y(n4799) );
  OAI22X1 U15937 ( .A0(top_core_EC_mc_n160), .A1(n2407), .B0(n2383), .B1(
        top_core_EC_mc_n161), .Y(top_core_EC_mix_out_82_) );
  XOR2X1 U15938 ( .A(top_core_EC_mc_n89), .B(top_core_EC_mc_n162), .Y(
        top_core_EC_mc_n161) );
  XNOR2X1 U15939 ( .A(top_core_EC_mc_mix_in_2_90_), .B(top_core_EC_mc_n163), 
        .Y(top_core_EC_mc_n160) );
  INVX1 U15940 ( .A(top_core_EC_mix_out_85_), .Y(n4788) );
  OAI22X1 U15941 ( .A0(top_core_EC_mc_n136), .A1(n2524), .B0(n2383), .B1(
        top_core_EC_mc_n137), .Y(top_core_EC_mix_out_85_) );
  XOR2X1 U15942 ( .A(top_core_EC_mc_n65), .B(top_core_EC_mc_n138), .Y(
        top_core_EC_mc_n137) );
  XNOR2X1 U15943 ( .A(top_core_EC_mc_mix_in_8[95]), .B(top_core_EC_mc_n139), 
        .Y(top_core_EC_mc_n136) );
  INVX1 U15944 ( .A(top_core_EC_mix_out_86_), .Y(n4784) );
  OAI22X1 U15945 ( .A0(top_core_EC_mc_n128), .A1(n2468), .B0(n2383), .B1(
        top_core_EC_mc_n129), .Y(top_core_EC_mix_out_86_) );
  XOR2X1 U15946 ( .A(top_core_EC_mc_n57), .B(top_core_EC_mc_n130), .Y(
        top_core_EC_mc_n129) );
  XNOR2X1 U15947 ( .A(n1535), .B(top_core_EC_mc_n131), .Y(top_core_EC_mc_n128)
         );
  INVX1 U15948 ( .A(top_core_EC_mix_out_87_), .Y(n4777) );
  OAI22X1 U15949 ( .A0(top_core_EC_mc_n120), .A1(n2467), .B0(n2383), .B1(
        top_core_EC_mc_n121), .Y(top_core_EC_mix_out_87_) );
  XOR2X1 U15950 ( .A(top_core_EC_mc_n49), .B(top_core_EC_mc_n122), .Y(
        top_core_EC_mc_n121) );
  XNOR2X1 U15951 ( .A(n1534), .B(top_core_EC_mc_n123), .Y(top_core_EC_mc_n120)
         );
  INVX1 U15952 ( .A(top_core_EC_mix_out_88_), .Y(n4801) );
  OAI22X1 U15953 ( .A0(top_core_EC_mc_n112), .A1(n2446), .B0(n2384), .B1(
        top_core_EC_mc_n113), .Y(top_core_EC_mix_out_88_) );
  XOR2X1 U15954 ( .A(top_core_EC_mc_n114), .B(top_core_EC_mc_n115), .Y(
        top_core_EC_mc_n113) );
  XNOR2X1 U15955 ( .A(n1533), .B(top_core_EC_mc_n116), .Y(top_core_EC_mc_n112)
         );
  INVX1 U15956 ( .A(top_core_EC_mix_out_90_), .Y(n4796) );
  OAI22X1 U15957 ( .A0(top_core_EC_mc_n87), .A1(n2398), .B0(n2384), .B1(
        top_core_EC_mc_n88), .Y(top_core_EC_mix_out_90_) );
  XOR2X1 U15958 ( .A(top_core_EC_mc_n89), .B(top_core_EC_mc_n90), .Y(
        top_core_EC_mc_n88) );
  XNOR2X1 U15959 ( .A(top_core_EC_mc_mix_in_2_90_), .B(top_core_EC_mc_n91), 
        .Y(top_core_EC_mc_n87) );
  INVX1 U15960 ( .A(top_core_EC_mix_out_93_), .Y(n4781) );
  OAI22X1 U15961 ( .A0(top_core_EC_mc_n63), .A1(n2448), .B0(n2380), .B1(
        top_core_EC_mc_n64), .Y(top_core_EC_mix_out_93_) );
  XOR2X1 U15962 ( .A(top_core_EC_mc_n65), .B(top_core_EC_mc_n66), .Y(
        top_core_EC_mc_n64) );
  XNOR2X1 U15963 ( .A(top_core_EC_mc_mix_in_8[95]), .B(top_core_EC_mc_n67), 
        .Y(top_core_EC_mc_n63) );
  INVX1 U15964 ( .A(top_core_EC_mix_out_94_), .Y(n4785) );
  OAI22X1 U15965 ( .A0(top_core_EC_mc_n55), .A1(n2395), .B0(n2375), .B1(
        top_core_EC_mc_n56), .Y(top_core_EC_mix_out_94_) );
  XOR2X1 U15966 ( .A(top_core_EC_mc_n57), .B(top_core_EC_mc_n58), .Y(
        top_core_EC_mc_n56) );
  XNOR2X1 U15967 ( .A(n1535), .B(top_core_EC_mc_n59), .Y(top_core_EC_mc_n55)
         );
  INVX1 U15968 ( .A(top_core_EC_mix_out_95_), .Y(n4802) );
  OAI22X1 U15969 ( .A0(top_core_EC_mc_n47), .A1(n2460), .B0(n2375), .B1(
        top_core_EC_mc_n48), .Y(top_core_EC_mix_out_95_) );
  XOR2X1 U15970 ( .A(top_core_EC_mc_n49), .B(top_core_EC_mc_n50), .Y(
        top_core_EC_mc_n48) );
  XNOR2X1 U15971 ( .A(n1534), .B(top_core_EC_mc_n51), .Y(top_core_EC_mc_n47)
         );
  INVX1 U15972 ( .A(top_core_EC_mix_out_96_), .Y(n5149) );
  OAI22X1 U15973 ( .A0(top_core_EC_mc_n38), .A1(n2418), .B0(n2375), .B1(
        top_core_EC_mc_n39), .Y(top_core_EC_mix_out_96_) );
  XOR2X1 U15974 ( .A(top_core_EC_mc_n40), .B(top_core_EC_mc_n41), .Y(
        top_core_EC_mc_n39) );
  XNOR2X1 U15975 ( .A(top_core_EC_mix_in[120]), .B(top_core_EC_mc_n42), .Y(
        top_core_EC_mc_n38) );
  INVX1 U15976 ( .A(top_core_EC_mix_out_97_), .Y(n5140) );
  OAI22X1 U15977 ( .A0(top_core_EC_mc_n29), .A1(n2410), .B0(n2375), .B1(
        top_core_EC_mc_n30), .Y(top_core_EC_mix_out_97_) );
  XOR2X1 U15978 ( .A(top_core_EC_mc_n31), .B(top_core_EC_mc_n32), .Y(
        top_core_EC_mc_n30) );
  XNOR2X1 U15979 ( .A(top_core_EC_mc_mix_in_2_122_), .B(top_core_EC_mc_n33), 
        .Y(top_core_EC_mc_n29) );
  INVX1 U15980 ( .A(top_core_EC_mix_out_98_), .Y(n5144) );
  OAI22X1 U15981 ( .A0(top_core_EC_mc_n20), .A1(n2409), .B0(n2379), .B1(
        top_core_EC_mc_n21), .Y(top_core_EC_mix_out_98_) );
  XOR2X1 U15982 ( .A(top_core_EC_mc_n22), .B(top_core_EC_mc_n23), .Y(
        top_core_EC_mc_n21) );
  XNOR2X1 U15983 ( .A(top_core_EC_mix_in[122]), .B(top_core_EC_mc_n24), .Y(
        top_core_EC_mc_n20) );
  INVX1 U15984 ( .A(top_core_EC_mix_out_99_), .Y(n5138) );
  OAI22X1 U15985 ( .A0(top_core_EC_mc_n11), .A1(n2476), .B0(n2377), .B1(
        top_core_EC_mc_n12), .Y(top_core_EC_mix_out_99_) );
  XOR2X1 U15986 ( .A(top_core_EC_mc_n13), .B(top_core_EC_mc_n14), .Y(
        top_core_EC_mc_n12) );
  XNOR2X1 U15987 ( .A(top_core_EC_mix_in[123]), .B(top_core_EC_mc_n15), .Y(
        top_core_EC_mc_n11) );
  INVX1 U15988 ( .A(top_core_EC_mix_out_100_), .Y(n5126) );
  OAI22X1 U15989 ( .A0(top_core_EC_mc_n914), .A1(n2491), .B0(n2375), .B1(
        top_core_EC_mc_n915), .Y(top_core_EC_mix_out_100_) );
  XOR2X1 U15990 ( .A(top_core_EC_mc_n916), .B(top_core_EC_mc_n917), .Y(
        top_core_EC_mc_n915) );
  XNOR2X1 U15991 ( .A(top_core_EC_mc_mix_in_8[127]), .B(top_core_EC_mc_n918), 
        .Y(top_core_EC_mc_n914) );
  INVX1 U15992 ( .A(top_core_EC_mix_out_101_), .Y(n5128) );
  OAI22X1 U15993 ( .A0(top_core_EC_mc_n906), .A1(n2415), .B0(n2375), .B1(
        top_core_EC_mc_n907), .Y(top_core_EC_mix_out_101_) );
  XOR2X1 U15994 ( .A(top_core_EC_mc_n908), .B(top_core_EC_mc_n909), .Y(
        top_core_EC_mc_n907) );
  XNOR2X1 U15995 ( .A(n1553), .B(top_core_EC_mc_n910), .Y(top_core_EC_mc_n906)
         );
  INVX1 U15996 ( .A(top_core_EC_mix_out_102_), .Y(n5130) );
  OAI22X1 U15997 ( .A0(top_core_EC_mc_n898), .A1(n2426), .B0(n2375), .B1(
        top_core_EC_mc_n899), .Y(top_core_EC_mix_out_102_) );
  XOR2X1 U15998 ( .A(top_core_EC_mc_n900), .B(top_core_EC_mc_n901), .Y(
        top_core_EC_mc_n899) );
  XNOR2X1 U15999 ( .A(n1552), .B(top_core_EC_mc_n902), .Y(top_core_EC_mc_n898)
         );
  INVX1 U16000 ( .A(top_core_EC_mix_out_103_), .Y(n5150) );
  OAI22X1 U16001 ( .A0(top_core_EC_mc_n890), .A1(n2489), .B0(n2375), .B1(
        top_core_EC_mc_n891), .Y(top_core_EC_mix_out_103_) );
  XOR2X1 U16002 ( .A(top_core_EC_mc_n892), .B(top_core_EC_mc_n893), .Y(
        top_core_EC_mc_n891) );
  XNOR2X1 U16003 ( .A(n1551), .B(top_core_EC_mc_n894), .Y(top_core_EC_mc_n890)
         );
  INVX1 U16004 ( .A(top_core_EC_mix_out_104_), .Y(n5154) );
  OAI22X1 U16005 ( .A0(top_core_EC_mc_n883), .A1(n2433), .B0(n2376), .B1(
        top_core_EC_mc_n884), .Y(top_core_EC_mix_out_104_) );
  XOR2X1 U16006 ( .A(top_core_EC_mc_n885), .B(top_core_EC_mc_n886), .Y(
        top_core_EC_mc_n884) );
  XNOR2X1 U16007 ( .A(n1554), .B(top_core_EC_mc_n887), .Y(top_core_EC_mc_n883)
         );
  INVX1 U16008 ( .A(top_core_EC_mix_out_106_), .Y(n5146) );
  OAI22X1 U16009 ( .A0(top_core_EC_mc_n869), .A1(n2427), .B0(n2376), .B1(
        top_core_EC_mc_n870), .Y(top_core_EC_mix_out_106_) );
  XOR2X1 U16010 ( .A(top_core_EC_mc_n871), .B(top_core_EC_mc_n872), .Y(
        top_core_EC_mc_n870) );
  XNOR2X1 U16011 ( .A(top_core_EC_mc_mix_in_2_106_), .B(top_core_EC_mc_n873), 
        .Y(top_core_EC_mc_n869) );
  INVX1 U16012 ( .A(top_core_EC_mix_out_109_), .Y(n5135) );
  OAI22X1 U16013 ( .A0(top_core_EC_mc_n852), .A1(n2478), .B0(n2376), .B1(
        top_core_EC_mc_n853), .Y(top_core_EC_mix_out_109_) );
  XOR2X1 U16014 ( .A(top_core_EC_mc_n854), .B(top_core_EC_mc_n855), .Y(
        top_core_EC_mc_n853) );
  XNOR2X1 U16015 ( .A(top_core_EC_mc_mix_in_8[111]), .B(top_core_EC_mc_n856), 
        .Y(top_core_EC_mc_n852) );
  INVX1 U16016 ( .A(top_core_EC_mix_out_110_), .Y(n5131) );
  OAI22X1 U16017 ( .A0(top_core_EC_mc_n840), .A1(n2434), .B0(n2376), .B1(
        top_core_EC_mc_n841), .Y(top_core_EC_mix_out_110_) );
  XOR2X1 U16018 ( .A(top_core_EC_mc_n842), .B(top_core_EC_mc_n843), .Y(
        top_core_EC_mc_n841) );
  XNOR2X1 U16019 ( .A(n1556), .B(top_core_EC_mc_n844), .Y(top_core_EC_mc_n840)
         );
  INVX1 U16020 ( .A(top_core_EC_mix_out_111_), .Y(n5123) );
  OAI22X1 U16021 ( .A0(top_core_EC_mc_n835), .A1(n2456), .B0(n2376), .B1(
        top_core_EC_mc_n836), .Y(top_core_EC_mix_out_111_) );
  XOR2X1 U16022 ( .A(top_core_EC_mc_n837), .B(top_core_EC_mc_n838), .Y(
        top_core_EC_mc_n836) );
  XNOR2X1 U16023 ( .A(n1555), .B(top_core_EC_mc_n839), .Y(top_core_EC_mc_n835)
         );
  INVX1 U16024 ( .A(top_core_EC_mix_out_112_), .Y(n5153) );
  OAI22X1 U16025 ( .A0(top_core_EC_mc_n829), .A1(n2454), .B0(n2376), .B1(
        top_core_EC_mc_n830), .Y(top_core_EC_mix_out_112_) );
  XOR2X1 U16026 ( .A(top_core_EC_mc_n767), .B(top_core_EC_mc_n831), .Y(
        top_core_EC_mc_n830) );
  XNOR2X1 U16027 ( .A(n1551), .B(top_core_EC_mc_n832), .Y(top_core_EC_mc_n829)
         );
  INVX1 U16028 ( .A(top_core_EC_mix_out_114_), .Y(n5143) );
  OAI22X1 U16029 ( .A0(top_core_EC_mc_n817), .A1(n2477), .B0(n2376), .B1(
        top_core_EC_mc_n818), .Y(top_core_EC_mix_out_114_) );
  XOR2X1 U16030 ( .A(top_core_EC_mc_n753), .B(top_core_EC_mc_n819), .Y(
        top_core_EC_mc_n818) );
  XNOR2X1 U16031 ( .A(top_core_EC_mc_mix_in_2_122_), .B(top_core_EC_mc_n820), 
        .Y(top_core_EC_mc_n817) );
  INVX1 U16032 ( .A(top_core_EC_mix_out_117_), .Y(n5129) );
  OAI22X1 U16033 ( .A0(top_core_EC_mc_n795), .A1(n2479), .B0(n2377), .B1(
        top_core_EC_mc_n796), .Y(top_core_EC_mix_out_117_) );
  XOR2X1 U16034 ( .A(top_core_EC_mc_n730), .B(top_core_EC_mc_n797), .Y(
        top_core_EC_mc_n796) );
  XNOR2X1 U16035 ( .A(top_core_EC_mc_mix_in_8[127]), .B(top_core_EC_mc_n798), 
        .Y(top_core_EC_mc_n795) );
  INVX1 U16036 ( .A(top_core_EC_mix_out_118_), .Y(n5132) );
  OAI22X1 U16037 ( .A0(top_core_EC_mc_n787), .A1(n2461), .B0(n2377), .B1(
        top_core_EC_mc_n788), .Y(top_core_EC_mix_out_118_) );
  XOR2X1 U16038 ( .A(top_core_EC_mc_n722), .B(top_core_EC_mc_n789), .Y(
        top_core_EC_mc_n788) );
  XNOR2X1 U16039 ( .A(n1553), .B(top_core_EC_mc_n790), .Y(top_core_EC_mc_n787)
         );
  INVX1 U16040 ( .A(top_core_EC_mix_out_119_), .Y(n5125) );
  OAI22X1 U16041 ( .A0(top_core_EC_mc_n779), .A1(n2414), .B0(n2377), .B1(
        top_core_EC_mc_n780), .Y(top_core_EC_mix_out_119_) );
  XOR2X1 U16042 ( .A(top_core_EC_mc_n714), .B(top_core_EC_mc_n781), .Y(
        top_core_EC_mc_n780) );
  XNOR2X1 U16043 ( .A(n1552), .B(top_core_EC_mc_n782), .Y(top_core_EC_mc_n779)
         );
  INVX1 U16044 ( .A(top_core_EC_mix_out_120_), .Y(n5148) );
  OAI22X1 U16045 ( .A0(top_core_EC_mc_n765), .A1(n2397), .B0(n2377), .B1(
        top_core_EC_mc_n766), .Y(top_core_EC_mix_out_120_) );
  XOR2X1 U16046 ( .A(top_core_EC_mc_n767), .B(top_core_EC_mc_n768), .Y(
        top_core_EC_mc_n766) );
  XNOR2X1 U16047 ( .A(n1551), .B(top_core_EC_mc_n769), .Y(top_core_EC_mc_n765)
         );
  INVX1 U16048 ( .A(top_core_EC_mix_out_122_), .Y(n5147) );
  OAI22X1 U16049 ( .A0(top_core_EC_mc_n751), .A1(n2417), .B0(n2377), .B1(
        top_core_EC_mc_n752), .Y(top_core_EC_mix_out_122_) );
  XOR2X1 U16050 ( .A(top_core_EC_mc_n753), .B(top_core_EC_mc_n754), .Y(
        top_core_EC_mc_n752) );
  XNOR2X1 U16051 ( .A(top_core_EC_mc_mix_in_2_122_), .B(top_core_EC_mc_n755), 
        .Y(top_core_EC_mc_n751) );
  INVX1 U16052 ( .A(top_core_EC_mix_out_125_), .Y(n5136) );
  OAI22X1 U16053 ( .A0(top_core_EC_mc_n728), .A1(n2485), .B0(n2377), .B1(
        top_core_EC_mc_n729), .Y(top_core_EC_mix_out_125_) );
  XOR2X1 U16054 ( .A(top_core_EC_mc_n730), .B(top_core_EC_mc_n731), .Y(
        top_core_EC_mc_n729) );
  XNOR2X1 U16055 ( .A(top_core_EC_mc_mix_in_8[127]), .B(top_core_EC_mc_n732), 
        .Y(top_core_EC_mc_n728) );
  INVX1 U16056 ( .A(top_core_EC_mix_out_126_), .Y(n5133) );
  OAI22X1 U16057 ( .A0(top_core_EC_mc_n720), .A1(n2437), .B0(n2377), .B1(
        top_core_EC_mc_n721), .Y(top_core_EC_mix_out_126_) );
  XOR2X1 U16058 ( .A(top_core_EC_mc_n722), .B(top_core_EC_mc_n723), .Y(
        top_core_EC_mc_n721) );
  XNOR2X1 U16059 ( .A(n1553), .B(top_core_EC_mc_n724), .Y(top_core_EC_mc_n720)
         );
  INVX1 U16060 ( .A(top_core_EC_mix_out_127_), .Y(n5124) );
  OAI22X1 U16061 ( .A0(top_core_EC_mc_n712), .A1(n2462), .B0(n2377), .B1(
        top_core_EC_mc_n713), .Y(top_core_EC_mix_out_127_) );
  XOR2X1 U16062 ( .A(top_core_EC_mc_n714), .B(top_core_EC_mc_n715), .Y(
        top_core_EC_mc_n713) );
  XNOR2X1 U16063 ( .A(n1552), .B(top_core_EC_mc_n716), .Y(top_core_EC_mc_n712)
         );
  XNOR2X1 U16064 ( .A(top_core_EC_mc_mix_in_2_74_), .B(top_core_EC_mc_n165), 
        .Y(top_core_EC_mc_n220) );
  XNOR2X1 U16065 ( .A(top_core_EC_mc_mix_in_2_106_), .B(top_core_EC_mc_n26), 
        .Y(top_core_EC_mc_n871) );
  BUFX3 U16066 ( .A(n699), .Y(n1138) );
  BUFX3 U16067 ( .A(n698), .Y(n999) );
  BUFX3 U16068 ( .A(n700), .Y(n943) );
  BUFX3 U16069 ( .A(n701), .Y(n1083) );
  BUFX3 U16070 ( .A(n702), .Y(n1069) );
  BUFX3 U16071 ( .A(n704), .Y(n929) );
  BUFX3 U16072 ( .A(n703), .Y(n1013) );
  BUFX3 U16073 ( .A(n705), .Y(n1097) );
  BUFX3 U16074 ( .A(n706), .Y(n1027) );
  BUFX3 U16075 ( .A(n707), .Y(n957) );
  BUFX3 U16076 ( .A(n708), .Y(n1111) );
  BUFX3 U16077 ( .A(n709), .Y(n1041) );
  BUFX3 U16078 ( .A(n710), .Y(n971) );
  BUFX3 U16079 ( .A(n711), .Y(n1125) );
  BUFX3 U16080 ( .A(n712), .Y(n1055) );
  BUFX3 U16081 ( .A(n713), .Y(n985) );
  CLKINVX3 U16082 ( .A(n1708), .Y(n1703) );
  CLKINVX3 U16083 ( .A(n1737), .Y(n1732) );
  CLKINVX3 U16084 ( .A(n1678), .Y(n1674) );
  CLKINVX3 U16085 ( .A(n1814), .Y(n1810) );
  CLKINVX3 U16086 ( .A(n1835), .Y(n1831) );
  CLKINVX3 U16087 ( .A(n1793), .Y(n1789) );
  BUFX3 U16088 ( .A(n6603), .Y(n1160) );
  INVXL U16089 ( .A(n6), .Y(n6603) );
  XNOR2X1 U16090 ( .A(top_core_EC_mix_in[88]), .B(top_core_EC_mc_n181), .Y(
        top_core_EC_mc_n300) );
  XNOR2X1 U16091 ( .A(top_core_EC_mix_in[90]), .B(top_core_EC_mc_n165), .Y(
        top_core_EC_mc_n284) );
  XNOR2X1 U16092 ( .A(top_core_EC_mix_in[91]), .B(top_core_EC_mc_n157), .Y(
        top_core_EC_mc_n276) );
  XNOR2X1 U16093 ( .A(top_core_EC_mix_in[120]), .B(top_core_EC_mc_n44), .Y(
        top_core_EC_mc_n40) );
  XNOR2X1 U16094 ( .A(top_core_EC_mix_in[122]), .B(top_core_EC_mc_n26), .Y(
        top_core_EC_mc_n22) );
  XNOR2X1 U16095 ( .A(top_core_EC_mix_in[123]), .B(top_core_EC_mc_n17), .Y(
        top_core_EC_mc_n13) );
  AND2X2 U16096 ( .A(n2866), .B(n1000), .Y(n633) );
  AND2X2 U16097 ( .A(n3467), .B(n1140), .Y(n634) );
  AND2X2 U16098 ( .A(n2624), .B(n944), .Y(n635) );
  AND2X2 U16099 ( .A(n3226), .B(n1084), .Y(n636) );
  AND2X2 U16100 ( .A(n3165), .B(n1070), .Y(n637) );
  AND2X2 U16101 ( .A(n2563), .B(n930), .Y(n638) );
  AND2X2 U16102 ( .A(n2927), .B(n1014), .Y(n639) );
  AND2X2 U16103 ( .A(n3287), .B(n1098), .Y(n640) );
  AND2X2 U16104 ( .A(n2988), .B(n1028), .Y(n641) );
  AND2X2 U16105 ( .A(n2685), .B(n958), .Y(n642) );
  AND2X2 U16106 ( .A(n3348), .B(n1112), .Y(n643) );
  AND2X2 U16107 ( .A(n3046), .B(n1042), .Y(n644) );
  AND2X2 U16108 ( .A(n2745), .B(n972), .Y(n645) );
  AND2X2 U16109 ( .A(n3406), .B(n1126), .Y(n646) );
  AND2X2 U16110 ( .A(n3107), .B(n1056), .Y(n647) );
  AND2X2 U16111 ( .A(n2806), .B(n986), .Y(n648) );
  XOR2X1 U16112 ( .A(n1541), .B(top_core_EC_mc_mix_in_4_58_), .Y(
        top_core_EC_mc_mix_in_8[59]) );
  XOR2X1 U16113 ( .A(n1535), .B(top_core_EC_mc_mix_in_4_90_), .Y(
        top_core_EC_mc_mix_in_8[91]) );
  XNOR2X1 U16114 ( .A(n1535), .B(top_core_EC_mc_n141), .Y(top_core_EC_mc_n260)
         );
  XNOR2X1 U16115 ( .A(n1534), .B(top_core_EC_mc_n133), .Y(top_core_EC_mc_n243)
         );
  XNOR2X1 U16116 ( .A(n1553), .B(top_core_EC_mc_n800), .Y(top_core_EC_mc_n908)
         );
  XNOR2X1 U16117 ( .A(n1552), .B(top_core_EC_mc_n792), .Y(top_core_EC_mc_n900)
         );
  XNOR2X1 U16118 ( .A(n1538), .B(top_core_EC_mc_n133), .Y(top_core_EC_mc_n200)
         );
  XNOR2X1 U16119 ( .A(n1537), .B(top_core_EC_mc_n125), .Y(top_core_EC_mc_n195)
         );
  XNOR2X1 U16120 ( .A(n1556), .B(top_core_EC_mc_n792), .Y(top_core_EC_mc_n842)
         );
  XNOR2X1 U16121 ( .A(n1555), .B(top_core_EC_mc_n784), .Y(top_core_EC_mc_n837)
         );
  XNOR2X1 U16122 ( .A(n1533), .B(top_core_EC_mc_n125), .Y(top_core_EC_mc_n235)
         );
  XNOR2X1 U16123 ( .A(n1551), .B(top_core_EC_mc_n784), .Y(top_core_EC_mc_n892)
         );
  XNOR2X1 U16124 ( .A(n1536), .B(top_core_EC_mc_n181), .Y(top_core_EC_mc_n230)
         );
  XNOR2X1 U16125 ( .A(n1554), .B(top_core_EC_mc_n44), .Y(top_core_EC_mc_n885)
         );
  XOR2X1 U16126 ( .A(n1553), .B(top_core_EC_mc_mix_in_4_123_), .Y(
        top_core_EC_mc_mix_in_8[124]) );
  XOR2X1 U16127 ( .A(n1541), .B(n1540), .Y(top_core_EC_mc_mix_in_8[57]) );
  XOR2X1 U16128 ( .A(n1541), .B(top_core_EC_mc_mix_in_4_59_), .Y(
        top_core_EC_mc_mix_in_8[60]) );
  XOR2X1 U16129 ( .A(n1535), .B(n1534), .Y(top_core_EC_mc_mix_in_8[89]) );
  XOR2X1 U16130 ( .A(n1535), .B(top_core_EC_mc_mix_in_4_91_), .Y(
        top_core_EC_mc_mix_in_8[92]) );
  INVX1 U16131 ( .A(n13765), .Y(n6516) );
  INVX1 U16132 ( .A(n11874), .Y(n6823) );
  INVX1 U16133 ( .A(top_core_KE_sb1_n303), .Y(n6799) );
  INVX1 U16134 ( .A(n12190), .Y(n6502) );
  INVX1 U16135 ( .A(n12505), .Y(n6527) );
  INVX1 U16136 ( .A(n13450), .Y(n6467) );
  INVX1 U16137 ( .A(n12820), .Y(n6770) );
  INVX1 U16138 ( .A(n13135), .Y(n6812) );
  AOI222X1 U16139 ( .A0(n17288), .A1(n2848), .B0(n5326), .B1(n17289), .C0(
        n2847), .C1(n17290), .Y(n17271) );
  OAI21XL U16140 ( .A0(n17291), .A1(n2851), .B0(n17292), .Y(n17290) );
  OAI221XL U16141 ( .A0(n2860), .A1(n17296), .B0(n17047), .B1(n17208), .C0(
        n17297), .Y(n17288) );
  AOI222X1 U16142 ( .A0(n14138), .A1(n3449), .B0(n6108), .B1(n14139), .C0(
        n3448), .C1(n14140), .Y(n14121) );
  OAI21XL U16143 ( .A0(n14141), .A1(n3452), .B0(n14142), .Y(n14140) );
  OAI221XL U16144 ( .A0(n3460), .A1(n14146), .B0(n13897), .B1(n14058), .C0(
        n14147), .Y(n14138) );
  AOI222X1 U16145 ( .A0(n15398), .A1(n3208), .B0(n5798), .B1(n15399), .C0(
        n3207), .C1(n15400), .Y(n15381) );
  OAI21XL U16146 ( .A0(n15401), .A1(n3211), .B0(n15402), .Y(n15400) );
  OAI221XL U16147 ( .A0(n3220), .A1(n15406), .B0(n15157), .B1(n15318), .C0(
        n15407), .Y(n15398) );
  AOI222X1 U16148 ( .A0(n18548), .A1(n2606), .B0(n4972), .B1(n18549), .C0(
        n2605), .C1(n18550), .Y(n18531) );
  OAI21XL U16149 ( .A0(n18551), .A1(n2609), .B0(n18552), .Y(n18550) );
  OAI221XL U16150 ( .A0(n2618), .A1(n18556), .B0(n18307), .B1(n18468), .C0(
        n18557), .Y(n18548) );
  AOI222X1 U16151 ( .A0(n15713), .A1(n3147), .B0(n5714), .B1(n15714), .C0(
        n3146), .C1(n15715), .Y(n15696) );
  OAI21XL U16152 ( .A0(n15716), .A1(n3150), .B0(n15717), .Y(n15715) );
  OAI221XL U16153 ( .A0(n3159), .A1(n15721), .B0(n15472), .B1(n15633), .C0(
        n15722), .Y(n15713) );
  AOI222X1 U16154 ( .A0(n16973), .A1(n2909), .B0(n5410), .B1(n16974), .C0(
        n2908), .C1(n16975), .Y(n16956) );
  OAI21XL U16155 ( .A0(n16976), .A1(n2912), .B0(n16977), .Y(n16975) );
  OAI221XL U16156 ( .A0(n2921), .A1(n16981), .B0(n16732), .B1(n16893), .C0(
        n16982), .Y(n16973) );
  AOI222X1 U16157 ( .A0(n18863), .A1(n2545), .B0(n4856), .B1(n18864), .C0(
        n2544), .C1(n18865), .Y(n18846) );
  OAI21XL U16158 ( .A0(n18866), .A1(n2548), .B0(n18867), .Y(n18865) );
  OAI221XL U16159 ( .A0(n2557), .A1(n18871), .B0(n18622), .B1(n18783), .C0(
        n18872), .Y(n18863) );
  AOI222X1 U16160 ( .A0(n15083), .A1(n3269), .B0(n5874), .B1(n15084), .C0(
        n3268), .C1(n15085), .Y(n15066) );
  OAI21XL U16161 ( .A0(n15086), .A1(n3272), .B0(n15087), .Y(n15085) );
  OAI221XL U16162 ( .A0(n3281), .A1(n15091), .B0(n14842), .B1(n15003), .C0(
        n15092), .Y(n15083) );
  AOI222X1 U16163 ( .A0(n16658), .A1(n2970), .B0(n5486), .B1(n16659), .C0(
        n2969), .C1(n16660), .Y(n16641) );
  OAI21XL U16164 ( .A0(n16661), .A1(n2973), .B0(n16662), .Y(n16660) );
  OAI221XL U16165 ( .A0(n2982), .A1(n16666), .B0(n16417), .B1(n16578), .C0(
        n16667), .Y(n16658) );
  AOI222X1 U16166 ( .A0(n18233), .A1(n2667), .B0(n5056), .B1(n18234), .C0(
        n2666), .C1(n18235), .Y(n18216) );
  OAI21XL U16167 ( .A0(n18236), .A1(n2670), .B0(n18237), .Y(n18235) );
  OAI221XL U16168 ( .A0(n2679), .A1(n18241), .B0(n17992), .B1(n18153), .C0(
        n18242), .Y(n18233) );
  AOI222X1 U16169 ( .A0(n14768), .A1(n3330), .B0(n5950), .B1(n14769), .C0(
        n3329), .C1(n14770), .Y(n14751) );
  OAI21XL U16170 ( .A0(n14771), .A1(n3333), .B0(n14772), .Y(n14770) );
  OAI221XL U16171 ( .A0(n3342), .A1(n14776), .B0(n14527), .B1(n14688), .C0(
        n14777), .Y(n14768) );
  AOI222X1 U16172 ( .A0(n16343), .A1(n3028), .B0(n5562), .B1(n16344), .C0(
        n3027), .C1(n16345), .Y(n16326) );
  OAI21XL U16173 ( .A0(n16346), .A1(n3031), .B0(n16347), .Y(n16345) );
  OAI221XL U16174 ( .A0(n3040), .A1(n16351), .B0(n16102), .B1(n16263), .C0(
        n16352), .Y(n16343) );
  AOI222X1 U16175 ( .A0(n17918), .A1(n2727), .B0(n5164), .B1(n17919), .C0(
        n2726), .C1(n17920), .Y(n17901) );
  OAI21XL U16176 ( .A0(n17921), .A1(n2730), .B0(n17922), .Y(n17920) );
  OAI221XL U16177 ( .A0(n2739), .A1(n17926), .B0(n17677), .B1(n17838), .C0(
        n17927), .Y(n17918) );
  AOI222X1 U16178 ( .A0(n14453), .A1(n3388), .B0(n6026), .B1(n14454), .C0(
        n3387), .C1(n14455), .Y(n14436) );
  OAI21XL U16179 ( .A0(n14456), .A1(n3391), .B0(n14457), .Y(n14455) );
  OAI221XL U16180 ( .A0(n3400), .A1(n14461), .B0(n14212), .B1(n14373), .C0(
        n14462), .Y(n14453) );
  AOI222X1 U16181 ( .A0(n16028), .A1(n3089), .B0(n5638), .B1(n16029), .C0(
        n3088), .C1(n16030), .Y(n16011) );
  OAI21XL U16182 ( .A0(n16031), .A1(n3092), .B0(n16032), .Y(n16030) );
  OAI221XL U16183 ( .A0(n3101), .A1(n16036), .B0(n15787), .B1(n15948), .C0(
        n16037), .Y(n16028) );
  AOI222X1 U16184 ( .A0(n17603), .A1(n2788), .B0(n5242), .B1(n17604), .C0(
        n2787), .C1(n17605), .Y(n17586) );
  OAI21XL U16185 ( .A0(n17606), .A1(n2791), .B0(n17607), .Y(n17605) );
  OAI221XL U16186 ( .A0(n2800), .A1(n17611), .B0(n17362), .B1(n17523), .C0(
        n17612), .Y(n17603) );
  OAI21XL U16187 ( .A0(n3501), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n145), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n265), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n318) );
  OAI222XL U16188 ( .A0(n3494), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n70), 
        .B0(n1327), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n68), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n131), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n74), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n317) );
  OAI21XL U16189 ( .A0(n2900), .A1(n9960), .B0(n10079), .Y(n10132) );
  OAI222XL U16190 ( .A0(n2893), .A1(n9888), .B0(n1245), .B1(n9886), .C0(n9946), 
        .C1(n9891), .Y(n10131) );
  OAI21XL U16191 ( .A0(n2657), .A1(n11128), .B0(n11247), .Y(n11300) );
  OAI222XL U16192 ( .A0(n2650), .A1(n11056), .B0(n1253), .B1(n11054), .C0(
        n11114), .C1(n11059), .Y(n11299) );
  OAI21XL U16193 ( .A0(n3260), .A1(n8208), .B0(n8327), .Y(n8380) );
  OAI222XL U16194 ( .A0(n3253), .A1(n8136), .B0(n1233), .B1(n8134), .C0(n8194), 
        .C1(n8139), .Y(n8379) );
  OAI21XL U16195 ( .A0(n2718), .A1(n10836), .B0(n10955), .Y(n11008) );
  OAI222XL U16196 ( .A0(n2711), .A1(n10764), .B0(n1251), .B1(n10762), .C0(
        n10822), .C1(n10767), .Y(n11007) );
  OAI21XL U16197 ( .A0(n3079), .A1(n9084), .B0(n9203), .Y(n9256) );
  OAI222XL U16198 ( .A0(n3072), .A1(n9012), .B0(n1239), .B1(n9010), .C0(n9070), 
        .C1(n9015), .Y(n9255) );
  OAI21XL U16199 ( .A0(n3440), .A1(n7332), .B0(n7451), .Y(n7504) );
  OAI222XL U16200 ( .A0(n3433), .A1(n7260), .B0(n1227), .B1(n7258), .C0(n7318), 
        .C1(n7263), .Y(n7503) );
  OAI21XL U16201 ( .A0(n2843), .A1(n10252), .B0(n10371), .Y(n10424) );
  OAI222XL U16202 ( .A0(n2833), .A1(n10180), .B0(n1247), .B1(n10178), .C0(
        n10238), .C1(n10183), .Y(n10423) );
  OAI21XL U16203 ( .A0(n3018), .A1(n9376), .B0(n9495), .Y(n9548) );
  OAI222XL U16204 ( .A0(n3015), .A1(n9304), .B0(n1241), .B1(n9302), .C0(n9362), 
        .C1(n9307), .Y(n9547) );
  OAI21XL U16205 ( .A0(n3199), .A1(n8500), .B0(n8619), .Y(n8672) );
  OAI222XL U16206 ( .A0(n3192), .A1(n8428), .B0(n1235), .B1(n8426), .C0(n8486), 
        .C1(n8431), .Y(n8671) );
  OAI21XL U16207 ( .A0(n3378), .A1(n7624), .B0(n7743), .Y(n7796) );
  OAI222XL U16208 ( .A0(n3375), .A1(n7552), .B0(n1229), .B1(n7550), .C0(n7610), 
        .C1(n7555), .Y(n7795) );
  OAI21XL U16209 ( .A0(n2596), .A1(n11420), .B0(n11539), .Y(n11592) );
  OAI222XL U16210 ( .A0(n2599), .A1(n11348), .B0(n1255), .B1(n11346), .C0(
        n11406), .C1(n11351), .Y(n11591) );
  OAI21XL U16211 ( .A0(n2781), .A1(n10544), .B0(n10663), .Y(n10716) );
  OAI222XL U16212 ( .A0(n2772), .A1(n10472), .B0(n1249), .B1(n10470), .C0(
        n10530), .C1(n10475), .Y(n10715) );
  OAI21XL U16213 ( .A0(n2961), .A1(n9668), .B0(n9787), .Y(n9840) );
  OAI222XL U16214 ( .A0(n2954), .A1(n9596), .B0(n1243), .B1(n9594), .C0(n9654), 
        .C1(n9599), .Y(n9839) );
  OAI21XL U16215 ( .A0(n3137), .A1(n8792), .B0(n8911), .Y(n8964) );
  OAI222XL U16216 ( .A0(n3134), .A1(n8720), .B0(n1237), .B1(n8718), .C0(n8778), 
        .C1(n8723), .Y(n8963) );
  OAI21XL U16217 ( .A0(n3323), .A1(n7916), .B0(n8035), .Y(n8088) );
  OAI222XL U16218 ( .A0(n3314), .A1(n7844), .B0(n1231), .B1(n7842), .C0(n7902), 
        .C1(n7847), .Y(n8087) );
  OAI2BB1X1 U16219 ( .A0N(n9913), .A1N(n135), .B0(n9999), .Y(n10031) );
  OAI222XL U16220 ( .A0(n2881), .A1(n15), .B0(n2893), .B1(n9944), .C0(n10032), 
        .C1(n2887), .Y(n10030) );
  OAI2BB1X1 U16221 ( .A0N(top_core_EC_ss_gen_tbox_0__sboxs_r_n97), .A1N(n136), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n185), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n217) );
  OAI222XL U16222 ( .A0(n3482), .A1(n14), .B0(n3494), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n129), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n218), .C1(n3489), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n216) );
  OAI2BB1X1 U16223 ( .A0N(n11081), .A1N(n137), .B0(n11167), .Y(n11199) );
  OAI222XL U16224 ( .A0(n2639), .A1(n16), .B0(n2650), .B1(n11112), .C0(n11200), 
        .C1(n2642), .Y(n11198) );
  OAI2BB1X1 U16225 ( .A0N(n8161), .A1N(n138), .B0(n8247), .Y(n8279) );
  OAI222XL U16226 ( .A0(n3241), .A1(n17), .B0(n3253), .B1(n8192), .C0(n8280), 
        .C1(n3251), .Y(n8278) );
  OAI2BB1X1 U16227 ( .A0N(n10789), .A1N(n139), .B0(n10875), .Y(n10907) );
  OAI222XL U16228 ( .A0(n2700), .A1(n18), .B0(n2711), .B1(n10820), .C0(n10908), 
        .C1(n2704), .Y(n10906) );
  OAI2BB1X1 U16229 ( .A0N(n9037), .A1N(n140), .B0(n9123), .Y(n9155) );
  OAI222XL U16230 ( .A0(n3061), .A1(n19), .B0(n3072), .B1(n9068), .C0(n9156), 
        .C1(n3065), .Y(n9154) );
  OAI2BB1X1 U16231 ( .A0N(n7285), .A1N(n141), .B0(n7371), .Y(n7403) );
  OAI222XL U16232 ( .A0(n3421), .A1(n20), .B0(n3433), .B1(n7316), .C0(n7404), 
        .C1(n3424), .Y(n7402) );
  OAI2BB1X1 U16233 ( .A0N(n10205), .A1N(n142), .B0(n10291), .Y(n10323) );
  OAI222XL U16234 ( .A0(n2821), .A1(n21), .B0(n2833), .B1(n10236), .C0(n10324), 
        .C1(n2825), .Y(n10322) );
  OAI2BB1X1 U16235 ( .A0N(n9329), .A1N(n143), .B0(n9415), .Y(n9447) );
  OAI222XL U16236 ( .A0(n3003), .A1(n22), .B0(n3015), .B1(n9360), .C0(n9448), 
        .C1(n3013), .Y(n9446) );
  OAI2BB1X1 U16237 ( .A0N(n8453), .A1N(n144), .B0(n8539), .Y(n8571) );
  OAI222XL U16238 ( .A0(n3180), .A1(n23), .B0(n3192), .B1(n8484), .C0(n8572), 
        .C1(n3184), .Y(n8570) );
  OAI2BB1X1 U16239 ( .A0N(n7577), .A1N(n145), .B0(n7663), .Y(n7695) );
  OAI222XL U16240 ( .A0(n3363), .A1(n24), .B0(n3375), .B1(n7608), .C0(n7696), 
        .C1(n3367), .Y(n7694) );
  OAI2BB1X1 U16241 ( .A0N(n11373), .A1N(n146), .B0(n11459), .Y(n11491) );
  OAI222XL U16242 ( .A0(n2578), .A1(n25), .B0(n2600), .B1(n11404), .C0(n11492), 
        .C1(n2582), .Y(n11490) );
  OAI2BB1X1 U16243 ( .A0N(n10497), .A1N(n147), .B0(n10583), .Y(n10615) );
  OAI222XL U16244 ( .A0(n2760), .A1(n26), .B0(n2772), .B1(n10528), .C0(n10616), 
        .C1(n2764), .Y(n10614) );
  OAI2BB1X1 U16245 ( .A0N(n9621), .A1N(n148), .B0(n9707), .Y(n9739) );
  OAI222XL U16246 ( .A0(n2942), .A1(n27), .B0(n2954), .B1(n9652), .C0(n9740), 
        .C1(n2946), .Y(n9738) );
  OAI2BB1X1 U16247 ( .A0N(n8745), .A1N(n149), .B0(n8831), .Y(n8863) );
  OAI222XL U16248 ( .A0(n3122), .A1(n28), .B0(n3134), .B1(n8776), .C0(n8864), 
        .C1(n3126), .Y(n8862) );
  OAI2BB1X1 U16249 ( .A0N(n7869), .A1N(n150), .B0(n7955), .Y(n7987) );
  OAI222XL U16250 ( .A0(n3302), .A1(n29), .B0(n3314), .B1(n7900), .C0(n7988), 
        .C1(n3312), .Y(n7986) );
  INVX1 U16251 ( .A(n11756), .Y(n6911) );
  INVX1 U16252 ( .A(top_core_KE_sb1_n184), .Y(n6865) );
  INVX1 U16253 ( .A(n12387), .Y(n6618) );
  INVX1 U16254 ( .A(n12072), .Y(n6571) );
  AND3X2 U16255 ( .A(n13894), .B(n13895), .C(n13896), .Y(n13893) );
  AND3X2 U16256 ( .A(n17044), .B(n17045), .C(n17046), .Y(n17043) );
  AND3X2 U16257 ( .A(n18304), .B(n18305), .C(n18306), .Y(n18303) );
  AND3X2 U16258 ( .A(n15154), .B(n15155), .C(n15156), .Y(n15153) );
  AND3X2 U16259 ( .A(n15469), .B(n15470), .C(n15471), .Y(n15468) );
  AND3X2 U16260 ( .A(n18619), .B(n18620), .C(n18621), .Y(n18618) );
  AND3X2 U16261 ( .A(n16729), .B(n16730), .C(n16731), .Y(n16728) );
  AND3X2 U16262 ( .A(n14839), .B(n14840), .C(n14841), .Y(n14838) );
  AND3X2 U16263 ( .A(n16414), .B(n16415), .C(n16416), .Y(n16413) );
  AND3X2 U16264 ( .A(n17989), .B(n17990), .C(n17991), .Y(n17988) );
  AND3X2 U16265 ( .A(n14524), .B(n14525), .C(n14526), .Y(n14523) );
  AND3X2 U16266 ( .A(n16099), .B(n16100), .C(n16101), .Y(n16098) );
  AND3X2 U16267 ( .A(n17674), .B(n17675), .C(n17676), .Y(n17673) );
  AND3X2 U16268 ( .A(n14209), .B(n14210), .C(n14211), .Y(n14208) );
  AND3X2 U16269 ( .A(n15784), .B(n15785), .C(n15786), .Y(n15783) );
  AND3X2 U16270 ( .A(n17359), .B(n17360), .C(n17361), .Y(n17358) );
  CLKINVX3 U16271 ( .A(n3705), .Y(n3704) );
  AOI221X1 U16272 ( .A0(n2858), .A1(n9971), .B0(n9972), .B1(n2864), .C0(n9973), 
        .Y(n9931) );
  NAND2X1 U16273 ( .A(n9947), .B(n9974), .Y(n9973) );
  OAI221XL U16274 ( .A0(n9976), .A1(n9970), .B0(n9945), .B1(n9918), .C0(n9949), 
        .Y(n9971) );
  OAI221XL U16275 ( .A0(n2881), .A1(n9887), .B0(n9893), .B1(n1245), .C0(n9975), 
        .Y(n9972) );
  AOI221X1 U16276 ( .A0(n3457), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n157), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n158), .B1(n3465), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n159), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n116) );
  NAND2X1 U16277 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n132), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n160), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n159) );
  OAI221XL U16278 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n162), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n130), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n102), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n134), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n157) );
  OAI221XL U16279 ( .A0(n3482), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n69), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n76), .B1(n1327), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n161), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n158) );
  AOI221X1 U16280 ( .A0(n2615), .A1(n11139), .B0(n11140), .B1(n2622), .C0(
        n11141), .Y(n11099) );
  NAND2X1 U16281 ( .A(n11115), .B(n11142), .Y(n11141) );
  OAI221XL U16282 ( .A0(n11144), .A1(n11138), .B0(n11113), .B1(n11086), .C0(
        n11117), .Y(n11139) );
  OAI221XL U16283 ( .A0(n2639), .A1(n11055), .B0(n11061), .B1(n1253), .C0(
        n11143), .Y(n11140) );
  AOI221X1 U16284 ( .A0(n3218), .A1(n8219), .B0(n8220), .B1(n3224), .C0(n8221), 
        .Y(n8179) );
  NAND2X1 U16285 ( .A(n8195), .B(n8222), .Y(n8221) );
  OAI221XL U16286 ( .A0(n8224), .A1(n8218), .B0(n8193), .B1(n8166), .C0(n8197), 
        .Y(n8219) );
  OAI221XL U16287 ( .A0(n3241), .A1(n8135), .B0(n8141), .B1(n1233), .C0(n8223), 
        .Y(n8220) );
  AOI221X1 U16288 ( .A0(n2677), .A1(n10847), .B0(n10848), .B1(n2683), .C0(
        n10849), .Y(n10807) );
  NAND2X1 U16289 ( .A(n10823), .B(n10850), .Y(n10849) );
  OAI221XL U16290 ( .A0(n10852), .A1(n10846), .B0(n10821), .B1(n10794), .C0(
        n10825), .Y(n10847) );
  OAI221XL U16291 ( .A0(n2700), .A1(n10763), .B0(n10769), .B1(n1251), .C0(
        n10851), .Y(n10848) );
  AOI221X1 U16292 ( .A0(n3037), .A1(n9095), .B0(n9096), .B1(n3044), .C0(n9097), 
        .Y(n9055) );
  NAND2X1 U16293 ( .A(n9071), .B(n9098), .Y(n9097) );
  OAI221XL U16294 ( .A0(n9100), .A1(n9094), .B0(n9069), .B1(n9042), .C0(n9073), 
        .Y(n9095) );
  OAI221XL U16295 ( .A0(n3061), .A1(n9011), .B0(n9017), .B1(n1239), .C0(n9099), 
        .Y(n9096) );
  AOI221X1 U16296 ( .A0(n3397), .A1(n7343), .B0(n7344), .B1(n3404), .C0(n7345), 
        .Y(n7303) );
  NAND2X1 U16297 ( .A(n7319), .B(n7346), .Y(n7345) );
  OAI221XL U16298 ( .A0(n7348), .A1(n7342), .B0(n7317), .B1(n7290), .C0(n7321), 
        .Y(n7343) );
  OAI221XL U16299 ( .A0(n3421), .A1(n7259), .B0(n7265), .B1(n1227), .C0(n7347), 
        .Y(n7344) );
  AOI221X1 U16300 ( .A0(n2797), .A1(n10263), .B0(n10264), .B1(n2804), .C0(
        n10265), .Y(n10223) );
  NAND2X1 U16301 ( .A(n10239), .B(n10266), .Y(n10265) );
  OAI221XL U16302 ( .A0(n10268), .A1(n10262), .B0(n10237), .B1(n10210), .C0(
        n10241), .Y(n10263) );
  OAI221XL U16303 ( .A0(n2821), .A1(n10179), .B0(n10185), .B1(n1247), .C0(
        n10267), .Y(n10264) );
  AOI221X1 U16304 ( .A0(n2979), .A1(n9387), .B0(n9388), .B1(n2986), .C0(n9389), 
        .Y(n9347) );
  NAND2X1 U16305 ( .A(n9363), .B(n9390), .Y(n9389) );
  OAI221XL U16306 ( .A0(n9392), .A1(n9386), .B0(n9361), .B1(n9334), .C0(n9365), 
        .Y(n9387) );
  OAI221XL U16307 ( .A0(n3003), .A1(n9303), .B0(n9309), .B1(n1241), .C0(n9391), 
        .Y(n9388) );
  AOI221X1 U16308 ( .A0(n3156), .A1(n8511), .B0(n8512), .B1(n3163), .C0(n8513), 
        .Y(n8471) );
  NAND2X1 U16309 ( .A(n8487), .B(n8514), .Y(n8513) );
  OAI221XL U16310 ( .A0(n8516), .A1(n8510), .B0(n8485), .B1(n8458), .C0(n8489), 
        .Y(n8511) );
  OAI221XL U16311 ( .A0(n3180), .A1(n8427), .B0(n8433), .B1(n1235), .C0(n8515), 
        .Y(n8512) );
  AOI221X1 U16312 ( .A0(n3339), .A1(n7635), .B0(n7636), .B1(n3346), .C0(n7637), 
        .Y(n7595) );
  NAND2X1 U16313 ( .A(n7611), .B(n7638), .Y(n7637) );
  OAI221XL U16314 ( .A0(n7640), .A1(n7634), .B0(n7609), .B1(n7582), .C0(n7613), 
        .Y(n7635) );
  OAI221XL U16315 ( .A0(n3363), .A1(n7551), .B0(n7557), .B1(n1229), .C0(n7639), 
        .Y(n7636) );
  AOI221X1 U16316 ( .A0(n2559), .A1(n11431), .B0(n11432), .B1(n2549), .C0(
        n11433), .Y(n11391) );
  NAND2X1 U16317 ( .A(n11407), .B(n11434), .Y(n11433) );
  OAI221XL U16318 ( .A0(n11436), .A1(n11430), .B0(n11405), .B1(n11378), .C0(
        n11409), .Y(n11431) );
  OAI221XL U16319 ( .A0(n2578), .A1(n11347), .B0(n11353), .B1(n1255), .C0(
        n11435), .Y(n11432) );
  AOI221X1 U16320 ( .A0(n2737), .A1(n10555), .B0(n10556), .B1(n2743), .C0(
        n10557), .Y(n10515) );
  NAND2X1 U16321 ( .A(n10531), .B(n10558), .Y(n10557) );
  OAI221XL U16322 ( .A0(n10560), .A1(n10554), .B0(n10529), .B1(n10502), .C0(
        n10533), .Y(n10555) );
  OAI221XL U16323 ( .A0(n2760), .A1(n10471), .B0(n10477), .B1(n1249), .C0(
        n10559), .Y(n10556) );
  AOI221X1 U16324 ( .A0(n2918), .A1(n9679), .B0(n9680), .B1(n2925), .C0(n9681), 
        .Y(n9639) );
  NAND2X1 U16325 ( .A(n9655), .B(n9682), .Y(n9681) );
  OAI221XL U16326 ( .A0(n9684), .A1(n9678), .B0(n9653), .B1(n9626), .C0(n9657), 
        .Y(n9679) );
  OAI221XL U16327 ( .A0(n2942), .A1(n9595), .B0(n9601), .B1(n1243), .C0(n9683), 
        .Y(n9680) );
  AOI221X1 U16328 ( .A0(n3099), .A1(n8803), .B0(n8804), .B1(n3105), .C0(n8805), 
        .Y(n8763) );
  NAND2X1 U16329 ( .A(n8779), .B(n8806), .Y(n8805) );
  OAI221XL U16330 ( .A0(n8808), .A1(n8802), .B0(n8777), .B1(n8750), .C0(n8781), 
        .Y(n8803) );
  OAI221XL U16331 ( .A0(n3122), .A1(n8719), .B0(n8725), .B1(n1237), .C0(n8807), 
        .Y(n8804) );
  AOI221X1 U16332 ( .A0(n3278), .A1(n7927), .B0(n7928), .B1(n3285), .C0(n7929), 
        .Y(n7887) );
  NAND2X1 U16333 ( .A(n7903), .B(n7930), .Y(n7929) );
  OAI221XL U16334 ( .A0(n7932), .A1(n7926), .B0(n7901), .B1(n7874), .C0(n7905), 
        .Y(n7927) );
  OAI221XL U16335 ( .A0(n3302), .A1(n7843), .B0(n7849), .B1(n1231), .C0(n7931), 
        .Y(n7928) );
  AOI221X1 U16336 ( .A0(n5321), .A1(n9936), .B0(n9909), .B1(n9937), .C0(n9938), 
        .Y(n9935) );
  AOI21X1 U16337 ( .A0(n9939), .A1(n9940), .B0(n2850), .Y(n9938) );
  OAI221XL U16338 ( .A0(n1004), .A1(n9917), .B0(n465), .B1(n9886), .C0(n9959), 
        .Y(n9937) );
  AOI221X1 U16339 ( .A0(n6105), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n121), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n93), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n122), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n123), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n120) );
  AOI21X1 U16340 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n124), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n125), .B0(n3451), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n123) );
  OAI221XL U16341 ( .A0(n1145), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n101), 
        .B0(n466), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n68), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n144), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n122) );
  AOI221X1 U16342 ( .A0(n4967), .A1(n11104), .B0(n11077), .B1(n11105), .C0(
        n11106), .Y(n11103) );
  AOI21X1 U16343 ( .A0(n11107), .A1(n11108), .B0(n2608), .Y(n11106) );
  OAI221XL U16344 ( .A0(n948), .A1(n11085), .B0(n467), .B1(n11054), .C0(n11127), .Y(n11105) );
  AOI221X1 U16345 ( .A0(n5793), .A1(n8184), .B0(n8157), .B1(n8185), .C0(n8186), 
        .Y(n8183) );
  AOI21X1 U16346 ( .A0(n8187), .A1(n8188), .B0(n3210), .Y(n8186) );
  OAI221XL U16347 ( .A0(n1088), .A1(n8165), .B0(n468), .B1(n8134), .C0(n8207), 
        .Y(n8185) );
  AOI221X1 U16348 ( .A0(n5051), .A1(n10812), .B0(n10785), .B1(n10813), .C0(
        n10814), .Y(n10811) );
  AOI21X1 U16349 ( .A0(n10815), .A1(n10816), .B0(n2669), .Y(n10814) );
  OAI221XL U16350 ( .A0(n962), .A1(n10793), .B0(n474), .B1(n10762), .C0(n10835), .Y(n10813) );
  AOI221X1 U16351 ( .A0(n5557), .A1(n9060), .B0(n9033), .B1(n9061), .C0(n9062), 
        .Y(n9059) );
  AOI21X1 U16352 ( .A0(n9063), .A1(n9064), .B0(n3030), .Y(n9062) );
  OAI221XL U16353 ( .A0(n1046), .A1(n9041), .B0(n476), .B1(n9010), .C0(n9083), 
        .Y(n9061) );
  AOI221X1 U16354 ( .A0(n6021), .A1(n7308), .B0(n7281), .B1(n7309), .C0(n7310), 
        .Y(n7307) );
  AOI21X1 U16355 ( .A0(n7311), .A1(n7312), .B0(n3390), .Y(n7310) );
  OAI221XL U16356 ( .A0(n1130), .A1(n7289), .B0(n478), .B1(n7258), .C0(n7331), 
        .Y(n7309) );
  AOI221X1 U16357 ( .A0(n5237), .A1(n10228), .B0(n10201), .B1(n10229), .C0(
        n10230), .Y(n10227) );
  AOI21X1 U16358 ( .A0(n10231), .A1(n10232), .B0(n2790), .Y(n10230) );
  OAI221XL U16359 ( .A0(n990), .A1(n10209), .B0(n480), .B1(n10178), .C0(n10251), .Y(n10229) );
  AOI221X1 U16360 ( .A0(n5481), .A1(n9352), .B0(n9325), .B1(n9353), .C0(n9354), 
        .Y(n9351) );
  AOI21X1 U16361 ( .A0(n9355), .A1(n9356), .B0(n2972), .Y(n9354) );
  OAI221XL U16362 ( .A0(n1032), .A1(n9333), .B0(n473), .B1(n9302), .C0(n9375), 
        .Y(n9353) );
  AOI221X1 U16363 ( .A0(n5709), .A1(n8476), .B0(n8449), .B1(n8477), .C0(n8478), 
        .Y(n8475) );
  AOI21X1 U16364 ( .A0(n8479), .A1(n8480), .B0(n3149), .Y(n8478) );
  OAI221XL U16365 ( .A0(n1074), .A1(n8457), .B0(n469), .B1(n8426), .C0(n8499), 
        .Y(n8477) );
  AOI221X1 U16366 ( .A0(n5945), .A1(n7600), .B0(n7573), .B1(n7601), .C0(n7602), 
        .Y(n7599) );
  AOI21X1 U16367 ( .A0(n7603), .A1(n7604), .B0(n3332), .Y(n7602) );
  OAI221XL U16368 ( .A0(n1116), .A1(n7581), .B0(n475), .B1(n7550), .C0(n7623), 
        .Y(n7601) );
  AOI221X1 U16369 ( .A0(n4851), .A1(n11396), .B0(n11369), .B1(n11397), .C0(
        n11398), .Y(n11395) );
  AOI21X1 U16370 ( .A0(n11399), .A1(n11400), .B0(n2547), .Y(n11398) );
  OAI221XL U16371 ( .A0(n934), .A1(n11377), .B0(n471), .B1(n11346), .C0(n11419), .Y(n11397) );
  AOI221X1 U16372 ( .A0(n5159), .A1(n10520), .B0(n10493), .B1(n10521), .C0(
        n10522), .Y(n10519) );
  AOI21X1 U16373 ( .A0(n10523), .A1(n10524), .B0(n2729), .Y(n10522) );
  OAI221XL U16374 ( .A0(n976), .A1(n10501), .B0(n477), .B1(n10470), .C0(n10543), .Y(n10521) );
  AOI221X1 U16375 ( .A0(n5405), .A1(n9644), .B0(n9617), .B1(n9645), .C0(n9646), 
        .Y(n9643) );
  AOI21X1 U16376 ( .A0(n9647), .A1(n9648), .B0(n2911), .Y(n9646) );
  OAI221XL U16377 ( .A0(n1018), .A1(n9625), .B0(n470), .B1(n9594), .C0(n9667), 
        .Y(n9645) );
  AOI221X1 U16378 ( .A0(n5633), .A1(n8768), .B0(n8741), .B1(n8769), .C0(n8770), 
        .Y(n8767) );
  AOI21X1 U16379 ( .A0(n8771), .A1(n8772), .B0(n3091), .Y(n8770) );
  OAI221XL U16380 ( .A0(n1060), .A1(n8749), .B0(n479), .B1(n8718), .C0(n8791), 
        .Y(n8769) );
  AOI221X1 U16381 ( .A0(n5869), .A1(n7892), .B0(n7865), .B1(n7893), .C0(n7894), 
        .Y(n7891) );
  AOI21X1 U16382 ( .A0(n7895), .A1(n7896), .B0(n3271), .Y(n7894) );
  OAI221XL U16383 ( .A0(n1102), .A1(n7873), .B0(n472), .B1(n7842), .C0(n7915), 
        .Y(n7893) );
  AND2X2 U16384 ( .A(n1802), .B(n1812), .Y(n665) );
  AND2X2 U16385 ( .A(n1823), .B(n1833), .Y(n666) );
  AND2X2 U16386 ( .A(n1760), .B(n1773), .Y(n667) );
  AND2X2 U16387 ( .A(n1781), .B(n1791), .Y(n668) );
  AND2X2 U16388 ( .A(n1651), .B(n1664), .Y(n669) );
  AND2X2 U16389 ( .A(n1680), .B(n1692), .Y(n670) );
  AND2X2 U16390 ( .A(n1738), .B(n1750), .Y(n671) );
  AND2X2 U16391 ( .A(n1709), .B(n1721), .Y(n672) );
  AOI221X1 U16392 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n65), .A1(n3454), 
        .B0(n3464), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n66), .C0(n6134), 
        .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n64) );
  INVX1 U16393 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n67), .Y(n6134) );
  OAI221XL U16394 ( .A0(n3482), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n71), 
        .B0(n1625), .B1(n14), .C0(top_core_EC_ss_gen_tbox_0__sboxs_r_n73), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n65) );
  OAI221XL U16395 ( .A0(n3499), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n68), 
        .B0(n3494), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n69), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n70), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n66) );
  AOI221X1 U16396 ( .A0(n9883), .A1(n2853), .B0(n2855), .B1(n9884), .C0(n5338), 
        .Y(n9882) );
  INVX1 U16397 ( .A(n9885), .Y(n5338) );
  OAI221XL U16398 ( .A0(n2881), .A1(n9889), .B0(n1615), .B1(n15), .C0(n9890), 
        .Y(n9883) );
  OAI221XL U16399 ( .A0(n2898), .A1(n9886), .B0(n2893), .B1(n9887), .C0(n9888), 
        .Y(n9884) );
  AOI221X1 U16400 ( .A0(n11051), .A1(n2611), .B0(n2613), .B1(n11052), .C0(
        n4984), .Y(n11050) );
  INVX1 U16401 ( .A(n11053), .Y(n4984) );
  OAI221XL U16402 ( .A0(n2639), .A1(n11057), .B0(n1611), .B1(n16), .C0(n11058), 
        .Y(n11051) );
  OAI221XL U16403 ( .A0(n2655), .A1(n11054), .B0(n2650), .B1(n11055), .C0(
        n11056), .Y(n11052) );
  AOI221X1 U16404 ( .A0(n8131), .A1(n3213), .B0(n3215), .B1(n8132), .C0(n5810), 
        .Y(n8130) );
  INVX1 U16405 ( .A(n8133), .Y(n5810) );
  OAI221XL U16406 ( .A0(n3241), .A1(n8137), .B0(n1621), .B1(n17), .C0(n8138), 
        .Y(n8131) );
  OAI221XL U16407 ( .A0(n3258), .A1(n8134), .B0(n3253), .B1(n8135), .C0(n8136), 
        .Y(n8132) );
  AOI221X1 U16408 ( .A0(n10759), .A1(n2672), .B0(n2674), .B1(n10760), .C0(
        n5068), .Y(n10758) );
  INVX1 U16409 ( .A(n10761), .Y(n5068) );
  OAI221XL U16410 ( .A0(n2700), .A1(n10765), .B0(n1612), .B1(n18), .C0(n10766), 
        .Y(n10759) );
  OAI221XL U16411 ( .A0(n2716), .A1(n10762), .B0(n2711), .B1(n10763), .C0(
        n10764), .Y(n10760) );
  AOI221X1 U16412 ( .A0(n9007), .A1(n3033), .B0(n3035), .B1(n9008), .C0(n5574), 
        .Y(n9006) );
  INVX1 U16413 ( .A(n9009), .Y(n5574) );
  OAI221XL U16414 ( .A0(n3061), .A1(n9013), .B0(n1618), .B1(n19), .C0(n9014), 
        .Y(n9007) );
  OAI221XL U16415 ( .A0(n3077), .A1(n9010), .B0(n3072), .B1(n9011), .C0(n9012), 
        .Y(n9008) );
  AOI221X1 U16416 ( .A0(n7255), .A1(n3393), .B0(n3395), .B1(n7256), .C0(n6038), 
        .Y(n7254) );
  INVX1 U16417 ( .A(n7257), .Y(n6038) );
  OAI221XL U16418 ( .A0(n3421), .A1(n7261), .B0(n1624), .B1(n20), .C0(n7262), 
        .Y(n7255) );
  OAI221XL U16419 ( .A0(n3438), .A1(n7258), .B0(n3433), .B1(n7259), .C0(n7260), 
        .Y(n7256) );
  AOI221X1 U16420 ( .A0(n10175), .A1(n2793), .B0(n2795), .B1(n10176), .C0(
        n5254), .Y(n10174) );
  INVX1 U16421 ( .A(n10177), .Y(n5254) );
  OAI221XL U16422 ( .A0(n2821), .A1(n10181), .B0(n1614), .B1(n21), .C0(n10182), 
        .Y(n10175) );
  OAI221XL U16423 ( .A0(n2841), .A1(n10178), .B0(n2833), .B1(n10179), .C0(
        n10180), .Y(n10176) );
  AOI221X1 U16424 ( .A0(n9299), .A1(n2975), .B0(n2977), .B1(n9300), .C0(n5498), 
        .Y(n9298) );
  INVX1 U16425 ( .A(n9301), .Y(n5498) );
  OAI221XL U16426 ( .A0(n3003), .A1(n9305), .B0(n1617), .B1(n22), .C0(n9306), 
        .Y(n9299) );
  OAI221XL U16427 ( .A0(n3022), .A1(n9302), .B0(n3015), .B1(n9303), .C0(n9304), 
        .Y(n9300) );
  AOI221X1 U16428 ( .A0(n8423), .A1(n3152), .B0(n3154), .B1(n8424), .C0(n5726), 
        .Y(n8422) );
  INVX1 U16429 ( .A(n8425), .Y(n5726) );
  OAI221XL U16430 ( .A0(n3180), .A1(n8429), .B0(n1620), .B1(n23), .C0(n8430), 
        .Y(n8423) );
  OAI221XL U16431 ( .A0(n3197), .A1(n8426), .B0(n3192), .B1(n8427), .C0(n8428), 
        .Y(n8424) );
  AOI221X1 U16432 ( .A0(n7547), .A1(n3335), .B0(n3337), .B1(n7548), .C0(n5962), 
        .Y(n7546) );
  INVX1 U16433 ( .A(n7549), .Y(n5962) );
  OAI221XL U16434 ( .A0(n3363), .A1(n7553), .B0(n1623), .B1(n24), .C0(n7554), 
        .Y(n7547) );
  OAI221XL U16435 ( .A0(n3382), .A1(n7550), .B0(n3375), .B1(n7551), .C0(n7552), 
        .Y(n7548) );
  AOI221X1 U16436 ( .A0(n11343), .A1(n2550), .B0(n2559), .B1(n11344), .C0(
        n4868), .Y(n11342) );
  INVX1 U16437 ( .A(n11345), .Y(n4868) );
  OAI221XL U16438 ( .A0(n2578), .A1(n11349), .B0(n1610), .B1(n25), .C0(n11350), 
        .Y(n11343) );
  OAI221XL U16439 ( .A0(n2594), .A1(n11346), .B0(n2590), .B1(n11347), .C0(
        n11348), .Y(n11344) );
  AOI221X1 U16440 ( .A0(n10467), .A1(n2732), .B0(n2734), .B1(n10468), .C0(
        n5176), .Y(n10466) );
  INVX1 U16441 ( .A(n10469), .Y(n5176) );
  OAI221XL U16442 ( .A0(n2760), .A1(n10473), .B0(n1613), .B1(n26), .C0(n10474), 
        .Y(n10467) );
  OAI221XL U16443 ( .A0(n2774), .A1(n10470), .B0(n2772), .B1(n10471), .C0(
        n10472), .Y(n10468) );
  AOI221X1 U16444 ( .A0(n9591), .A1(n2914), .B0(n2916), .B1(n9592), .C0(n5422), 
        .Y(n9590) );
  INVX1 U16445 ( .A(n9593), .Y(n5422) );
  OAI221XL U16446 ( .A0(n2942), .A1(n9597), .B0(n1616), .B1(n27), .C0(n9598), 
        .Y(n9591) );
  OAI221XL U16447 ( .A0(n2959), .A1(n9594), .B0(n2954), .B1(n9595), .C0(n9596), 
        .Y(n9592) );
  AOI221X1 U16448 ( .A0(n8715), .A1(n3094), .B0(n3096), .B1(n8716), .C0(n5650), 
        .Y(n8714) );
  INVX1 U16449 ( .A(n8717), .Y(n5650) );
  OAI221XL U16450 ( .A0(n3122), .A1(n8721), .B0(n1619), .B1(n28), .C0(n8722), 
        .Y(n8715) );
  OAI221XL U16451 ( .A0(n3141), .A1(n8718), .B0(n3134), .B1(n8719), .C0(n8720), 
        .Y(n8716) );
  AOI221X1 U16452 ( .A0(n7839), .A1(n3274), .B0(n3276), .B1(n7840), .C0(n5886), 
        .Y(n7838) );
  INVX1 U16453 ( .A(n7841), .Y(n5886) );
  OAI221XL U16454 ( .A0(n3302), .A1(n7845), .B0(n1622), .B1(n29), .C0(n7846), 
        .Y(n7839) );
  OAI221XL U16455 ( .A0(n3321), .A1(n7842), .B0(n3314), .B1(n7843), .C0(n7844), 
        .Y(n7840) );
  AOI222X1 U16456 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n320), .A1(n3454), 
        .B0(n3455), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n321), .C0(n1139), 
        .C1(n6119), .Y(top_core_EC_ss_gen_tbox_0__sboxs_r_n306) );
  NAND3X1 U16457 ( .A(top_core_EC_ss_gen_tbox_0__sboxs_r_n323), .B(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n274), .C(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n324), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n320) );
  OAI221XL U16458 ( .A0(n530), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n102), 
        .B0(n1625), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n218), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n322), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n321) );
  AOI222X1 U16459 ( .A0(n10134), .A1(n2853), .B0(n2863), .B1(n10135), .C0(n996), .C1(n5333), .Y(n10120) );
  NAND3X1 U16460 ( .A(n10137), .B(n10088), .C(n10138), .Y(n10134) );
  OAI221XL U16461 ( .A0(n529), .A1(n9918), .B0(n1615), .B1(n10032), .C0(n10136), .Y(n10135) );
  AOI222X1 U16462 ( .A0(n11302), .A1(n2611), .B0(n2621), .B1(n11303), .C0(n940), .C1(n4979), .Y(n11288) );
  NAND3X1 U16463 ( .A(n11305), .B(n11256), .C(n11306), .Y(n11302) );
  OAI221XL U16464 ( .A0(n531), .A1(n11086), .B0(n1611), .B1(n11200), .C0(
        n11304), .Y(n11303) );
  AOI222X1 U16465 ( .A0(n8382), .A1(n3213), .B0(n3223), .B1(n8383), .C0(n1080), 
        .C1(n5805), .Y(n8368) );
  NAND3X1 U16466 ( .A(n8385), .B(n8336), .C(n8386), .Y(n8382) );
  OAI221XL U16467 ( .A0(n532), .A1(n8166), .B0(n1621), .B1(n8280), .C0(n8384), 
        .Y(n8383) );
  AOI222X1 U16468 ( .A0(n11010), .A1(n2672), .B0(n2682), .B1(n11011), .C0(n954), .C1(n5063), .Y(n10996) );
  NAND3X1 U16469 ( .A(n11013), .B(n10964), .C(n11014), .Y(n11010) );
  OAI221XL U16470 ( .A0(n533), .A1(n10794), .B0(n1612), .B1(n10908), .C0(
        n11012), .Y(n11011) );
  AOI222X1 U16471 ( .A0(n9258), .A1(n3033), .B0(n3043), .B1(n9259), .C0(n1038), 
        .C1(n5569), .Y(n9244) );
  NAND3X1 U16472 ( .A(n9261), .B(n9212), .C(n9262), .Y(n9258) );
  OAI221XL U16473 ( .A0(n534), .A1(n9042), .B0(n1618), .B1(n9156), .C0(n9260), 
        .Y(n9259) );
  AOI222X1 U16474 ( .A0(n7506), .A1(n3393), .B0(n3403), .B1(n7507), .C0(n1122), 
        .C1(n6033), .Y(n7492) );
  NAND3X1 U16475 ( .A(n7509), .B(n7460), .C(n7510), .Y(n7506) );
  OAI221XL U16476 ( .A0(n535), .A1(n7290), .B0(n1624), .B1(n7404), .C0(n7508), 
        .Y(n7507) );
  AOI222X1 U16477 ( .A0(n10426), .A1(n2793), .B0(n2803), .B1(n10427), .C0(n982), .C1(n5249), .Y(n10412) );
  NAND3X1 U16478 ( .A(n10429), .B(n10380), .C(n10430), .Y(n10426) );
  OAI221XL U16479 ( .A0(n536), .A1(n10210), .B0(n1614), .B1(n10324), .C0(
        n10428), .Y(n10427) );
  AOI222X1 U16480 ( .A0(n9550), .A1(n2975), .B0(n2985), .B1(n9551), .C0(n1024), 
        .C1(n5493), .Y(n9536) );
  NAND3X1 U16481 ( .A(n9553), .B(n9504), .C(n9554), .Y(n9550) );
  OAI221XL U16482 ( .A0(n537), .A1(n9334), .B0(n1617), .B1(n9448), .C0(n9552), 
        .Y(n9551) );
  AOI222X1 U16483 ( .A0(n8674), .A1(n3152), .B0(n3162), .B1(n8675), .C0(n1066), 
        .C1(n5721), .Y(n8660) );
  NAND3X1 U16484 ( .A(n8677), .B(n8628), .C(n8678), .Y(n8674) );
  OAI221XL U16485 ( .A0(n538), .A1(n8458), .B0(n1620), .B1(n8572), .C0(n8676), 
        .Y(n8675) );
  AOI222X1 U16486 ( .A0(n7798), .A1(n3335), .B0(n3345), .B1(n7799), .C0(n1108), 
        .C1(n5957), .Y(n7784) );
  NAND3X1 U16487 ( .A(n7801), .B(n7752), .C(n7802), .Y(n7798) );
  OAI221XL U16488 ( .A0(n539), .A1(n7582), .B0(n1623), .B1(n7696), .C0(n7800), 
        .Y(n7799) );
  AOI222X1 U16489 ( .A0(n11594), .A1(n2550), .B0(n2560), .B1(n11595), .C0(n926), .C1(n4863), .Y(n11580) );
  NAND3X1 U16490 ( .A(n11597), .B(n11548), .C(n11598), .Y(n11594) );
  OAI221XL U16491 ( .A0(n540), .A1(n11378), .B0(n1610), .B1(n11492), .C0(
        n11596), .Y(n11595) );
  AOI222X1 U16492 ( .A0(n10718), .A1(n2732), .B0(n2742), .B1(n10719), .C0(n968), .C1(n5171), .Y(n10704) );
  NAND3X1 U16493 ( .A(n10721), .B(n10672), .C(n10722), .Y(n10718) );
  OAI221XL U16494 ( .A0(n541), .A1(n10502), .B0(n1613), .B1(n10616), .C0(
        n10720), .Y(n10719) );
  AOI222X1 U16495 ( .A0(n9842), .A1(n2914), .B0(n2924), .B1(n9843), .C0(n1010), 
        .C1(n5417), .Y(n9828) );
  NAND3X1 U16496 ( .A(n9845), .B(n9796), .C(n9846), .Y(n9842) );
  OAI221XL U16497 ( .A0(n542), .A1(n9626), .B0(n1616), .B1(n9740), .C0(n9844), 
        .Y(n9843) );
  AOI222X1 U16498 ( .A0(n8966), .A1(n3094), .B0(n3104), .B1(n8967), .C0(n1052), 
        .C1(n5645), .Y(n8952) );
  NAND3X1 U16499 ( .A(n8969), .B(n8920), .C(n8970), .Y(n8966) );
  OAI221XL U16500 ( .A0(n543), .A1(n8750), .B0(n1619), .B1(n8864), .C0(n8968), 
        .Y(n8967) );
  AOI222X1 U16501 ( .A0(n8090), .A1(n3274), .B0(n3284), .B1(n8091), .C0(n1094), 
        .C1(n5881), .Y(n8076) );
  NAND3X1 U16502 ( .A(n8093), .B(n8044), .C(n8094), .Y(n8090) );
  OAI221XL U16503 ( .A0(n544), .A1(n7874), .B0(n1622), .B1(n7988), .C0(n8092), 
        .Y(n8091) );
  INVX1 U16504 ( .A(n11799), .Y(n6912) );
  INVX1 U16505 ( .A(top_core_KE_sb1_n227), .Y(n6866) );
  INVX1 U16506 ( .A(n12430), .Y(n6619) );
  INVX1 U16507 ( .A(n12115), .Y(n6572) );
  AOI222X1 U16508 ( .A0(n2854), .A1(n17283), .B0(n17284), .B1(n2851), .C0(
        n5328), .C1(n2887), .Y(n17282) );
  NAND4X1 U16509 ( .A(n17114), .B(n17073), .C(n17286), .D(n17287), .Y(n17283)
         );
  OAI211XL U16510 ( .A0(n17285), .A1(n17072), .B0(n17036), .C0(n17026), .Y(
        n17284) );
  AOI222X1 U16511 ( .A0(n5363), .A1(top_core_EC_ss_in[80]), .B0(n17175), .B1(
        n417), .C0(n5380), .C1(n386), .Y(n17287) );
  AOI222X1 U16512 ( .A0(n3463), .A1(n14133), .B0(n14134), .B1(n3452), .C0(
        n6112), .C1(n3487), .Y(n14132) );
  NAND4X1 U16513 ( .A(n13964), .B(n13923), .C(n14136), .D(n14137), .Y(n14133)
         );
  OAI211XL U16514 ( .A0(n14135), .A1(n13922), .B0(n13886), .C0(n13876), .Y(
        n14134) );
  AOI222X1 U16515 ( .A0(n6131), .A1(n3503), .B0(n14025), .B1(n418), .C0(n6151), 
        .C1(n385), .Y(n14137) );
  AOI222X1 U16516 ( .A0(n3214), .A1(n15393), .B0(n15394), .B1(n3211), .C0(
        n5800), .C1(n3250), .Y(n15392) );
  NAND4X1 U16517 ( .A(n15224), .B(n15183), .C(n15396), .D(n15397), .Y(n15393)
         );
  OAI211XL U16518 ( .A0(n15395), .A1(n15182), .B0(n15146), .C0(n15136), .Y(
        n15394) );
  AOI222X1 U16519 ( .A0(n5835), .A1(top_core_EC_ss_in[32]), .B0(n15285), .B1(
        n420), .C0(n5852), .C1(n388), .Y(n15397) );
  AOI222X1 U16520 ( .A0(n2620), .A1(n18543), .B0(n18544), .B1(n2622), .C0(
        n4974), .C1(n2642), .Y(n18542) );
  NAND4X1 U16521 ( .A(n18374), .B(n18333), .C(n18546), .D(n18547), .Y(n18543)
         );
  OAI211XL U16522 ( .A0(n18545), .A1(n18332), .B0(n18296), .C0(n18286), .Y(
        n18544) );
  AOI222X1 U16523 ( .A0(n5009), .A1(n2651), .B0(n18435), .B1(n419), .C0(n5026), 
        .C1(n387), .Y(n18547) );
  AOI222X1 U16524 ( .A0(n3161), .A1(n15708), .B0(n15709), .B1(n3150), .C0(
        n5716), .C1(n3184), .Y(n15707) );
  NAND4X1 U16525 ( .A(n15539), .B(n15498), .C(n15711), .D(n15712), .Y(n15708)
         );
  OAI211XL U16526 ( .A0(n15710), .A1(n15497), .B0(n15461), .C0(n15451), .Y(
        n15709) );
  AOI222X1 U16527 ( .A0(n5751), .A1(top_core_EC_ss_in[40]), .B0(n15600), .B1(
        n426), .C0(n5768), .C1(n389), .Y(n15712) );
  AOI222X1 U16528 ( .A0(n2923), .A1(n16968), .B0(n16969), .B1(n2912), .C0(
        n5412), .C1(n2946), .Y(n16967) );
  NAND4X1 U16529 ( .A(n16799), .B(n16758), .C(n16971), .D(n16972), .Y(n16968)
         );
  OAI211XL U16530 ( .A0(n16970), .A1(n16757), .B0(n16721), .C0(n16711), .Y(
        n16969) );
  AOI222X1 U16531 ( .A0(n5447), .A1(top_core_EC_ss_in[72]), .B0(n16860), .B1(
        n430), .C0(n5464), .C1(n391), .Y(n16972) );
  AOI222X1 U16532 ( .A0(n2558), .A1(n18858), .B0(n18859), .B1(n2548), .C0(
        n4858), .C1(n2582), .Y(n18857) );
  NAND4X1 U16533 ( .A(n18689), .B(n18648), .C(n18861), .D(n18862), .Y(n18858)
         );
  OAI211XL U16534 ( .A0(n18860), .A1(n18647), .B0(n18611), .C0(n18601), .Y(
        n18859) );
  AOI222X1 U16535 ( .A0(n4893), .A1(n2590), .B0(n18750), .B1(n428), .C0(n4910), 
        .C1(n390), .Y(n18862) );
  AOI222X1 U16536 ( .A0(n3283), .A1(n15078), .B0(n15079), .B1(n3272), .C0(
        n5876), .C1(n3311), .Y(n15077) );
  NAND4X1 U16537 ( .A(n14909), .B(n14868), .C(n15081), .D(n15082), .Y(n15078)
         );
  OAI211XL U16538 ( .A0(n15080), .A1(n14867), .B0(n14831), .C0(n14821), .Y(
        n15079) );
  AOI222X1 U16539 ( .A0(n5911), .A1(n3325), .B0(n14970), .B1(n432), .C0(n5928), 
        .C1(n392), .Y(n15082) );
  AOI222X1 U16540 ( .A0(n2984), .A1(n16653), .B0(n16654), .B1(n2973), .C0(
        n5488), .C1(n3012), .Y(n16652) );
  NAND4X1 U16541 ( .A(n16484), .B(n16443), .C(n16656), .D(n16657), .Y(n16653)
         );
  OAI211XL U16542 ( .A0(n16655), .A1(n16442), .B0(n16406), .C0(n16396), .Y(
        n16654) );
  AOI222X1 U16543 ( .A0(n5523), .A1(n3016), .B0(n16545), .B1(n425), .C0(n5540), 
        .C1(n393), .Y(n16657) );
  AOI222X1 U16544 ( .A0(n2673), .A1(n18228), .B0(n18229), .B1(n2670), .C0(
        n5058), .C1(n2704), .Y(n18227) );
  NAND4X1 U16545 ( .A(n18059), .B(n18018), .C(n18231), .D(n18232), .Y(n18228)
         );
  OAI211XL U16546 ( .A0(n18230), .A1(n18017), .B0(n17981), .C0(n17971), .Y(
        n18229) );
  AOI222X1 U16547 ( .A0(n5093), .A1(top_core_EC_ss_in[104]), .B0(n18120), .B1(
        n421), .C0(n5110), .C1(n394), .Y(n18232) );
  AOI222X1 U16548 ( .A0(n3344), .A1(n14763), .B0(n14764), .B1(n3346), .C0(
        n5952), .C1(n3367), .Y(n14762) );
  NAND4X1 U16549 ( .A(n14594), .B(n14553), .C(n14766), .D(n14767), .Y(n14763)
         );
  OAI211XL U16550 ( .A0(n14765), .A1(n14552), .B0(n14516), .C0(n14506), .Y(
        n14764) );
  AOI222X1 U16551 ( .A0(n5987), .A1(n3376), .B0(n14655), .B1(n427), .C0(n6004), 
        .C1(n395), .Y(n14767) );
  AOI222X1 U16552 ( .A0(n3042), .A1(n16338), .B0(n16339), .B1(n3044), .C0(
        n5564), .C1(n3065), .Y(n16337) );
  NAND4X1 U16553 ( .A(n16169), .B(n16128), .C(n16341), .D(n16342), .Y(n16338)
         );
  OAI211XL U16554 ( .A0(n16340), .A1(n16127), .B0(n16091), .C0(n16081), .Y(
        n16339) );
  AOI222X1 U16555 ( .A0(n5599), .A1(n3073), .B0(n16230), .B1(n422), .C0(n5616), 
        .C1(n396), .Y(n16342) );
  AOI222X1 U16556 ( .A0(n2733), .A1(n17913), .B0(n17914), .B1(n2730), .C0(
        n5166), .C1(n2764), .Y(n17912) );
  NAND4X1 U16557 ( .A(n17744), .B(n17703), .C(n17916), .D(n17917), .Y(n17913)
         );
  OAI211XL U16558 ( .A0(n17915), .A1(n17702), .B0(n17666), .C0(n17656), .Y(
        n17914) );
  AOI222X1 U16559 ( .A0(n5201), .A1(n2773), .B0(n17805), .B1(n429), .C0(n5218), 
        .C1(n397), .Y(n17917) );
  AOI222X1 U16560 ( .A0(n3402), .A1(n14448), .B0(n14449), .B1(n3404), .C0(
        n6028), .C1(n3424), .Y(n14447) );
  NAND4X1 U16561 ( .A(n14279), .B(n14238), .C(n14451), .D(n14452), .Y(n14448)
         );
  OAI211XL U16562 ( .A0(n14450), .A1(n14237), .B0(n14201), .C0(n14191), .Y(
        n14449) );
  AOI222X1 U16563 ( .A0(n6063), .A1(top_core_EC_ss_in[8]), .B0(n14340), .B1(
        n423), .C0(n6080), .C1(n398), .Y(n14452) );
  AOI222X1 U16564 ( .A0(n3095), .A1(n16023), .B0(n16024), .B1(n3092), .C0(
        n5640), .C1(n3126), .Y(n16022) );
  NAND4X1 U16565 ( .A(n15854), .B(n15813), .C(n16026), .D(n16027), .Y(n16023)
         );
  OAI211XL U16566 ( .A0(n16025), .A1(n15812), .B0(n15776), .C0(n15766), .Y(
        n16024) );
  AOI222X1 U16567 ( .A0(n5675), .A1(n3135), .B0(n15915), .B1(n431), .C0(n5692), 
        .C1(n399), .Y(n16027) );
  AOI222X1 U16568 ( .A0(n2802), .A1(n17598), .B0(n17599), .B1(n2791), .C0(
        n5244), .C1(n2825), .Y(n17597) );
  NAND4X1 U16569 ( .A(n17429), .B(n17388), .C(n17601), .D(n17602), .Y(n17598)
         );
  OAI211XL U16570 ( .A0(n17600), .A1(n17387), .B0(n17351), .C0(n17341), .Y(
        n17599) );
  AOI222X1 U16571 ( .A0(n5279), .A1(n2834), .B0(n17490), .B1(n424), .C0(n5296), 
        .C1(n400), .Y(n17602) );
  OAI21XL U16572 ( .A0(n9970), .A1(n9912), .B0(n9886), .Y(n10106) );
  OAI21XL U16573 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n156), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n96), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n68), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n292) );
  OAI21XL U16574 ( .A0(n8218), .A1(n8160), .B0(n8134), .Y(n8354) );
  OAI21XL U16575 ( .A0(n11138), .A1(n11080), .B0(n11054), .Y(n11274) );
  OAI21XL U16576 ( .A0(n10846), .A1(n10788), .B0(n10762), .Y(n10982) );
  OAI21XL U16577 ( .A0(n7342), .A1(n7284), .B0(n7258), .Y(n7478) );
  OAI21XL U16578 ( .A0(n9094), .A1(n9036), .B0(n9010), .Y(n9230) );
  OAI21XL U16579 ( .A0(n10262), .A1(n10204), .B0(n10178), .Y(n10398) );
  OAI21XL U16580 ( .A0(n9386), .A1(n9328), .B0(n9302), .Y(n9522) );
  OAI21XL U16581 ( .A0(n8510), .A1(n8452), .B0(n8426), .Y(n8646) );
  OAI21XL U16582 ( .A0(n7634), .A1(n7576), .B0(n7550), .Y(n7770) );
  OAI21XL U16583 ( .A0(n11430), .A1(n11372), .B0(n11346), .Y(n11566) );
  OAI21XL U16584 ( .A0(n10554), .A1(n10496), .B0(n10470), .Y(n10690) );
  OAI21XL U16585 ( .A0(n9678), .A1(n9620), .B0(n9594), .Y(n9814) );
  OAI21XL U16586 ( .A0(n8802), .A1(n8744), .B0(n8718), .Y(n8938) );
  OAI21XL U16587 ( .A0(n7926), .A1(n7868), .B0(n7842), .Y(n8062) );
  AOI21X1 U16588 ( .A0(n9919), .A1(n9914), .B0(n2899), .Y(n9987) );
  AOI21X1 U16589 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n104), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n98), .B0(n3506), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n173) );
  AOI21X1 U16590 ( .A0(n11087), .A1(n11082), .B0(n2656), .Y(n11155) );
  AOI21X1 U16591 ( .A0(n8167), .A1(n8162), .B0(n3259), .Y(n8235) );
  AOI21X1 U16592 ( .A0(n10795), .A1(n10790), .B0(n2717), .Y(n10863) );
  AOI21X1 U16593 ( .A0(n9043), .A1(n9038), .B0(n3078), .Y(n9111) );
  AOI21X1 U16594 ( .A0(n7291), .A1(n7286), .B0(n3439), .Y(n7359) );
  AOI21X1 U16595 ( .A0(n10211), .A1(n10206), .B0(n2842), .Y(n10279) );
  AOI21X1 U16596 ( .A0(n9335), .A1(n9330), .B0(n3023), .Y(n9403) );
  AOI21X1 U16597 ( .A0(n8459), .A1(n8454), .B0(n3198), .Y(n8527) );
  AOI21X1 U16598 ( .A0(n7583), .A1(n7578), .B0(n3383), .Y(n7651) );
  AOI21X1 U16599 ( .A0(n11379), .A1(n11374), .B0(n2595), .Y(n11447) );
  AOI21X1 U16600 ( .A0(n10503), .A1(n10498), .B0(n2780), .Y(n10571) );
  AOI21X1 U16601 ( .A0(n9627), .A1(n9622), .B0(n2960), .Y(n9695) );
  AOI21X1 U16602 ( .A0(n8751), .A1(n8746), .B0(n3142), .Y(n8819) );
  AOI21X1 U16603 ( .A0(n7875), .A1(n7870), .B0(n3322), .Y(n7943) );
  AND2X2 U16604 ( .A(n1806), .B(n1815), .Y(n673) );
  AND2X2 U16605 ( .A(n1827), .B(n1836), .Y(n674) );
  AND2X2 U16606 ( .A(n1762), .B(n1770), .Y(n675) );
  AND2X2 U16607 ( .A(n1785), .B(n1794), .Y(n676) );
  AND2X2 U16608 ( .A(n1685), .B(n1689), .Y(n677) );
  AND2X2 U16609 ( .A(n1743), .B(n1747), .Y(n678) );
  AND2X2 U16610 ( .A(n1654), .B(n1660), .Y(n679) );
  AND2X2 U16611 ( .A(n1714), .B(n1718), .Y(n680) );
  AOI222X1 U16612 ( .A0(n2906), .A1(n5353), .B0(n417), .B1(n17153), .C0(n633), 
        .C1(n465), .Y(n17151) );
  AOI222X1 U16613 ( .A0(n3504), .A1(n6121), .B0(n418), .B1(n14003), .C0(n634), 
        .C1(n466), .Y(n14001) );
  AOI222X1 U16614 ( .A0(n2651), .A1(n4999), .B0(n419), .B1(n18413), .C0(n635), 
        .C1(n467), .Y(n18411) );
  AOI222X1 U16615 ( .A0(n3266), .A1(n5825), .B0(n420), .B1(n15263), .C0(n636), 
        .C1(n468), .Y(n15261) );
  AOI222X1 U16616 ( .A0(n3205), .A1(n5741), .B0(n426), .B1(n15578), .C0(n637), 
        .C1(n469), .Y(n15576) );
  AOI222X1 U16617 ( .A0(n2590), .A1(n4883), .B0(n428), .B1(n18728), .C0(n638), 
        .C1(n471), .Y(n18726) );
  AOI222X1 U16618 ( .A0(n2967), .A1(n5437), .B0(n430), .B1(n16838), .C0(n639), 
        .C1(n470), .Y(n16836) );
  AOI222X1 U16619 ( .A0(top_core_EC_ss_in[24]), .A1(n5901), .B0(n432), .B1(
        n14948), .C0(n640), .C1(n472), .Y(n14946) );
  AOI222X1 U16620 ( .A0(n3016), .A1(n5513), .B0(n425), .B1(n16523), .C0(n641), 
        .C1(n473), .Y(n16521) );
  AOI222X1 U16621 ( .A0(n2721), .A1(n5083), .B0(n421), .B1(n18098), .C0(n642), 
        .C1(n474), .Y(n18096) );
  AOI222X1 U16622 ( .A0(n3376), .A1(n5977), .B0(n427), .B1(n14633), .C0(n643), 
        .C1(n475), .Y(n14631) );
  AOI222X1 U16623 ( .A0(n3073), .A1(n5589), .B0(n422), .B1(n16208), .C0(n644), 
        .C1(n476), .Y(n16206) );
  AOI222X1 U16624 ( .A0(n2773), .A1(n5191), .B0(n429), .B1(n17783), .C0(n645), 
        .C1(n477), .Y(n17781) );
  AOI222X1 U16625 ( .A0(n3443), .A1(n6053), .B0(n423), .B1(n14318), .C0(n646), 
        .C1(n478), .Y(n14316) );
  AOI222X1 U16626 ( .A0(n3135), .A1(n5665), .B0(n431), .B1(n15893), .C0(n647), 
        .C1(n479), .Y(n15891) );
  AOI222X1 U16627 ( .A0(n2834), .A1(n5269), .B0(n424), .B1(n17468), .C0(n648), 
        .C1(n480), .Y(n17466) );
  CLKINVX3 U16628 ( .A(n2262), .Y(n2261) );
  AND2X2 U16629 ( .A(n1802), .B(n1813), .Y(n681) );
  AND2X2 U16630 ( .A(n1823), .B(n1834), .Y(n682) );
  AND2X2 U16631 ( .A(n1760), .B(n1773), .Y(n683) );
  AND2X2 U16632 ( .A(n1781), .B(n1792), .Y(n684) );
  AND2X2 U16633 ( .A(n1651), .B(n1661), .Y(n685) );
  AND2X2 U16634 ( .A(n1680), .B(n1691), .Y(n686) );
  AND2X2 U16635 ( .A(n1709), .B(n1720), .Y(n687) );
  AND2X2 U16636 ( .A(n1738), .B(n1749), .Y(n688) );
  AND2X2 U16637 ( .A(n1804), .B(n1811), .Y(n689) );
  AND2X2 U16638 ( .A(n1825), .B(n1832), .Y(n690) );
  AND2X2 U16639 ( .A(n1762), .B(n1772), .Y(n691) );
  AND2X2 U16640 ( .A(n1686), .B(n1693), .Y(n692) );
  AND2X2 U16641 ( .A(n1783), .B(n1790), .Y(n693) );
  AND2X2 U16642 ( .A(n1744), .B(n1751), .Y(n694) );
  AND2X2 U16643 ( .A(n1654), .B(n1660), .Y(n695) );
  AND2X2 U16644 ( .A(n1715), .B(n1722), .Y(n696) );
  INVX1 U16645 ( .A(top_core_KE_n1359), .Y(n6336) );
  INVX1 U16646 ( .A(n17201), .Y(n5324) );
  AOI22X1 U16647 ( .A0(n5325), .A1(n17202), .B0(n5326), .B1(n17203), .Y(n17201) );
  NAND4XL U16648 ( .A(n17163), .B(n17075), .C(n17081), .D(n17204), .Y(n17203)
         );
  NAND4BXL U16649 ( .AN(n17206), .B(n17027), .C(n17143), .D(n17207), .Y(n17202) );
  INVX1 U16650 ( .A(n14051), .Y(n6106) );
  AOI22X1 U16651 ( .A0(n6107), .A1(n14052), .B0(n6108), .B1(n14053), .Y(n14051) );
  NAND4XL U16652 ( .A(n14013), .B(n13925), .C(n13931), .D(n14054), .Y(n14053)
         );
  NAND4BXL U16653 ( .AN(n14056), .B(n13877), .C(n13993), .D(n14057), .Y(n14052) );
  INVX1 U16654 ( .A(n18461), .Y(n4970) );
  AOI22X1 U16655 ( .A0(n4971), .A1(n18462), .B0(n4972), .B1(n18463), .Y(n18461) );
  NAND4XL U16656 ( .A(n18423), .B(n18335), .C(n18341), .D(n18464), .Y(n18463)
         );
  NAND4BXL U16657 ( .AN(n18466), .B(n18287), .C(n18403), .D(n18467), .Y(n18462) );
  INVX1 U16658 ( .A(n15311), .Y(n5796) );
  AOI22X1 U16659 ( .A0(n5797), .A1(n15312), .B0(n5798), .B1(n15313), .Y(n15311) );
  NAND4XL U16660 ( .A(n15273), .B(n15185), .C(n15191), .D(n15314), .Y(n15313)
         );
  NAND4BXL U16661 ( .AN(n15316), .B(n15137), .C(n15253), .D(n15317), .Y(n15312) );
  INVX1 U16662 ( .A(n15626), .Y(n5712) );
  AOI22X1 U16663 ( .A0(n5713), .A1(n15627), .B0(n5714), .B1(n15628), .Y(n15626) );
  NAND4XL U16664 ( .A(n15588), .B(n15500), .C(n15506), .D(n15629), .Y(n15628)
         );
  NAND4BXL U16665 ( .AN(n15631), .B(n15452), .C(n15568), .D(n15632), .Y(n15627) );
  INVX1 U16666 ( .A(n16886), .Y(n5408) );
  AOI22X1 U16667 ( .A0(n5409), .A1(n16887), .B0(n5410), .B1(n16888), .Y(n16886) );
  NAND4XL U16668 ( .A(n16848), .B(n16760), .C(n16766), .D(n16889), .Y(n16888)
         );
  NAND4BXL U16669 ( .AN(n16891), .B(n16712), .C(n16828), .D(n16892), .Y(n16887) );
  INVX1 U16670 ( .A(n18776), .Y(n4854) );
  AOI22X1 U16671 ( .A0(n4855), .A1(n18777), .B0(n4856), .B1(n18778), .Y(n18776) );
  NAND4XL U16672 ( .A(n18738), .B(n18650), .C(n18656), .D(n18779), .Y(n18778)
         );
  NAND4BXL U16673 ( .AN(n18781), .B(n18602), .C(n18718), .D(n18782), .Y(n18777) );
  INVX1 U16674 ( .A(n14996), .Y(n5872) );
  AOI22X1 U16675 ( .A0(n5873), .A1(n14997), .B0(n5874), .B1(n14998), .Y(n14996) );
  NAND4XL U16676 ( .A(n14958), .B(n14870), .C(n14876), .D(n14999), .Y(n14998)
         );
  NAND4BXL U16677 ( .AN(n15001), .B(n14822), .C(n14938), .D(n15002), .Y(n14997) );
  INVX1 U16678 ( .A(n16571), .Y(n5484) );
  AOI22X1 U16679 ( .A0(n5485), .A1(n16572), .B0(n5486), .B1(n16573), .Y(n16571) );
  NAND4XL U16680 ( .A(n16533), .B(n16445), .C(n16451), .D(n16574), .Y(n16573)
         );
  NAND4BXL U16681 ( .AN(n16576), .B(n16397), .C(n16513), .D(n16577), .Y(n16572) );
  INVX1 U16682 ( .A(n18146), .Y(n5054) );
  AOI22X1 U16683 ( .A0(n5055), .A1(n18147), .B0(n5056), .B1(n18148), .Y(n18146) );
  NAND4XL U16684 ( .A(n18108), .B(n18020), .C(n18026), .D(n18149), .Y(n18148)
         );
  NAND4BXL U16685 ( .AN(n18151), .B(n17972), .C(n18088), .D(n18152), .Y(n18147) );
  INVX1 U16686 ( .A(n14681), .Y(n5948) );
  AOI22X1 U16687 ( .A0(n5949), .A1(n14682), .B0(n5950), .B1(n14683), .Y(n14681) );
  NAND4XL U16688 ( .A(n14643), .B(n14555), .C(n14561), .D(n14684), .Y(n14683)
         );
  NAND4BXL U16689 ( .AN(n14686), .B(n14507), .C(n14623), .D(n14687), .Y(n14682) );
  INVX1 U16690 ( .A(n16256), .Y(n5560) );
  AOI22X1 U16691 ( .A0(n5561), .A1(n16257), .B0(n5562), .B1(n16258), .Y(n16256) );
  NAND4XL U16692 ( .A(n16218), .B(n16130), .C(n16136), .D(n16259), .Y(n16258)
         );
  NAND4BXL U16693 ( .AN(n16261), .B(n16082), .C(n16198), .D(n16262), .Y(n16257) );
  INVX1 U16694 ( .A(n17831), .Y(n5162) );
  AOI22X1 U16695 ( .A0(n5163), .A1(n17832), .B0(n5164), .B1(n17833), .Y(n17831) );
  NAND4XL U16696 ( .A(n17793), .B(n17705), .C(n17711), .D(n17834), .Y(n17833)
         );
  NAND4BXL U16697 ( .AN(n17836), .B(n17657), .C(n17773), .D(n17837), .Y(n17832) );
  INVX1 U16698 ( .A(n14366), .Y(n6024) );
  AOI22X1 U16699 ( .A0(n6025), .A1(n14367), .B0(n6026), .B1(n14368), .Y(n14366) );
  NAND4XL U16700 ( .A(n14328), .B(n14240), .C(n14246), .D(n14369), .Y(n14368)
         );
  NAND4BXL U16701 ( .AN(n14371), .B(n14192), .C(n14308), .D(n14372), .Y(n14367) );
  INVX1 U16702 ( .A(n15941), .Y(n5636) );
  AOI22X1 U16703 ( .A0(n5637), .A1(n15942), .B0(n5638), .B1(n15943), .Y(n15941) );
  NAND4XL U16704 ( .A(n15903), .B(n15815), .C(n15821), .D(n15944), .Y(n15943)
         );
  NAND4BXL U16705 ( .AN(n15946), .B(n15767), .C(n15883), .D(n15947), .Y(n15942) );
  INVX1 U16706 ( .A(n17516), .Y(n5240) );
  AOI22X1 U16707 ( .A0(n5241), .A1(n17517), .B0(n5242), .B1(n17518), .Y(n17516) );
  NAND4XL U16708 ( .A(n17478), .B(n17390), .C(n17396), .D(n17519), .Y(n17518)
         );
  NAND4BXL U16709 ( .AN(n17521), .B(n17342), .C(n17458), .D(n17522), .Y(n17517) );
  INVX1 U16710 ( .A(n3960), .Y(n3907) );
  INVX1 U16711 ( .A(n3938), .Y(n3960) );
  INVX1 U16712 ( .A(n3906), .Y(n3947) );
  INVX1 U16713 ( .A(n2286), .Y(n2304) );
  INVX1 U16714 ( .A(n2286), .Y(n2303) );
  INVX1 U16715 ( .A(n2286), .Y(n2302) );
  INVX1 U16716 ( .A(n3231), .Y(n3233) );
  INVX1 U16717 ( .A(n3170), .Y(n3172) );
  INVX1 U16718 ( .A(n3353), .Y(n3355) );
  INVX1 U16719 ( .A(n2750), .Y(n2752) );
  INVX1 U16720 ( .A(top_core_EC_ss_in[2]), .Y(n3480) );
  INVX1 U16721 ( .A(top_core_EC_ss_in[82]), .Y(n2879) );
  INVX1 U16722 ( .A(n237), .Y(n3627) );
  INVX1 U16723 ( .A(top_core_EC_ss_in[114]), .Y(n2637) );
  INVX1 U16724 ( .A(top_core_EC_ss_in[34]), .Y(n3239) );
  INVX1 U16725 ( .A(top_core_EC_ss_in[42]), .Y(n3178) );
  INVX1 U16726 ( .A(top_core_EC_ss_in[122]), .Y(n2576) );
  INVX1 U16727 ( .A(top_core_EC_ss_in[74]), .Y(n2940) );
  INVX1 U16728 ( .A(top_core_EC_ss_in[66]), .Y(n3001) );
  INVX1 U16729 ( .A(top_core_EC_ss_in[106]), .Y(n2698) );
  INVX1 U16730 ( .A(top_core_EC_ss_in[18]), .Y(n3361) );
  INVX1 U16731 ( .A(top_core_EC_ss_in[58]), .Y(n3059) );
  INVX1 U16732 ( .A(top_core_EC_ss_in[98]), .Y(n2758) );
  INVX1 U16733 ( .A(top_core_EC_ss_in[10]), .Y(n3419) );
  INVX1 U16734 ( .A(top_core_EC_ss_in[50]), .Y(n3120) );
  INVX1 U16735 ( .A(top_core_EC_ss_in[26]), .Y(n3300) );
  INVX1 U16736 ( .A(top_core_EC_ss_in[90]), .Y(n2819) );
  INVX1 U16737 ( .A(n2220), .Y(n2235) );
  INVX1 U16738 ( .A(n2525), .Y(n2521) );
  INVX1 U16739 ( .A(n4089), .Y(n4104) );
  INVX1 U16740 ( .A(n4115), .Y(n4097) );
  INVX1 U16741 ( .A(n4112), .Y(n4105) );
  INVX1 U16742 ( .A(n4113), .Y(n4102) );
  INVX1 U16743 ( .A(n4111), .Y(n4107) );
  INVX1 U16744 ( .A(n4074), .Y(n4099) );
  INVX1 U16745 ( .A(n4072), .Y(n4100) );
  INVX1 U16746 ( .A(n4066), .Y(n4101) );
  INVX1 U16747 ( .A(n4115), .Y(n4096) );
  INVX1 U16748 ( .A(n4112), .Y(n4106) );
  INVX1 U16749 ( .A(n4114), .Y(n4098) );
  INVX1 U16750 ( .A(n4113), .Y(n4103) );
  INVX1 U16751 ( .A(n4094), .Y(n4108) );
  INVX1 U16752 ( .A(n4085), .Y(n4109) );
  INVX1 U16753 ( .A(n3653), .Y(n3679) );
  INVX1 U16754 ( .A(n3686), .Y(n3680) );
  INVX1 U16755 ( .A(n3686), .Y(n3681) );
  INVX1 U16756 ( .A(n3644), .Y(n3682) );
  INVX1 U16757 ( .A(n3644), .Y(n3683) );
  INVX1 U16758 ( .A(n3644), .Y(n3684) );
  INVX1 U16759 ( .A(n3686), .Y(n3685) );
  INVX1 U16760 ( .A(n3962), .Y(n3956) );
  INVX1 U16761 ( .A(n3928), .Y(n3954) );
  INVX1 U16762 ( .A(n3962), .Y(n3955) );
  INVX1 U16763 ( .A(n3913), .Y(n3957) );
  INVX1 U16764 ( .A(n3961), .Y(n3958) );
  INVX1 U16765 ( .A(n3961), .Y(n3959) );
  INVX1 U16766 ( .A(n3910), .Y(n3948) );
  INVX1 U16767 ( .A(n3913), .Y(n3952) );
  INVX1 U16768 ( .A(n3962), .Y(n3949) );
  INVX1 U16769 ( .A(n3918), .Y(n3950) );
  INVX1 U16770 ( .A(n3907), .Y(n3951) );
  INVX1 U16771 ( .A(n3962), .Y(n3953) );
  INVX1 U16772 ( .A(n4025), .Y(n4029) );
  INVX1 U16773 ( .A(n2542), .Y(n2536) );
  INVX1 U16774 ( .A(n2542), .Y(n2537) );
  INVX1 U16775 ( .A(n2542), .Y(n2535) );
  INVX1 U16776 ( .A(n2216), .Y(n2204) );
  INVX1 U16778 ( .A(n2284), .Y(n2305) );
  INVX1 U16779 ( .A(n4026), .Y(n4030) );
  INVX1 U16780 ( .A(n2289), .Y(n2291) );
  INVX1 U16781 ( .A(top_core_KE_n1876), .Y(n2272) );
  INVX1 U16782 ( .A(n2286), .Y(n2292) );
  INVX1 U16783 ( .A(top_core_EC_n870), .Y(n3553) );
  INVX1 U16784 ( .A(n2538), .Y(n2525) );
  INVX1 U16785 ( .A(n2391), .Y(n2523) );
  INVX1 U16786 ( .A(n2385), .Y(n2522) );
  INVX1 U16787 ( .A(n2538), .Y(n2524) );
  INVX1 U16788 ( .A(top_core_EC_ss_in[0]), .Y(n3506) );
  INVX1 U16789 ( .A(top_core_EC_ss_in[80]), .Y(n2904) );
  INVX1 U16790 ( .A(top_core_EC_ss_in[112]), .Y(n2662) );
  INVX1 U16791 ( .A(top_core_EC_ss_in[32]), .Y(n3264) );
  INVX1 U16792 ( .A(top_core_EC_ss_in[81]), .Y(n2890) );
  INVX1 U16793 ( .A(top_core_EC_ss_in[1]), .Y(n3491) );
  INVX1 U16794 ( .A(n2906), .Y(n2905) );
  INVX1 U16795 ( .A(top_core_EC_ss_in[33]), .Y(n3250) );
  INVX1 U16796 ( .A(top_core_EC_ss_in[113]), .Y(n2648) );
  INVX1 U16797 ( .A(n2661), .Y(n2663) );
  INVX1 U16798 ( .A(n3266), .Y(n3265) );
  INVX1 U16799 ( .A(top_core_EC_ss_in[40]), .Y(n3203) );
  INVX1 U16800 ( .A(top_core_EC_ss_in[120]), .Y(n2601) );
  INVX1 U16801 ( .A(top_core_EC_ss_in[72]), .Y(n2965) );
  INVX1 U16802 ( .A(top_core_Addr[3]), .Y(n3974) );
  INVX1 U16803 ( .A(top_core_EC_ss_in[64]), .Y(n3024) );
  INVX1 U16804 ( .A(top_core_EC_ss_in[16]), .Y(n3384) );
  INVX1 U16805 ( .A(top_core_EC_ss_in[48]), .Y(n3143) );
  INVX1 U16806 ( .A(top_core_EC_ss_in[88]), .Y(n2845) );
  INVX1 U16807 ( .A(n3205), .Y(n3204) );
  INVX1 U16808 ( .A(n2724), .Y(n2723) );
  INVX1 U16809 ( .A(top_core_EC_ss_in[104]), .Y(n2722) );
  INVX1 U16810 ( .A(top_core_EC_ss_in[105]), .Y(n2709) );
  INVX1 U16811 ( .A(top_core_EC_ss_in[56]), .Y(n3084) );
  INVX1 U16812 ( .A(n3083), .Y(n3085) );
  INVX1 U16813 ( .A(n2967), .Y(n2966) );
  INVX1 U16814 ( .A(top_core_EC_ss_in[8]), .Y(n3444) );
  INVX1 U16815 ( .A(n3446), .Y(n3445) );
  INVX1 U16816 ( .A(top_core_EC_ss_in[57]), .Y(n3070) );
  INVX1 U16817 ( .A(n2600), .Y(n2602) );
  INVX1 U16818 ( .A(top_core_EC_ss_in[9]), .Y(n3430) );
  INVX1 U16819 ( .A(top_core_EC_ss_in[89]), .Y(n2830) );
  INVX1 U16820 ( .A(top_core_EC_ss_in[65]), .Y(n3012) );
  INVX1 U16821 ( .A(top_core_EC_ss_in[17]), .Y(n3373) );
  INVX1 U16822 ( .A(top_core_EC_ss_in[97]), .Y(n2770) );
  INVX1 U16823 ( .A(top_core_Addr[2]), .Y(n3987) );
  INVX1 U16824 ( .A(top_core_EC_ss_in[49]), .Y(n3132) );
  INVX1 U16825 ( .A(top_core_EC_ss_in[25]), .Y(n3311) );
  INVX1 U16826 ( .A(n3984), .Y(n3986) );
  INVX1 U16827 ( .A(n3970), .Y(n3973) );
  INVX1 U16828 ( .A(top_core_EC_ss_in[41]), .Y(n3190) );
  INVX1 U16829 ( .A(top_core_EC_ss_in[121]), .Y(n2588) );
  INVX1 U16830 ( .A(top_core_EC_ss_in[73]), .Y(n2951) );
  INVX1 U16831 ( .A(n2539), .Y(n2534) );
  INVX1 U16832 ( .A(top_core_KE_n874), .Y(n1896) );
  INVX1 U16833 ( .A(top_core_KE_n877), .Y(n1936) );
  INVX1 U16834 ( .A(top_core_KE_n880), .Y(n1976) );
  INVX1 U16835 ( .A(top_core_KE_n886), .Y(n2056) );
  INVX1 U16836 ( .A(top_core_KE_n889), .Y(n2096) );
  INVX1 U16837 ( .A(top_core_KE_n891), .Y(n2136) );
  INVX1 U16838 ( .A(n1880), .Y(n1893) );
  INVX1 U16839 ( .A(n1920), .Y(n1933) );
  INVX1 U16840 ( .A(n1960), .Y(n1973) );
  INVX1 U16841 ( .A(n2040), .Y(n2053) );
  INVX1 U16842 ( .A(n2079), .Y(n2093) );
  INVX1 U16843 ( .A(n2119), .Y(n2133) );
  INVX1 U16844 ( .A(n1878), .Y(n1895) );
  INVX1 U16845 ( .A(n1918), .Y(n1935) );
  INVX1 U16846 ( .A(n1958), .Y(n1975) );
  INVX1 U16847 ( .A(n2038), .Y(n2055) );
  INVX1 U16848 ( .A(n2087), .Y(n2095) );
  INVX1 U16849 ( .A(n2117), .Y(n2135) );
  INVX1 U16850 ( .A(top_core_KE_n874), .Y(n1894) );
  INVX1 U16851 ( .A(top_core_KE_n877), .Y(n1934) );
  INVX1 U16852 ( .A(top_core_KE_n880), .Y(n1974) );
  INVX1 U16853 ( .A(top_core_KE_n886), .Y(n2054) );
  INVX1 U16854 ( .A(top_core_KE_n889), .Y(n2094) );
  INVX1 U16855 ( .A(top_core_KE_n891), .Y(n2134) );
  INVX1 U16856 ( .A(top_core_KE_n882), .Y(n2016) );
  INVX1 U16857 ( .A(n1999), .Y(n2013) );
  INVX1 U16858 ( .A(n1997), .Y(n2015) );
  INVX1 U16859 ( .A(top_core_KE_n882), .Y(n2014) );
  INVX1 U16860 ( .A(top_core_EC_n730), .Y(n3524) );
  INVX1 U16861 ( .A(n4257), .Y(n1605) );
  INVX1 U16862 ( .A(n4257), .Y(n1606) );
  INVX1 U16863 ( .A(n4257), .Y(n1607) );
  INVX1 U16864 ( .A(n4257), .Y(n1608) );
  INVX1 U16865 ( .A(top_core_Addr[1]), .Y(n4028) );
  INVX1 U16866 ( .A(top_core_Addr[3]), .Y(n3975) );
  INVX1 U16867 ( .A(top_core_EC_ss_in[4]), .Y(n3471) );
  INVX1 U16868 ( .A(top_core_EC_ss_in[84]), .Y(n2870) );
  INVX1 U16869 ( .A(top_core_EC_ss_in[116]), .Y(n2628) );
  INVX1 U16870 ( .A(top_core_EC_ss_in[36]), .Y(n3230) );
  INVX1 U16871 ( .A(top_core_EC_ss_in[44]), .Y(n3169) );
  INVX1 U16872 ( .A(top_core_EC_ss_in[124]), .Y(n2567) );
  INVX1 U16873 ( .A(top_core_EC_ss_in[76]), .Y(n2931) );
  INVX1 U16874 ( .A(top_core_EC_ss_in[28]), .Y(n3291) );
  INVX1 U16875 ( .A(top_core_EC_ss_in[68]), .Y(n2992) );
  INVX1 U16876 ( .A(top_core_EC_ss_in[108]), .Y(n2689) );
  INVX1 U16877 ( .A(top_core_EC_ss_in[20]), .Y(n3352) );
  INVX1 U16878 ( .A(top_core_EC_ss_in[60]), .Y(n3050) );
  INVX1 U16879 ( .A(top_core_EC_ss_in[12]), .Y(n3410) );
  INVX1 U16880 ( .A(top_core_EC_ss_in[52]), .Y(n3111) );
  INVX1 U16881 ( .A(top_core_EC_ss_in[92]), .Y(n2810) );
  NOR2X2 U16882 ( .A(n4127), .B(n4128), .Y(top_core_io_n177) );
  NOR2X1 U16883 ( .A(n4136), .B(n4124), .Y(top_core_io_n166) );
  AND2X2 U16884 ( .A(top_core_io_n621), .B(top_core_io_n188), .Y(
        top_core_io_n528) );
  AND2X2 U16885 ( .A(top_core_io_n621), .B(top_core_io_n177), .Y(
        top_core_io_n517) );
  AND2X2 U16886 ( .A(top_core_io_n621), .B(top_core_io_n166), .Y(
        top_core_io_n506) );
  AND2X2 U16887 ( .A(top_core_io_n621), .B(top_core_io_n155), .Y(
        top_core_io_n495) );
  AND2X2 U16888 ( .A(top_core_io_n324), .B(top_core_io_n177), .Y(
        top_core_io_n222) );
  AND2X2 U16889 ( .A(top_core_io_n324), .B(top_core_io_n188), .Y(
        top_core_io_n233) );
  AND2X2 U16890 ( .A(top_core_io_n324), .B(top_core_io_n166), .Y(
        top_core_io_n211) );
  AND2X2 U16891 ( .A(top_core_io_n324), .B(top_core_io_n155), .Y(
        top_core_io_n200) );
  AND2X2 U16892 ( .A(top_core_io_n154), .B(top_core_io_n177), .Y(
        top_core_io_n49) );
  AND2X2 U16893 ( .A(top_core_io_n188), .B(top_core_io_n154), .Y(
        top_core_io_n60) );
  AND2X2 U16894 ( .A(top_core_io_n166), .B(top_core_io_n154), .Y(
        top_core_io_n38) );
  AND2X2 U16895 ( .A(top_core_io_n154), .B(top_core_io_n155), .Y(
        top_core_io_n27) );
  CLKINVX3 U16896 ( .A(n4125), .Y(n4119) );
  CLKINVX3 U16897 ( .A(n4125), .Y(n4117) );
  CLKINVX3 U16898 ( .A(n4125), .Y(n4118) );
  CLKINVX3 U16899 ( .A(n4137), .Y(n4128) );
  CLKINVX3 U16900 ( .A(n4126), .Y(n4124) );
  NOR2X1 U16901 ( .A(n4136), .B(n4126), .Y(top_core_io_n155) );
  CLKINVX3 U16902 ( .A(n4127), .Y(n4122) );
  CLKINVX3 U16903 ( .A(n4125), .Y(n4123) );
  CLKINVX3 U16904 ( .A(n4125), .Y(n4121) );
  CLKINVX3 U16905 ( .A(n4127), .Y(n4120) );
  CLKINVX3 U16906 ( .A(n4127), .Y(n4116) );
  CLKINVX3 U16907 ( .A(n4143), .Y(n4141) );
  CLKINVX3 U16908 ( .A(n4137), .Y(n4129) );
  CLKINVX3 U16909 ( .A(n4136), .Y(n4130) );
  CLKINVX3 U16910 ( .A(n4137), .Y(n4135) );
  CLKINVX3 U16911 ( .A(n4136), .Y(n4133) );
  CLKINVX3 U16912 ( .A(n4136), .Y(n4134) );
  CLKINVX3 U16913 ( .A(n4137), .Y(n4132) );
  CLKINVX3 U16914 ( .A(n4137), .Y(n4131) );
  CLKINVX3 U16915 ( .A(n4140), .Y(n4139) );
  CLKINVX3 U16916 ( .A(n_DIN[7]), .Y(n1557) );
  CLKINVX3 U16917 ( .A(n_DIN[6]), .Y(n1560) );
  CLKINVX3 U16918 ( .A(n_DIN[5]), .Y(n1563) );
  CLKINVX3 U16919 ( .A(n_DIN[4]), .Y(n1566) );
  CLKINVX3 U16920 ( .A(n_DIN[3]), .Y(n1569) );
  CLKINVX3 U16921 ( .A(n_DIN[7]), .Y(n1558) );
  CLKINVX3 U16922 ( .A(n_DIN[6]), .Y(n1561) );
  CLKINVX3 U16923 ( .A(n_DIN[5]), .Y(n1564) );
  CLKINVX3 U16924 ( .A(n_DIN[4]), .Y(n1567) );
  CLKINVX3 U16925 ( .A(n_DIN[3]), .Y(n1570) );
  CLKINVX3 U16926 ( .A(n_DIN[2]), .Y(n1573) );
  CLKINVX3 U16927 ( .A(n_DIN[1]), .Y(n1576) );
  CLKINVX3 U16928 ( .A(n_DIN[7]), .Y(n1559) );
  CLKINVX3 U16929 ( .A(n_DIN[6]), .Y(n1562) );
  CLKINVX3 U16930 ( .A(n_DIN[5]), .Y(n1565) );
  CLKINVX3 U16931 ( .A(n_DIN[4]), .Y(n1568) );
  CLKINVX3 U16932 ( .A(n_DIN[3]), .Y(n1571) );
  CLKINVX3 U16933 ( .A(n_DIN[2]), .Y(n1574) );
  CLKINVX3 U16934 ( .A(n_DIN[1]), .Y(n1577) );
  OAI22X2 U16935 ( .A0(n2486), .A1(top_core_EC_ss_n156), .B0(n2373), .B1(n155), 
        .Y(top_core_EC_mc_mix_in_8[79]) );
  OAI22X2 U16936 ( .A0(n2534), .A1(top_core_EC_ss_n248), .B0(n2367), .B1(n161), 
        .Y(top_core_EC_mc_mix_in_8[111]) );
  OAI22X2 U16937 ( .A0(n2440), .A1(top_core_EC_ss_n161), .B0(n2373), .B1(n153), 
        .Y(top_core_EC_mc_mix_in_2_64_) );
  OAI22X2 U16938 ( .A0(n2469), .A1(top_core_EC_ss_n253), .B0(n2367), .B1(n159), 
        .Y(top_core_EC_mc_mix_in_2_96_) );
  OAI22X2 U16939 ( .A0(n2523), .A1(top_core_EC_ss_n142), .B0(n2374), .B1(n157), 
        .Y(top_core_EC_mc_mix_in_2_90_) );
  OAI22X2 U16940 ( .A0(n2526), .A1(top_core_EC_ss_n233), .B0(n2537), .B1(n163), 
        .Y(top_core_EC_mc_mix_in_2_122_) );
  NOR2X2 U16941 ( .A(n6964), .B(n1797), .Y(n11652) );
  NOR2X2 U16942 ( .A(n6958), .B(n1818), .Y(top_core_KE_sb1_n77) );
  NOR2X2 U16943 ( .A(n1171), .B(top_core_KE_prev_key1_reg_29_), .Y(n12284) );
  NOR2X2 U16944 ( .A(n6670), .B(n1776), .Y(n11968) );
  NOR2X2 U16945 ( .A(n1643), .B(n1640), .Y(n13544) );
  OAI22X2 U16946 ( .A0(n2440), .A1(top_core_EC_ss_n159), .B0(n2373), .B1(n154), 
        .Y(top_core_EC_mc_mix_in_2_74_) );
  OAI22X2 U16947 ( .A0(n2475), .A1(top_core_EC_ss_n251), .B0(n2367), .B1(n160), 
        .Y(top_core_EC_mc_mix_in_2_106_) );
  AOI32X1 U16948 ( .A0(top_core_EC_n1022), .A1(n3975), .A2(n3986), .B0(n2511), 
        .B1(n6306), .Y(top_core_EC_n1024) );
  OAI22X2 U16949 ( .A0(n2447), .A1(top_core_EC_ss_n147), .B0(n2374), .B1(n156), 
        .Y(top_core_EC_mc_mix_in_8[87]) );
  OAI22X2 U16950 ( .A0(n2428), .A1(top_core_EC_ss_n239), .B0(n2538), .B1(n162), 
        .Y(top_core_EC_mc_mix_in_8[119]) );
  OAI22X2 U16951 ( .A0(n2438), .A1(top_core_EC_ss_n165), .B0(n2372), .B1(n152), 
        .Y(top_core_EC_mc_mix_in_8[71]) );
  OAI22X2 U16952 ( .A0(n2445), .A1(top_core_EC_ss_n256), .B0(n2367), .B1(n158), 
        .Y(top_core_EC_mc_mix_in_8[103]) );
  NAND2X2 U16953 ( .A(top_core_EC_ss_in[2]), .B(n1517), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n104) );
  NAND2X2 U16954 ( .A(n2878), .B(n1505), .Y(n9919) );
  NAND2X2 U16955 ( .A(n2636), .B(n1529), .Y(n11087) );
  NAND2X2 U16956 ( .A(n3236), .B(n1519), .Y(n8167) );
  NAND2X2 U16957 ( .A(n2696), .B(n1531), .Y(n10795) );
  NAND2X2 U16958 ( .A(n3417), .B(n1527), .Y(n7291) );
  NAND2X2 U16959 ( .A(n3058), .B(n1512), .Y(n9043) );
  NAND2X2 U16960 ( .A(n2813), .B(n1503), .Y(n10211) );
  NAND2X2 U16961 ( .A(n2999), .B(n1510), .Y(n9335) );
  NAND2X2 U16962 ( .A(n3175), .B(n1516), .Y(n8459) );
  NAND2X2 U16963 ( .A(n3358), .B(n1523), .Y(n7583) );
  NAND2X2 U16964 ( .A(n2575), .B(n1526), .Y(n11379) );
  NAND2X2 U16965 ( .A(n2755), .B(n1501), .Y(n10503) );
  NAND2X2 U16966 ( .A(n2938), .B(n1508), .Y(n9627) );
  NAND2X2 U16967 ( .A(n3119), .B(n1514), .Y(n8751) );
  NAND2X2 U16968 ( .A(n3294), .B(n1521), .Y(n7875) );
  NAND2X2 U16969 ( .A(n6598), .B(n1648), .Y(n13608) );
  NAND2X2 U16970 ( .A(n2866), .B(n1505), .Y(n9886) );
  NAND2X2 U16971 ( .A(n3467), .B(n1517), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n68) );
  NAND2X2 U16972 ( .A(n2624), .B(n1529), .Y(n11054) );
  NAND2X2 U16973 ( .A(n3226), .B(n1519), .Y(n8134) );
  NAND2X2 U16974 ( .A(n2685), .B(n1531), .Y(n10762) );
  NAND2X2 U16975 ( .A(n3046), .B(n1512), .Y(n9010) );
  NAND2X2 U16976 ( .A(n3406), .B(n1527), .Y(n7258) );
  NAND2X2 U16977 ( .A(n2806), .B(n1503), .Y(n10178) );
  NAND2X2 U16978 ( .A(n2988), .B(n1510), .Y(n9302) );
  NAND2X2 U16979 ( .A(n3165), .B(n1516), .Y(n8426) );
  NAND2X2 U16980 ( .A(n3348), .B(n1523), .Y(n7550) );
  NAND2X2 U16981 ( .A(n2563), .B(n1526), .Y(n11346) );
  NAND2X2 U16982 ( .A(n2745), .B(n1501), .Y(n10470) );
  NAND2X2 U16983 ( .A(n2927), .B(n1508), .Y(n9594) );
  NAND2X2 U16984 ( .A(n3107), .B(n1514), .Y(n8718) );
  NAND2X2 U16985 ( .A(n3287), .B(n1521), .Y(n7842) );
  NOR2X2 U16986 ( .A(n11797), .B(n11811), .Y(n11849) );
  NOR2X2 U16987 ( .A(top_core_KE_sb1_n225), .B(top_core_KE_sb1_n239), .Y(
        top_core_KE_sb1_n278) );
  NOR2X2 U16988 ( .A(n12428), .B(n12442), .Y(n12480) );
  NOR2X2 U16989 ( .A(n13373), .B(n13387), .Y(n13425) );
  NOR2X2 U16990 ( .A(n12113), .B(n12127), .Y(n12165) );
  NOR2X2 U16991 ( .A(n12743), .B(n12757), .Y(n12795) );
  NOR2X2 U16992 ( .A(n13688), .B(n13702), .Y(n13740) );
  NOR2X2 U16993 ( .A(n13058), .B(n13072), .Y(n13110) );
  NOR2X2 U16994 ( .A(n2871), .B(n1505), .Y(n17153) );
  NOR2X2 U16995 ( .A(n3472), .B(n1517), .Y(n14003) );
  NOR2X2 U16996 ( .A(n2629), .B(n1529), .Y(n18413) );
  NOR2X2 U16997 ( .A(n3231), .B(n1519), .Y(n15263) );
  NOR2X2 U16998 ( .A(n3170), .B(n1516), .Y(n15578) );
  NOR2X2 U16999 ( .A(n2932), .B(n1508), .Y(n16838) );
  NOR2X2 U17000 ( .A(n2568), .B(n1526), .Y(n18728) );
  NOR2X2 U17001 ( .A(n3292), .B(n1521), .Y(n14948) );
  NOR2X2 U17002 ( .A(n2993), .B(n1510), .Y(n16523) );
  NOR2X2 U17003 ( .A(n2690), .B(n1531), .Y(n18098) );
  NOR2X2 U17004 ( .A(n3353), .B(n1523), .Y(n14633) );
  NOR2X2 U17005 ( .A(n3051), .B(n1512), .Y(n16208) );
  NOR2X2 U17006 ( .A(n2750), .B(n1501), .Y(n17783) );
  NOR2X2 U17007 ( .A(n3411), .B(n1527), .Y(n14318) );
  NOR2X2 U17008 ( .A(n3112), .B(n1514), .Y(n15893) );
  NOR2X2 U17009 ( .A(n2811), .B(n1503), .Y(n17468) );
  NAND2X2 U17010 ( .A(top_core_KE_prev_key1_reg_13_), .B(n1211), .Y(n11679) );
  NAND2X2 U17011 ( .A(top_core_KE_prev_key1_reg_5_), .B(n1210), .Y(
        top_core_KE_sb1_n104) );
  NAND2X2 U17012 ( .A(n1757), .B(n1171), .Y(n12310) );
  NAND2X2 U17013 ( .A(top_core_KE_prev_key1_reg_21_), .B(n1170), .Y(n11995) );
  NAND2X2 U17014 ( .A(top_core_KE_prev_key1_reg_93_), .B(n1643), .Y(n13571) );
  NAND2X2 U17015 ( .A(n1505), .B(n2870), .Y(n9918) );
  NAND2X2 U17016 ( .A(n1517), .B(n3469), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n102) );
  NAND2X2 U17017 ( .A(n1529), .B(n2628), .Y(n11086) );
  NAND2X2 U17018 ( .A(n1519), .B(n3230), .Y(n8166) );
  NAND2X2 U17019 ( .A(n1531), .B(n2689), .Y(n10794) );
  NAND2X2 U17020 ( .A(n1512), .B(n3048), .Y(n9042) );
  NAND2X2 U17021 ( .A(n1527), .B(n3408), .Y(n7290) );
  NAND2X2 U17022 ( .A(n1503), .B(n2810), .Y(n10210) );
  NAND2X2 U17023 ( .A(n1510), .B(n2992), .Y(n9334) );
  NAND2X2 U17024 ( .A(n1516), .B(n3169), .Y(n8458) );
  NAND2X2 U17025 ( .A(n1523), .B(n3352), .Y(n7582) );
  NAND2X2 U17026 ( .A(n1526), .B(n2567), .Y(n11378) );
  NAND2X2 U17027 ( .A(n1501), .B(n2749), .Y(n10502) );
  NAND2X2 U17028 ( .A(n1508), .B(n2931), .Y(n9626) );
  NAND2X2 U17029 ( .A(n1514), .B(n3111), .Y(n8750) );
  NAND2X2 U17030 ( .A(n1521), .B(n3291), .Y(n7874) );
  NAND2X2 U17031 ( .A(n1163), .B(n1171), .Y(n12483) );
  NAND2X2 U17032 ( .A(n1171), .B(n1752), .Y(n12305) );
  NOR2X1 U17033 ( .A(n11718), .B(n11679), .Y(n11712) );
  NOR2X1 U17034 ( .A(top_core_KE_sb1_n145), .B(top_core_KE_sb1_n104), .Y(
        top_core_KE_sb1_n138) );
  NOR2X1 U17035 ( .A(n12349), .B(n12310), .Y(n12343) );
  NOR2X1 U17036 ( .A(n13295), .B(n13256), .Y(n13289) );
  NOR2X1 U17037 ( .A(n12034), .B(n11995), .Y(n12028) );
  NOR2X1 U17038 ( .A(n12980), .B(n12941), .Y(n12974) );
  NOR2X1 U17039 ( .A(n13610), .B(n13571), .Y(n13604) );
  NOR2X1 U17040 ( .A(n12665), .B(n12626), .Y(n12659) );
  OAI22X1 U17041 ( .A0(n2542), .A1(top_core_EC_ss_n132), .B0(n2375), .B1(n219), 
        .Y(top_core_EC_mix_in[98]) );
  OAI22X1 U17042 ( .A0(n2527), .A1(top_core_EC_ss_n134), .B0(n2374), .B1(n217), 
        .Y(top_core_EC_mix_in[96]) );
  OAI22X1 U17043 ( .A0(n2493), .A1(top_core_EC_ss_n131), .B0(n2375), .B1(n220), 
        .Y(top_core_EC_mix_in[99]) );
  AOI22X1 U17044 ( .A0(n1643), .A1(n1660), .B0(n1645), .B1(n631), .Y(n13609)
         );
  OAI22X1 U17045 ( .A0(n2440), .A1(top_core_EC_ss_n160), .B0(n2373), .B1(n201), 
        .Y(top_core_EC_mix_in[72]) );
  OAI22X1 U17046 ( .A0(n2429), .A1(top_core_EC_ss_n158), .B0(n2373), .B1(n202), 
        .Y(top_core_EC_mix_in[74]) );
  OAI22X1 U17047 ( .A0(n2485), .A1(top_core_EC_ss_n157), .B0(n2373), .B1(n203), 
        .Y(top_core_EC_mix_in[75]) );
  OAI22X1 U17048 ( .A0(n2468), .A1(top_core_EC_ss_n149), .B0(n2373), .B1(n209), 
        .Y(top_core_EC_mix_in[82]) );
  OAI22X1 U17049 ( .A0(n2440), .A1(top_core_EC_ss_n151), .B0(n2373), .B1(n207), 
        .Y(top_core_EC_mix_in[80]) );
  OAI22X1 U17050 ( .A0(n2476), .A1(top_core_EC_ss_n148), .B0(n2373), .B1(n210), 
        .Y(top_core_EC_mix_in[83]) );
  OAI22X1 U17051 ( .A0(n2438), .A1(top_core_EC_ss_n167), .B0(n2372), .B1(n199), 
        .Y(top_core_EC_mix_in[66]) );
  OAI22X1 U17052 ( .A0(n2427), .A1(top_core_EC_ss_n241), .B0(n2392), .B1(n229), 
        .Y(top_core_EC_mix_in[114]) );
  OAI22X1 U17053 ( .A0(n2467), .A1(top_core_EC_ss_n169), .B0(n2372), .B1(n197), 
        .Y(top_core_EC_mix_in[64]) );
  OAI22X1 U17054 ( .A0(n2438), .A1(top_core_EC_ss_n166), .B0(n2372), .B1(n200), 
        .Y(top_core_EC_mix_in[67]) );
  OAI22X1 U17055 ( .A0(n2427), .A1(top_core_EC_ss_n243), .B0(n2512), .B1(n227), 
        .Y(top_core_EC_mix_in[112]) );
  OAI22X1 U17056 ( .A0(n2428), .A1(top_core_EC_ss_n240), .B0(n2496), .B1(n230), 
        .Y(top_core_EC_mix_in[115]) );
  OAI22X1 U17057 ( .A0(n2532), .A1(top_core_EC_ss_n252), .B0(n2367), .B1(n221), 
        .Y(top_core_EC_mix_in[104]) );
  OAI22X1 U17058 ( .A0(n2414), .A1(top_core_EC_ss_n250), .B0(n2367), .B1(n222), 
        .Y(top_core_EC_mix_in[106]) );
  OAI22X1 U17059 ( .A0(n2444), .A1(top_core_EC_ss_n249), .B0(n2367), .B1(n223), 
        .Y(top_core_EC_mix_in[107]) );
  NOR2X1 U17060 ( .A(n3476), .B(n1517), .Y(n13869) );
  NOR2X1 U17061 ( .A(n2874), .B(n1505), .Y(n17019) );
  NOR2X1 U17062 ( .A(n2632), .B(n1529), .Y(n18279) );
  NOR2X1 U17063 ( .A(n3235), .B(n1519), .Y(n15129) );
  NOR2X1 U17064 ( .A(n3174), .B(n1516), .Y(n15444) );
  NOR2X1 U17065 ( .A(n2571), .B(n1526), .Y(n18594) );
  NOR2X1 U17066 ( .A(n2935), .B(n1508), .Y(n16704) );
  NOR2X1 U17067 ( .A(n3295), .B(n1521), .Y(n14814) );
  NOR2X1 U17068 ( .A(n2996), .B(n1510), .Y(n16389) );
  NOR2X1 U17069 ( .A(n2693), .B(n1531), .Y(n17964) );
  NOR2X1 U17070 ( .A(n3357), .B(n1523), .Y(n14499) );
  NOR2X1 U17071 ( .A(n3054), .B(n1512), .Y(n16074) );
  NOR2X1 U17072 ( .A(n2754), .B(n1501), .Y(n17649) );
  NOR2X1 U17073 ( .A(n3414), .B(n1527), .Y(n14184) );
  NOR2X1 U17074 ( .A(n3115), .B(n1514), .Y(n15759) );
  NOR2X1 U17075 ( .A(n2814), .B(n1503), .Y(n17334) );
  NOR2X1 U17076 ( .A(n1166), .B(n1673), .Y(n13387) );
  NOR2X1 U17077 ( .A(n1206), .B(n1731), .Y(n12757) );
  NOR2X1 U17078 ( .A(n1208), .B(n1702), .Y(n13072) );
  NOR2X1 U17079 ( .A(n1168), .B(n1649), .Y(n13702) );
  NOR2X1 U17080 ( .A(n1211), .B(n1209), .Y(n11704) );
  NOR2X1 U17081 ( .A(n1210), .B(n1207), .Y(top_core_KE_sb1_n129) );
  NOR2X1 U17082 ( .A(n1676), .B(n1166), .Y(n13281) );
  NOR2X1 U17083 ( .A(n1170), .B(n1167), .Y(n12020) );
  NOR2X1 U17084 ( .A(n1734), .B(n1206), .Y(n12651) );
  NOR2X1 U17085 ( .A(n1643), .B(n1168), .Y(n13596) );
  NOR2X1 U17086 ( .A(n1705), .B(n1208), .Y(n12966) );
  NOR2X1 U17087 ( .A(n1171), .B(n1169), .Y(n12335) );
  NOR2X1 U17088 ( .A(n11705), .B(n77), .Y(n11681) );
  NOR2X1 U17089 ( .A(top_core_KE_sb1_n130), .B(n78), .Y(top_core_KE_sb1_n106)
         );
  NOR2X1 U17090 ( .A(n12336), .B(n184), .Y(n12312) );
  NOR2X1 U17091 ( .A(n12021), .B(n79), .Y(n11997) );
  NOR2X1 U17092 ( .A(n11779), .B(n681), .Y(n11664) );
  NOR2X1 U17093 ( .A(top_core_KE_sb1_n207), .B(n682), .Y(top_core_KE_sb1_n89)
         );
  NOR2X1 U17094 ( .A(n12410), .B(n683), .Y(n12295) );
  NOR2X1 U17095 ( .A(n12095), .B(n684), .Y(n11980) );
  NAND2X1 U17096 ( .A(n760), .B(n1171), .Y(n12337) );
  NOR2BX1 U17097 ( .AN(n11652), .B(n1209), .Y(n11827) );
  NOR2BX1 U17098 ( .AN(top_core_KE_sb1_n77), .B(n1207), .Y(
        top_core_KE_sb1_n256) );
  NOR2BX1 U17099 ( .AN(n12284), .B(n1169), .Y(n12458) );
  NOR2BX1 U17100 ( .AN(n13229), .B(n1166), .Y(n13403) );
  NOR2BX1 U17101 ( .AN(n11968), .B(n1167), .Y(n12143) );
  NOR2BX1 U17102 ( .AN(n12599), .B(n1206), .Y(n12773) );
  NOR2BX1 U17103 ( .AN(n13544), .B(n1168), .Y(n13718) );
  NOR2BX1 U17104 ( .AN(n12914), .B(n1208), .Y(n13088) );
  AND2X2 U17105 ( .A(top_core_KE_n2699), .B(top_core_KE_n896), .Y(
        top_core_KE_n1876) );
  NOR3XL U17106 ( .A(top_core_KE_n1865), .B(top_core_KE_N0), .C(
        top_core_KE_n2704), .Y(top_core_KE_n1871) );
  AOI22X1 U17107 ( .A0(top_core_EC_ss_sbox_out_r[1]), .A1(n2463), .B0(
        top_core_EC_ss_sbox_out[1]), .B1(n2390), .Y(top_core_EC_ss_n218) );
  OAI2BB2X1 U17108 ( .B0(n1506), .B1(n14093), .A0N(n1506), .A1N(n14094), .Y(
        top_core_EC_ss_sbox_out[1]) );
  OAI222XL U17109 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n305), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n276), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n306), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n278), .C0(n1506), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n307), .Y(
        top_core_EC_ss_sbox_out_r[1]) );
  AOI222X1 U17110 ( .A0(n14109), .A1(n3449), .B0(n6107), .B1(n14110), .C0(
        n6108), .C1(n14111), .Y(n14093) );
  AOI22X1 U17111 ( .A0(top_core_EC_ss_sbox_out_r[82]), .A1(n2463), .B0(
        top_core_EC_ss_sbox_out[82]), .B1(n2519), .Y(top_core_EC_ss_n220) );
  OAI222XL U17112 ( .A0(n17210), .A1(n16987), .B0(n17211), .B1(n16989), .C0(
        n1504), .C1(n17212), .Y(top_core_EC_ss_sbox_out[82]) );
  OAI222XL U17113 ( .A0(n10089), .A1(n10090), .B0(n10091), .B1(n10092), .C0(
        n1504), .C1(n10093), .Y(top_core_EC_ss_sbox_out_r[82]) );
  AOI221X1 U17114 ( .A0(n17183), .A1(n2888), .B0(n2863), .B1(n17228), .C0(
        n17229), .Y(n17211) );
  AOI22X1 U17115 ( .A0(top_core_EC_ss_sbox_out_r[2]), .A1(n2478), .B0(
        top_core_EC_ss_sbox_out[2]), .B1(n2521), .Y(top_core_EC_ss_n207) );
  OAI222XL U17116 ( .A0(n14060), .A1(n13837), .B0(n14061), .B1(n13839), .C0(
        n1506), .C1(n14062), .Y(top_core_EC_ss_sbox_out[2]) );
  OAI222XL U17117 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n275), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n276), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n277), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n278), .C0(n1506), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n279), .Y(
        top_core_EC_ss_sbox_out_r[2]) );
  AOI221X1 U17118 ( .A0(n14033), .A1(n3492), .B0(n3459), .B1(n14078), .C0(
        n14079), .Y(n14061) );
  AOI22X1 U17119 ( .A0(top_core_EC_ss_sbox_out_r[34]), .A1(n2441), .B0(
        top_core_EC_ss_sbox_out[34]), .B1(n2374), .Y(top_core_EC_ss_n202) );
  OAI222XL U17120 ( .A0(n15320), .A1(n15097), .B0(n15321), .B1(n15099), .C0(
        n1518), .C1(n15322), .Y(top_core_EC_ss_sbox_out[34]) );
  OAI222XL U17121 ( .A0(n8337), .A1(n8338), .B0(n8339), .B1(n8340), .C0(n1518), 
        .C1(n8341), .Y(top_core_EC_ss_sbox_out_r[34]) );
  AOI221X1 U17122 ( .A0(n15293), .A1(n3250), .B0(n3223), .B1(n15338), .C0(
        n15339), .Y(n15321) );
  AOI22X1 U17123 ( .A0(top_core_EC_ss_sbox_out_r[114]), .A1(n2446), .B0(
        top_core_EC_ss_sbox_out[114]), .B1(n2536), .Y(top_core_EC_ss_n184) );
  OAI222XL U17124 ( .A0(n18470), .A1(n18247), .B0(n18471), .B1(n18249), .C0(
        n1528), .C1(n18472), .Y(top_core_EC_ss_sbox_out[114]) );
  OAI222XL U17125 ( .A0(n11257), .A1(n11258), .B0(n11259), .B1(n11260), .C0(
        n1528), .C1(n11261), .Y(top_core_EC_ss_sbox_out_r[114]) );
  AOI221X1 U17126 ( .A0(n18443), .A1(n2642), .B0(n2621), .B1(n18488), .C0(
        n18489), .Y(n18471) );
  AOI22X1 U17127 ( .A0(top_core_EC_ss_sbox_out_r[80]), .A1(n2464), .B0(
        top_core_EC_ss_sbox_out[80]), .B1(n2369), .Y(top_core_EC_ss_n222) );
  OAI21XL U17128 ( .A0(n1504), .A1(n10144), .B0(n10145), .Y(
        top_core_EC_ss_sbox_out_r[80]) );
  OAI22X1 U17129 ( .A0(n17271), .A1(n992), .B0(n1504), .B1(n17272), .Y(
        top_core_EC_ss_sbox_out[80]) );
  AOI222X1 U17130 ( .A0(n2847), .A1(n10159), .B0(n9909), .B1(n10160), .C0(
        n5321), .C1(n10161), .Y(n10144) );
  AOI22X1 U17131 ( .A0(top_core_EC_ss_sbox_out_r[0]), .A1(n2476), .B0(
        top_core_EC_ss_sbox_out[0]), .B1(n2535), .Y(top_core_EC_ss_n257) );
  OAI21XL U17132 ( .A0(n1506), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n330), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n331), .Y(
        top_core_EC_ss_sbox_out_r[0]) );
  OAI22X1 U17133 ( .A0(n14121), .A1(n1132), .B0(n1506), .B1(n14122), .Y(
        top_core_EC_ss_sbox_out[0]) );
  AOI222X1 U17134 ( .A0(n3448), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n345), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n93), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n346), .C0(n6105), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n347), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n330) );
  AOI22X1 U17135 ( .A0(top_core_EC_ss_sbox_out_r[83]), .A1(n2463), .B0(
        top_core_EC_ss_sbox_out[83]), .B1(n2516), .Y(top_core_EC_ss_n219) );
  OAI21XL U17136 ( .A0(n1504), .A1(n17176), .B0(n17177), .Y(
        top_core_EC_ss_sbox_out[83]) );
  OAI22X1 U17137 ( .A0(n10056), .A1(n992), .B0(n1504), .B1(n10057), .Y(
        top_core_EC_ss_sbox_out_r[83]) );
  AOI211X1 U17138 ( .A0(n17051), .A1(n17196), .B0(n5324), .C0(n17197), .Y(
        n17176) );
  AOI22X1 U17139 ( .A0(top_core_EC_ss_sbox_out_r[7]), .A1(n2454), .B0(
        top_core_EC_ss_sbox_out[7]), .B1(n2502), .Y(top_core_EC_ss_n152) );
  OAI22X1 U17140 ( .A0(n1506), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n59), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n60), .B1(n1132), .Y(
        top_core_EC_ss_sbox_out_r[7]) );
  OAI222XL U17141 ( .A0(n13836), .A1(n13837), .B0(n13838), .B1(n13839), .C0(
        n1506), .C1(n13840), .Y(top_core_EC_ss_sbox_out[7]) );
  AOI222X1 U17142 ( .A0(n3448), .A1(top_core_EC_ss_gen_tbox_0__sboxs_r_n92), 
        .B0(top_core_EC_ss_gen_tbox_0__sboxs_r_n93), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n94), .C0(n6105), .C1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n95), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n59) );
  AOI22X1 U17143 ( .A0(top_core_EC_ss_sbox_out_r[3]), .A1(n2443), .B0(
        top_core_EC_ss_sbox_out[3]), .B1(n2367), .Y(top_core_EC_ss_n196) );
  OAI21XL U17144 ( .A0(n1506), .A1(n14026), .B0(n14027), .Y(
        top_core_EC_ss_sbox_out[3]) );
  OAI22X1 U17145 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n242), .A1(n1132), 
        .B0(n1506), .B1(top_core_EC_ss_gen_tbox_0__sboxs_r_n243), .Y(
        top_core_EC_ss_sbox_out_r[3]) );
  AOI211X1 U17146 ( .A0(n13901), .A1(n14046), .B0(n6106), .C0(n14047), .Y(
        n14026) );
  AOI22X1 U17147 ( .A0(top_core_EC_ss_sbox_out_r[32]), .A1(n2441), .B0(
        top_core_EC_ss_sbox_out[32]), .B1(n2394), .Y(top_core_EC_ss_n204) );
  OAI21XL U17148 ( .A0(n1518), .A1(n8392), .B0(n8393), .Y(
        top_core_EC_ss_sbox_out_r[32]) );
  OAI22X1 U17149 ( .A0(n15381), .A1(n1076), .B0(n1518), .B1(n15382), .Y(
        top_core_EC_ss_sbox_out[32]) );
  AOI222X1 U17150 ( .A0(n3207), .A1(n8407), .B0(n8157), .B1(n8408), .C0(n5793), 
        .C1(n8409), .Y(n8392) );
  AOI22X1 U17151 ( .A0(top_core_EC_ss_sbox_out_r[112]), .A1(n2445), .B0(
        top_core_EC_ss_sbox_out[112]), .B1(n2537), .Y(top_core_EC_ss_n187) );
  OAI21XL U17152 ( .A0(n1528), .A1(n11312), .B0(n11313), .Y(
        top_core_EC_ss_sbox_out_r[112]) );
  OAI22X1 U17153 ( .A0(n18531), .A1(n936), .B0(n1528), .B1(n18532), .Y(
        top_core_EC_ss_sbox_out[112]) );
  AOI222X1 U17154 ( .A0(n2605), .A1(n11327), .B0(n11077), .B1(n11328), .C0(
        n4967), .C1(n11329), .Y(n11312) );
  AOI22X1 U17155 ( .A0(top_core_EC_ss_sbox_out_r[115]), .A1(n2447), .B0(
        top_core_EC_ss_sbox_out[115]), .B1(n2494), .Y(top_core_EC_ss_n183) );
  OAI21XL U17156 ( .A0(n1528), .A1(n18436), .B0(n18437), .Y(
        top_core_EC_ss_sbox_out[115]) );
  OAI22X1 U17157 ( .A0(n11224), .A1(n936), .B0(n1528), .B1(n11225), .Y(
        top_core_EC_ss_sbox_out_r[115]) );
  AOI211X1 U17158 ( .A0(n18311), .A1(n18456), .B0(n4970), .C0(n18457), .Y(
        n18436) );
  AOI22X1 U17159 ( .A0(top_core_EC_ss_sbox_out_r[35]), .A1(n2442), .B0(
        top_core_EC_ss_sbox_out[35]), .B1(n2393), .Y(top_core_EC_ss_n201) );
  OAI21XL U17160 ( .A0(n1518), .A1(n15286), .B0(n15287), .Y(
        top_core_EC_ss_sbox_out[35]) );
  OAI22X1 U17161 ( .A0(n8304), .A1(n1076), .B0(n1518), .B1(n8305), .Y(
        top_core_EC_ss_sbox_out_r[35]) );
  AOI211X1 U17162 ( .A0(n15161), .A1(n15306), .B0(n5796), .C0(n15307), .Y(
        n15286) );
  AOI22X1 U17163 ( .A0(top_core_EC_ss_sbox_out_r[81]), .A1(n2464), .B0(
        top_core_EC_ss_sbox_out[81]), .B1(n2494), .Y(top_core_EC_ss_n221) );
  OAI2BB2X1 U17164 ( .B0(n1504), .B1(n17243), .A0N(n1504), .A1N(n17244), .Y(
        top_core_EC_ss_sbox_out[81]) );
  OAI222XL U17165 ( .A0(n10119), .A1(n10090), .B0(n10120), .B1(n10092), .C0(
        n1504), .C1(n10121), .Y(top_core_EC_ss_sbox_out_r[81]) );
  AOI222X1 U17166 ( .A0(n17259), .A1(n2848), .B0(n5325), .B1(n17260), .C0(
        n5326), .C1(n17261), .Y(n17243) );
  AOI22X1 U17167 ( .A0(top_core_EC_ss_sbox_out_r[106]), .A1(n2472), .B0(
        top_core_EC_ss_sbox_out[42]), .B1(n2388), .Y(top_core_EC_ss_n246) );
  OAI222XL U17168 ( .A0(n15635), .A1(n15412), .B0(n15636), .B1(n15414), .C0(
        n1515), .C1(n15637), .Y(top_core_EC_ss_sbox_out[42]) );
  OAI222XL U17169 ( .A0(n10965), .A1(n10966), .B0(n10967), .B1(n10968), .C0(
        n1530), .C1(n10969), .Y(top_core_EC_ss_sbox_out_r[106]) );
  AOI221X1 U17170 ( .A0(n15608), .A1(n3183), .B0(n3162), .B1(n15653), .C0(
        n15654), .Y(n15636) );
  AOI22X1 U17171 ( .A0(top_core_EC_ss_sbox_out_r[107]), .A1(n2468), .B0(
        top_core_EC_ss_sbox_out[43]), .B1(n2387), .Y(top_core_EC_ss_n235) );
  OAI21XL U17172 ( .A0(n1515), .A1(n15601), .B0(n15602), .Y(
        top_core_EC_ss_sbox_out[43]) );
  OAI22X1 U17173 ( .A0(n10932), .A1(n950), .B0(n1530), .B1(n10933), .Y(
        top_core_EC_ss_sbox_out_r[107]) );
  AOI211X1 U17174 ( .A0(n15476), .A1(n15621), .B0(n5712), .C0(n15622), .Y(
        n15601) );
  AOI22X1 U17175 ( .A0(top_core_EC_ss_sbox_out_r[85]), .A1(n2462), .B0(
        top_core_EC_ss_sbox_out[85]), .B1(n2515), .Y(top_core_EC_ss_n216) );
  OAI222XL U17176 ( .A0(n17102), .A1(n16989), .B0(n1504), .B1(n17103), .C0(
        n17104), .C1(n16987), .Y(top_core_EC_ss_sbox_out[85]) );
  OAI222XL U17177 ( .A0(n9977), .A1(n9932), .B0(n9978), .B1(n9934), .C0(n9979), 
        .C1(n992), .Y(top_core_EC_ss_sbox_out_r[85]) );
  AOI222X1 U17178 ( .A0(n2862), .A1(n17105), .B0(n17106), .B1(n2864), .C0(
        n5330), .C1(n17107), .Y(n17104) );
  AOI22X1 U17179 ( .A0(top_core_EC_ss_sbox_out_r[5]), .A1(n2533), .B0(
        top_core_EC_ss_sbox_out[5]), .B1(n2518), .Y(top_core_EC_ss_n174) );
  OAI222XL U17180 ( .A0(n13952), .A1(n13839), .B0(n1506), .B1(n13953), .C0(
        n13954), .C1(n13837), .Y(top_core_EC_ss_sbox_out[5]) );
  OAI222XL U17181 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n163), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n117), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n164), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n119), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n165), .C1(n1132), .Y(
        top_core_EC_ss_sbox_out_r[5]) );
  AOI222X1 U17182 ( .A0(n3458), .A1(n13955), .B0(n13956), .B1(n3465), .C0(
        n6114), .C1(n13957), .Y(n13954) );
  AOI22X1 U17183 ( .A0(top_core_EC_ss_sbox_out_r[86]), .A1(n2522), .B0(
        top_core_EC_ss_sbox_out[86]), .B1(n2517), .Y(top_core_EC_ss_n215) );
  OAI22X1 U17184 ( .A0(n1504), .A1(n17048), .B0(n17049), .B1(n992), .Y(
        top_core_EC_ss_sbox_out[86]) );
  OAI222XL U17185 ( .A0(n9931), .A1(n9932), .B0(n9933), .B1(n9934), .C0(n9935), 
        .C1(n992), .Y(top_core_EC_ss_sbox_out_r[86]) );
  AOI211X1 U17186 ( .A0(n17078), .A1(n2850), .B0(n17079), .C0(n17080), .Y(
        n17048) );
  AOI22X1 U17187 ( .A0(top_core_EC_ss_sbox_out_r[6]), .A1(n2451), .B0(
        top_core_EC_ss_sbox_out[6]), .B1(n2508), .Y(top_core_EC_ss_n163) );
  OAI22X1 U17188 ( .A0(n1506), .A1(n13898), .B0(n13899), .B1(n1132), .Y(
        top_core_EC_ss_sbox_out[6]) );
  OAI222XL U17189 ( .A0(top_core_EC_ss_gen_tbox_0__sboxs_r_n116), .A1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n117), .B0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n118), .B1(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n119), .C0(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n120), .C1(n1132), .Y(
        top_core_EC_ss_sbox_out_r[6]) );
  AOI211X1 U17190 ( .A0(n13928), .A1(n3451), .B0(n13929), .C0(n13930), .Y(
        n13898) );
  AOI22X1 U17191 ( .A0(top_core_EC_ss_sbox_out_r[87]), .A1(n2452), .B0(
        top_core_EC_ss_sbox_out[87]), .B1(n2518), .Y(top_core_EC_ss_n214) );
  OAI22X1 U17192 ( .A0(n1504), .A1(n9877), .B0(n9878), .B1(n992), .Y(
        top_core_EC_ss_sbox_out_r[87]) );
  OAI222XL U17193 ( .A0(n16986), .A1(n16987), .B0(n16988), .B1(n16989), .C0(
        n1504), .C1(n16990), .Y(top_core_EC_ss_sbox_out[87]) );
  AOI222X1 U17194 ( .A0(n2847), .A1(n9908), .B0(n9909), .B1(n9910), .C0(n5321), 
        .C1(n9911), .Y(n9877) );
  AOI22X1 U17195 ( .A0(top_core_EC_ss_sbox_out_r[113]), .A1(n2446), .B0(
        top_core_EC_ss_sbox_out[113]), .B1(n2365), .Y(top_core_EC_ss_n186) );
  OAI2BB2X1 U17196 ( .B0(n1528), .B1(n18503), .A0N(n1528), .A1N(n18504), .Y(
        top_core_EC_ss_sbox_out[113]) );
  OAI222XL U17197 ( .A0(n11287), .A1(n11258), .B0(n11288), .B1(n11260), .C0(
        n1528), .C1(n11289), .Y(top_core_EC_ss_sbox_out_r[113]) );
  AOI222X1 U17198 ( .A0(n18519), .A1(n2606), .B0(n4971), .B1(n18520), .C0(
        n4972), .C1(n18521), .Y(n18503) );
  AOI22X1 U17199 ( .A0(top_core_EC_ss_sbox_out_r[33]), .A1(n2441), .B0(
        top_core_EC_ss_sbox_out[33]), .B1(n2389), .Y(top_core_EC_ss_n203) );
  OAI2BB2X1 U17200 ( .B0(n1518), .B1(n15353), .A0N(n1518), .A1N(n15354), .Y(
        top_core_EC_ss_sbox_out[33]) );
  OAI222XL U17201 ( .A0(n8367), .A1(n8338), .B0(n8368), .B1(n8340), .C0(n1518), 
        .C1(n8369), .Y(top_core_EC_ss_sbox_out_r[33]) );
  AOI222X1 U17202 ( .A0(n15369), .A1(n3208), .B0(n5797), .B1(n15370), .C0(
        n5798), .C1(n15371), .Y(n15353) );
  AOI22X1 U17203 ( .A0(top_core_EC_ss_sbox_out_r[117]), .A1(n2447), .B0(
        top_core_EC_ss_sbox_out[117]), .B1(n2382), .Y(top_core_EC_ss_n181) );
  OAI222XL U17204 ( .A0(n18362), .A1(n18249), .B0(n1528), .B1(n18363), .C0(
        n18364), .C1(n18247), .Y(top_core_EC_ss_sbox_out[117]) );
  OAI222XL U17205 ( .A0(n11145), .A1(n11100), .B0(n11146), .B1(n11102), .C0(
        n11147), .C1(n936), .Y(top_core_EC_ss_sbox_out_r[117]) );
  AOI222X1 U17206 ( .A0(n2619), .A1(n18365), .B0(n18366), .B1(n2623), .C0(
        n4976), .C1(n18367), .Y(n18364) );
  AOI22X1 U17207 ( .A0(top_core_EC_ss_sbox_out_r[118]), .A1(n2448), .B0(
        top_core_EC_ss_sbox_out[118]), .B1(n2514), .Y(top_core_EC_ss_n180) );
  OAI22X1 U17208 ( .A0(n1528), .A1(n18308), .B0(n18309), .B1(n936), .Y(
        top_core_EC_ss_sbox_out[118]) );
  OAI222XL U17209 ( .A0(n11099), .A1(n11100), .B0(n11101), .B1(n11102), .C0(
        n11103), .C1(n936), .Y(top_core_EC_ss_sbox_out_r[118]) );
  AOI211X1 U17210 ( .A0(n18338), .A1(n2608), .B0(n18339), .C0(n18340), .Y(
        n18308) );
  AOI22X1 U17211 ( .A0(top_core_EC_ss_sbox_out_r[37]), .A1(n2442), .B0(
        top_core_EC_ss_sbox_out[37]), .B1(n2391), .Y(top_core_EC_ss_n199) );
  OAI222XL U17212 ( .A0(n15212), .A1(n15099), .B0(n1518), .B1(n15213), .C0(
        n15214), .C1(n15097), .Y(top_core_EC_ss_sbox_out[37]) );
  OAI222XL U17213 ( .A0(n8225), .A1(n8180), .B0(n8226), .B1(n8182), .C0(n8227), 
        .C1(n1076), .Y(top_core_EC_ss_sbox_out_r[37]) );
  AOI222X1 U17214 ( .A0(n3222), .A1(n15215), .B0(n15216), .B1(n3224), .C0(
        n5802), .C1(n15217), .Y(n15214) );
  AOI22X1 U17215 ( .A0(top_core_EC_ss_sbox_out_r[119]), .A1(n2448), .B0(
        top_core_EC_ss_sbox_out[119]), .B1(n2495), .Y(top_core_EC_ss_n179) );
  OAI22X1 U17216 ( .A0(n1528), .A1(n11045), .B0(n11046), .B1(n936), .Y(
        top_core_EC_ss_sbox_out_r[119]) );
  OAI222XL U17217 ( .A0(n18246), .A1(n18247), .B0(n18248), .B1(n18249), .C0(
        n1528), .C1(n18250), .Y(top_core_EC_ss_sbox_out[119]) );
  AOI222X1 U17218 ( .A0(n2605), .A1(n11076), .B0(n11077), .B1(n11078), .C0(
        n4967), .C1(n11079), .Y(n11045) );
  AOI22X1 U17219 ( .A0(top_core_EC_ss_sbox_out_r[39]), .A1(n2443), .B0(
        top_core_EC_ss_sbox_out[39]), .B1(n2385), .Y(top_core_EC_ss_n197) );
  OAI22X1 U17220 ( .A0(n1518), .A1(n8125), .B0(n8126), .B1(n1076), .Y(
        top_core_EC_ss_sbox_out_r[39]) );
  OAI222XL U17221 ( .A0(n15096), .A1(n15097), .B0(n15098), .B1(n15099), .C0(
        n1518), .C1(n15100), .Y(top_core_EC_ss_sbox_out[39]) );
  AOI222X1 U17222 ( .A0(n3207), .A1(n8156), .B0(n8157), .B1(n8158), .C0(n5793), 
        .C1(n8159), .Y(n8125) );
  AOI22X1 U17223 ( .A0(top_core_EC_ss_sbox_out_r[38]), .A1(n2443), .B0(
        top_core_EC_ss_sbox_out[38]), .B1(n2390), .Y(top_core_EC_ss_n198) );
  OAI22X1 U17224 ( .A0(n1518), .A1(n15158), .B0(n15159), .B1(n1076), .Y(
        top_core_EC_ss_sbox_out[38]) );
  OAI222XL U17225 ( .A0(n8179), .A1(n8180), .B0(n8181), .B1(n8182), .C0(n8183), 
        .C1(n1076), .Y(top_core_EC_ss_sbox_out_r[38]) );
  AOI211X1 U17226 ( .A0(n15188), .A1(n3210), .B0(n15189), .C0(n15190), .Y(
        n15158) );
  AOI22X1 U17227 ( .A0(top_core_EC_ss_sbox_out_r[111]), .A1(n2464), .B0(
        top_core_EC_ss_sbox_out[47]), .B1(n2365), .Y(top_core_EC_ss_n223) );
  OAI22X1 U17228 ( .A0(n1530), .A1(n10753), .B0(n10754), .B1(n950), .Y(
        top_core_EC_ss_sbox_out_r[111]) );
  OAI222XL U17229 ( .A0(n15411), .A1(n15412), .B0(n15413), .B1(n15414), .C0(
        n1515), .C1(n15415), .Y(top_core_EC_ss_sbox_out[47]) );
  AOI222X1 U17230 ( .A0(n2666), .A1(n10784), .B0(n10785), .B1(n10786), .C0(
        n5051), .C1(n10787), .Y(n10753) );
  AOI22X1 U17231 ( .A0(top_core_EC_ss_sbox_out_r[104]), .A1(n2458), .B0(
        top_core_EC_ss_sbox_out[40]), .B1(n2394), .Y(top_core_EC_ss_n141) );
  OAI21XL U17232 ( .A0(n1530), .A1(n11020), .B0(n11021), .Y(
        top_core_EC_ss_sbox_out_r[104]) );
  OAI22X1 U17233 ( .A0(n15696), .A1(n1062), .B0(n1515), .B1(n15697), .Y(
        top_core_EC_ss_sbox_out[40]) );
  AOI222X1 U17234 ( .A0(n2666), .A1(n11035), .B0(n10785), .B1(n11036), .C0(
        n5051), .C1(n11037), .Y(n11020) );
  AOI22X1 U17235 ( .A0(top_core_EC_ss_sbox_out_r[109]), .A1(n2465), .B0(
        top_core_EC_ss_sbox_out[45]), .B1(n2377), .Y(top_core_EC_ss_n225) );
  OAI222XL U17236 ( .A0(n15527), .A1(n15414), .B0(n1515), .B1(n15528), .C0(
        n15529), .C1(n15412), .Y(top_core_EC_ss_sbox_out[45]) );
  OAI222XL U17237 ( .A0(n10853), .A1(n10808), .B0(n10854), .B1(n10810), .C0(
        n10855), .C1(n950), .Y(top_core_EC_ss_sbox_out_r[109]) );
  AOI222X1 U17238 ( .A0(n3160), .A1(n15530), .B0(n15531), .B1(n3163), .C0(
        n5718), .C1(n15532), .Y(n15529) );
  AOI22X1 U17239 ( .A0(top_core_EC_ss_sbox_out_r[110]), .A1(n2465), .B0(
        top_core_EC_ss_sbox_out[46]), .B1(n2500), .Y(top_core_EC_ss_n224) );
  OAI22X1 U17240 ( .A0(n1515), .A1(n15473), .B0(n15474), .B1(n1062), .Y(
        top_core_EC_ss_sbox_out[46]) );
  OAI222XL U17241 ( .A0(n10807), .A1(n10808), .B0(n10809), .B1(n10810), .C0(
        n10811), .C1(n950), .Y(top_core_EC_ss_sbox_out_r[110]) );
  AOI211X1 U17242 ( .A0(n15503), .A1(n3149), .B0(n15504), .C0(n15505), .Y(
        n15473) );
  AOI22X1 U17243 ( .A0(top_core_EC_ss_sbox_out_r[63]), .A1(n2479), .B0(
        top_core_EC_ss_sbox_out[127]), .B1(n2386), .Y(top_core_EC_ss_n205) );
  OAI22X1 U17244 ( .A0(n1511), .A1(n9001), .B0(n9002), .B1(n1034), .Y(
        top_core_EC_ss_sbox_out_r[63]) );
  OAI222XL U17245 ( .A0(n18561), .A1(n18562), .B0(n18563), .B1(n18564), .C0(
        n1525), .C1(n18565), .Y(top_core_EC_ss_sbox_out[127]) );
  AOI222X1 U17246 ( .A0(n3027), .A1(n9032), .B0(n9033), .B1(n9034), .C0(n5557), 
        .C1(n9035), .Y(n9001) );
  AOI22X1 U17247 ( .A0(top_core_EC_ss_sbox_out_r[61]), .A1(n2434), .B0(
        top_core_EC_ss_sbox_out[125]), .B1(n2495), .Y(top_core_EC_ss_n208) );
  OAI222XL U17248 ( .A0(n18677), .A1(n18564), .B0(n1525), .B1(n18678), .C0(
        n18679), .C1(n18562), .Y(top_core_EC_ss_sbox_out[125]) );
  OAI222XL U17249 ( .A0(n9101), .A1(n9056), .B0(n9102), .B1(n9058), .C0(n9103), 
        .C1(n1034), .Y(top_core_EC_ss_sbox_out_r[61]) );
  AOI222X1 U17250 ( .A0(n2559), .A1(n18680), .B0(n18681), .B1(n2561), .C0(
        n4860), .C1(n18682), .Y(n18679) );
  AOI22X1 U17251 ( .A0(top_core_EC_ss_sbox_out_r[62]), .A1(n2462), .B0(
        top_core_EC_ss_sbox_out[126]), .B1(n2388), .Y(top_core_EC_ss_n206) );
  OAI22X1 U17252 ( .A0(n1525), .A1(n18623), .B0(n18624), .B1(n922), .Y(
        top_core_EC_ss_sbox_out[126]) );
  OAI222XL U17253 ( .A0(n9055), .A1(n9056), .B0(n9057), .B1(n9058), .C0(n9059), 
        .C1(n1034), .Y(top_core_EC_ss_sbox_out_r[62]) );
  AOI211X1 U17254 ( .A0(n18653), .A1(n2547), .B0(n18654), .C0(n18655), .Y(
        n18623) );
  AOI22X1 U17255 ( .A0(top_core_EC_ss_sbox_out_r[15]), .A1(n2445), .B0(
        top_core_EC_ss_sbox_out[79]), .B1(n2379), .Y(top_core_EC_ss_n188) );
  OAI22X1 U17256 ( .A0(n1524), .A1(n7249), .B0(n7250), .B1(n1118), .Y(
        top_core_EC_ss_sbox_out_r[15]) );
  OAI222XL U17257 ( .A0(n16671), .A1(n16672), .B0(n16673), .B1(n16674), .C0(
        n1507), .C1(n16675), .Y(top_core_EC_ss_sbox_out[79]) );
  AOI222X1 U17258 ( .A0(n3387), .A1(n7280), .B0(n7281), .B1(n7282), .C0(n6021), 
        .C1(n7283), .Y(n7249) );
  AOI22X1 U17259 ( .A0(top_core_EC_ss_sbox_out_r[8]), .A1(n2444), .B0(
        top_core_EC_ss_sbox_out[72]), .B1(n2387), .Y(top_core_EC_ss_n195) );
  OAI21XL U17260 ( .A0(n1524), .A1(n7516), .B0(n7517), .Y(
        top_core_EC_ss_sbox_out_r[8]) );
  OAI22X1 U17261 ( .A0(n16956), .A1(n1006), .B0(n1507), .B1(n16957), .Y(
        top_core_EC_ss_sbox_out[72]) );
  AOI222X1 U17262 ( .A0(n3387), .A1(n7531), .B0(n7281), .B1(n7532), .C0(n6021), 
        .C1(n7533), .Y(n7516) );
  AOI22X1 U17263 ( .A0(top_core_EC_ss_sbox_out_r[10]), .A1(n2444), .B0(
        top_core_EC_ss_sbox_out[74]), .B1(n2519), .Y(top_core_EC_ss_n193) );
  OAI222XL U17264 ( .A0(n16895), .A1(n16672), .B0(n16896), .B1(n16674), .C0(
        n1507), .C1(n16897), .Y(top_core_EC_ss_sbox_out[74]) );
  OAI222XL U17265 ( .A0(n7461), .A1(n7462), .B0(n7463), .B1(n7464), .C0(n1524), 
        .C1(n7465), .Y(top_core_EC_ss_sbox_out_r[10]) );
  AOI221X1 U17266 ( .A0(n16868), .A1(n2946), .B0(n2924), .B1(n16913), .C0(
        n16914), .Y(n16896) );
  AOI22X1 U17267 ( .A0(top_core_EC_ss_sbox_out_r[11]), .A1(n2523), .B0(
        top_core_EC_ss_sbox_out[75]), .B1(n2521), .Y(top_core_EC_ss_n192) );
  OAI21XL U17268 ( .A0(n1507), .A1(n16861), .B0(n16862), .Y(
        top_core_EC_ss_sbox_out[75]) );
  OAI22X1 U17269 ( .A0(n7428), .A1(n1118), .B0(n1524), .B1(n7429), .Y(
        top_core_EC_ss_sbox_out_r[11]) );
  AOI211X1 U17270 ( .A0(n16736), .A1(n16881), .B0(n5408), .C0(n16882), .Y(
        n16861) );
  AOI22X1 U17271 ( .A0(top_core_EC_ss_sbox_out_r[13]), .A1(n2430), .B0(
        top_core_EC_ss_sbox_out[77]), .B1(n2516), .Y(top_core_EC_ss_n190) );
  OAI222XL U17272 ( .A0(n16787), .A1(n16674), .B0(n1507), .B1(n16788), .C0(
        n16789), .C1(n16672), .Y(top_core_EC_ss_sbox_out[77]) );
  OAI222XL U17273 ( .A0(n7349), .A1(n7304), .B0(n7350), .B1(n7306), .C0(n7351), 
        .C1(n1118), .Y(top_core_EC_ss_sbox_out_r[13]) );
  AOI222X1 U17274 ( .A0(n2922), .A1(n16790), .B0(n16791), .B1(n2925), .C0(
        n5414), .C1(n16792), .Y(n16789) );
  AOI22X1 U17275 ( .A0(top_core_EC_ss_sbox_out_r[14]), .A1(n2445), .B0(
        top_core_EC_ss_sbox_out[78]), .B1(n2515), .Y(top_core_EC_ss_n189) );
  OAI22X1 U17276 ( .A0(n1507), .A1(n16733), .B0(n16734), .B1(n1006), .Y(
        top_core_EC_ss_sbox_out[78]) );
  OAI222XL U17277 ( .A0(n7303), .A1(n7304), .B0(n7305), .B1(n7306), .C0(n7307), 
        .C1(n1118), .Y(top_core_EC_ss_sbox_out_r[14]) );
  AOI211X1 U17278 ( .A0(n16763), .A1(n2911), .B0(n16764), .C0(n16765), .Y(
        n16733) );
  AOI22X1 U17279 ( .A0(top_core_EC_ss_sbox_out_r[56]), .A1(n2408), .B0(
        top_core_EC_ss_sbox_out[120]), .B1(n2513), .Y(top_core_EC_ss_n213) );
  OAI21XL U17280 ( .A0(n1511), .A1(n9268), .B0(n9269), .Y(
        top_core_EC_ss_sbox_out_r[56]) );
  OAI22X1 U17281 ( .A0(n18846), .A1(n922), .B0(n1525), .B1(n18847), .Y(
        top_core_EC_ss_sbox_out[120]) );
  AOI222X1 U17282 ( .A0(n3027), .A1(n9283), .B0(n9033), .B1(n9284), .C0(n5557), 
        .C1(n9285), .Y(n9268) );
  AOI22X1 U17283 ( .A0(top_core_EC_ss_sbox_out_r[58]), .A1(n2482), .B0(
        top_core_EC_ss_sbox_out[122]), .B1(n2509), .Y(top_core_EC_ss_n211) );
  OAI222XL U17284 ( .A0(n18785), .A1(n18562), .B0(n18786), .B1(n18564), .C0(
        n1525), .C1(n18787), .Y(top_core_EC_ss_sbox_out[122]) );
  OAI222XL U17285 ( .A0(n9213), .A1(n9214), .B0(n9215), .B1(n9216), .C0(n1511), 
        .C1(n9217), .Y(top_core_EC_ss_sbox_out_r[58]) );
  AOI221X1 U17286 ( .A0(n18758), .A1(n2581), .B0(n2560), .B1(n18803), .C0(
        n18804), .Y(n18786) );
  AOI22X1 U17287 ( .A0(top_core_EC_ss_sbox_out_r[59]), .A1(n2483), .B0(
        top_core_EC_ss_sbox_out[123]), .B1(n2510), .Y(top_core_EC_ss_n210) );
  OAI21XL U17288 ( .A0(n1525), .A1(n18751), .B0(n18752), .Y(
        top_core_EC_ss_sbox_out[123]) );
  OAI22X1 U17289 ( .A0(n9180), .A1(n1034), .B0(n1511), .B1(n9181), .Y(
        top_core_EC_ss_sbox_out_r[59]) );
  AOI211X1 U17290 ( .A0(n18626), .A1(n18771), .B0(n4854), .C0(n18772), .Y(
        n18751) );
  AOI22X1 U17291 ( .A0(top_core_EC_ss_sbox_out_r[105]), .A1(n2461), .B0(
        top_core_EC_ss_sbox_out[41]), .B1(n2393), .Y(top_core_EC_ss_n130) );
  OAI2BB2X1 U17292 ( .B0(n1515), .B1(n15668), .A0N(n1515), .A1N(n15669), .Y(
        top_core_EC_ss_sbox_out[41]) );
  OAI222XL U17293 ( .A0(n10995), .A1(n10966), .B0(n10996), .B1(n10968), .C0(
        n1530), .C1(n10997), .Y(top_core_EC_ss_sbox_out_r[105]) );
  AOI222X1 U17294 ( .A0(n15684), .A1(n3147), .B0(n5713), .B1(n15685), .C0(
        n5714), .C1(n15686), .Y(n15668) );
  AOI22X1 U17295 ( .A0(top_core_EC_ss_sbox_out_r[57]), .A1(n2405), .B0(
        top_core_EC_ss_sbox_out[121]), .B1(n2503), .Y(top_core_EC_ss_n212) );
  OAI2BB2X1 U17296 ( .B0(n1525), .B1(n18818), .A0N(n1525), .A1N(n18819), .Y(
        top_core_EC_ss_sbox_out[121]) );
  OAI222XL U17297 ( .A0(n9243), .A1(n9214), .B0(n9244), .B1(n9216), .C0(n1511), 
        .C1(n9245), .Y(top_core_EC_ss_sbox_out_r[57]) );
  AOI222X1 U17298 ( .A0(n18834), .A1(n2545), .B0(n4855), .B1(n18835), .C0(
        n4856), .C1(n18836), .Y(n18818) );
  AOI22X1 U17299 ( .A0(top_core_EC_ss_sbox_out_r[88]), .A1(n2448), .B0(
        top_core_EC_ss_sbox_out[24]), .B1(n2513), .Y(top_core_EC_ss_n178) );
  OAI21XL U17300 ( .A0(n1502), .A1(n10436), .B0(n10437), .Y(
        top_core_EC_ss_sbox_out_r[88]) );
  OAI22X1 U17301 ( .A0(n15066), .A1(n1090), .B0(n1520), .B1(n15067), .Y(
        top_core_EC_ss_sbox_out[24]) );
  AOI222X1 U17302 ( .A0(n2787), .A1(n10451), .B0(n10201), .B1(n10452), .C0(
        n5237), .C1(n10453), .Y(n10436) );
  AOI22X1 U17303 ( .A0(top_core_EC_ss_sbox_out_r[9]), .A1(n2444), .B0(
        top_core_EC_ss_sbox_out[73]), .B1(n2392), .Y(top_core_EC_ss_n194) );
  OAI2BB2X1 U17304 ( .B0(n1507), .B1(n16928), .A0N(n1507), .A1N(n16929), .Y(
        top_core_EC_ss_sbox_out[73]) );
  OAI222XL U17305 ( .A0(n7491), .A1(n7462), .B0(n7492), .B1(n7464), .C0(n1524), 
        .C1(n7493), .Y(top_core_EC_ss_sbox_out_r[9]) );
  AOI222X1 U17306 ( .A0(n16944), .A1(n2909), .B0(n5409), .B1(n16945), .C0(
        n5410), .C1(n16946), .Y(n16928) );
  AOI22X1 U17307 ( .A0(top_core_EC_ss_sbox_out_r[89]), .A1(n2526), .B0(
        top_core_EC_ss_sbox_out[25]), .B1(n2509), .Y(top_core_EC_ss_n177) );
  OAI2BB2X1 U17308 ( .B0(n1520), .B1(n15038), .A0N(n1520), .A1N(n15039), .Y(
        top_core_EC_ss_sbox_out[25]) );
  OAI222XL U17309 ( .A0(n10411), .A1(n10382), .B0(n10412), .B1(n10384), .C0(
        n1502), .C1(n10413), .Y(top_core_EC_ss_sbox_out_r[89]) );
  AOI222X1 U17310 ( .A0(n15054), .A1(n3269), .B0(n5873), .B1(n15055), .C0(
        n5874), .C1(n15056), .Y(n15038) );
  AOI22X1 U17311 ( .A0(top_core_EC_ss_sbox_out_r[90]), .A1(n2531), .B0(
        top_core_EC_ss_sbox_out[26]), .B1(n2510), .Y(top_core_EC_ss_n176) );
  OAI222XL U17312 ( .A0(n15005), .A1(n14782), .B0(n15006), .B1(n14784), .C0(
        n1520), .C1(n15007), .Y(top_core_EC_ss_sbox_out[26]) );
  OAI222XL U17313 ( .A0(n10381), .A1(n10382), .B0(n10383), .B1(n10384), .C0(
        n1502), .C1(n10385), .Y(top_core_EC_ss_sbox_out_r[90]) );
  AOI221X1 U17314 ( .A0(n14978), .A1(n3311), .B0(n3284), .B1(n15023), .C0(
        n15024), .Y(n15006) );
  AOI22X1 U17315 ( .A0(top_core_EC_ss_sbox_out_r[91]), .A1(n2528), .B0(
        top_core_EC_ss_sbox_out[27]), .B1(n2503), .Y(top_core_EC_ss_n175) );
  OAI21XL U17316 ( .A0(n1520), .A1(n14971), .B0(n14972), .Y(
        top_core_EC_ss_sbox_out[27]) );
  OAI22X1 U17317 ( .A0(n10348), .A1(n978), .B0(n1502), .B1(n10349), .Y(
        top_core_EC_ss_sbox_out_r[91]) );
  AOI211X1 U17318 ( .A0(n14846), .A1(n14991), .B0(n5872), .C0(n14992), .Y(
        n14971) );
  AOI22X1 U17319 ( .A0(top_core_EC_ss_sbox_out_r[93]), .A1(n2475), .B0(
        top_core_EC_ss_sbox_out[29]), .B1(n2504), .Y(top_core_EC_ss_n172) );
  OAI222XL U17320 ( .A0(n14897), .A1(n14784), .B0(n1520), .B1(n14898), .C0(
        n14899), .C1(n14782), .Y(top_core_EC_ss_sbox_out[29]) );
  OAI222XL U17321 ( .A0(n10269), .A1(n10224), .B0(n10270), .B1(n10226), .C0(
        n10271), .C1(n978), .Y(top_core_EC_ss_sbox_out_r[93]) );
  AOI222X1 U17322 ( .A0(n3282), .A1(n14900), .B0(n14901), .B1(n3285), .C0(
        n5878), .C1(n14902), .Y(n14899) );
  AOI22X1 U17323 ( .A0(top_core_EC_ss_sbox_out_r[94]), .A1(n2474), .B0(
        top_core_EC_ss_sbox_out[30]), .B1(n2501), .Y(top_core_EC_ss_n171) );
  OAI22X1 U17324 ( .A0(n1520), .A1(n14843), .B0(n14844), .B1(n1090), .Y(
        top_core_EC_ss_sbox_out[30]) );
  OAI222XL U17325 ( .A0(n10223), .A1(n10224), .B0(n10225), .B1(n10226), .C0(
        n10227), .C1(n978), .Y(top_core_EC_ss_sbox_out_r[94]) );
  AOI211X1 U17326 ( .A0(n14873), .A1(n3271), .B0(n14874), .C0(n14875), .Y(
        n14843) );
  AOI22X1 U17327 ( .A0(top_core_EC_ss_sbox_out_r[95]), .A1(n2473), .B0(
        top_core_EC_ss_sbox_out[31]), .B1(n2502), .Y(top_core_EC_ss_n170) );
  OAI22X1 U17328 ( .A0(n1502), .A1(n10169), .B0(n10170), .B1(n978), .Y(
        top_core_EC_ss_sbox_out_r[95]) );
  OAI222XL U17329 ( .A0(n14781), .A1(n14782), .B0(n14783), .B1(n14784), .C0(
        n1520), .C1(n14785), .Y(top_core_EC_ss_sbox_out[31]) );
  AOI222X1 U17330 ( .A0(n2787), .A1(n10200), .B0(n10201), .B1(n10202), .C0(
        n5237), .C1(n10203), .Y(n10169) );
  AOI22X1 U17331 ( .A0(top_core_EC_ss_sbox_out_r[64]), .A1(n2449), .B0(
        top_core_EC_ss_sbox_out[64]), .B1(n2508), .Y(top_core_EC_ss_n169) );
  OAI21XL U17332 ( .A0(n1509), .A1(n9560), .B0(n9561), .Y(
        top_core_EC_ss_sbox_out_r[64]) );
  OAI22X1 U17333 ( .A0(n16641), .A1(n1020), .B0(n1509), .B1(n16642), .Y(
        top_core_EC_ss_sbox_out[64]) );
  AOI222X1 U17334 ( .A0(n2969), .A1(n9575), .B0(n9325), .B1(n9576), .C0(n5481), 
        .C1(n9577), .Y(n9560) );
  AOI22X1 U17335 ( .A0(top_core_EC_ss_sbox_out_r[65]), .A1(n2449), .B0(
        top_core_EC_ss_sbox_out[65]), .B1(n2507), .Y(top_core_EC_ss_n168) );
  OAI2BB2X1 U17336 ( .B0(n1509), .B1(n16613), .A0N(n1509), .A1N(n16614), .Y(
        top_core_EC_ss_sbox_out[65]) );
  OAI222XL U17337 ( .A0(n9535), .A1(n9506), .B0(n9536), .B1(n9508), .C0(n1509), 
        .C1(n9537), .Y(top_core_EC_ss_sbox_out_r[65]) );
  AOI222X1 U17338 ( .A0(n16629), .A1(n2970), .B0(n5485), .B1(n16630), .C0(
        n5486), .C1(n16631), .Y(n16613) );
  AOI22X1 U17339 ( .A0(top_core_EC_ss_sbox_out_r[66]), .A1(n2449), .B0(
        top_core_EC_ss_sbox_out[66]), .B1(n2506), .Y(top_core_EC_ss_n167) );
  OAI222XL U17340 ( .A0(n16580), .A1(n16357), .B0(n16581), .B1(n16359), .C0(
        n1509), .C1(n16582), .Y(top_core_EC_ss_sbox_out[66]) );
  OAI222XL U17341 ( .A0(n9505), .A1(n9506), .B0(n9507), .B1(n9508), .C0(n1509), 
        .C1(n9509), .Y(top_core_EC_ss_sbox_out_r[66]) );
  AOI221X1 U17342 ( .A0(n16553), .A1(n3012), .B0(n2985), .B1(n16598), .C0(
        n16599), .Y(n16581) );
  AOI22X1 U17343 ( .A0(top_core_EC_ss_sbox_out_r[67]), .A1(n2450), .B0(
        top_core_EC_ss_sbox_out[67]), .B1(n2505), .Y(top_core_EC_ss_n166) );
  OAI21XL U17344 ( .A0(n1509), .A1(n16546), .B0(n16547), .Y(
        top_core_EC_ss_sbox_out[67]) );
  OAI22X1 U17345 ( .A0(n9472), .A1(n1020), .B0(n1509), .B1(n9473), .Y(
        top_core_EC_ss_sbox_out_r[67]) );
  AOI211X1 U17346 ( .A0(n16421), .A1(n16566), .B0(n5484), .C0(n16567), .Y(
        n16546) );
  AOI22X1 U17347 ( .A0(top_core_EC_ss_sbox_out_r[69]), .A1(n2450), .B0(
        top_core_EC_ss_sbox_out[69]), .B1(n2507), .Y(top_core_EC_ss_n164) );
  OAI222XL U17348 ( .A0(n16472), .A1(n16359), .B0(n1509), .B1(n16473), .C0(
        n16474), .C1(n16357), .Y(top_core_EC_ss_sbox_out[69]) );
  OAI222XL U17349 ( .A0(n9393), .A1(n9348), .B0(n9394), .B1(n9350), .C0(n9395), 
        .C1(n1020), .Y(top_core_EC_ss_sbox_out_r[69]) );
  AOI222X1 U17350 ( .A0(n2983), .A1(n16475), .B0(n16476), .B1(n2986), .C0(
        n5490), .C1(n16477), .Y(n16474) );
  AOI22X1 U17351 ( .A0(top_core_EC_ss_sbox_out_r[70]), .A1(n2451), .B0(
        top_core_EC_ss_sbox_out[70]), .B1(n2506), .Y(top_core_EC_ss_n162) );
  OAI22X1 U17352 ( .A0(n1509), .A1(n16418), .B0(n16419), .B1(n1020), .Y(
        top_core_EC_ss_sbox_out[70]) );
  OAI222XL U17353 ( .A0(n9347), .A1(n9348), .B0(n9349), .B1(n9350), .C0(n9351), 
        .C1(n1020), .Y(top_core_EC_ss_sbox_out_r[70]) );
  AOI211X1 U17354 ( .A0(n16448), .A1(n2972), .B0(n16449), .C0(n16450), .Y(
        n16418) );
  AOI22X1 U17355 ( .A0(top_core_EC_ss_sbox_out_r[71]), .A1(n2451), .B0(
        top_core_EC_ss_sbox_out[71]), .B1(n2505), .Y(top_core_EC_ss_n161) );
  OAI22X1 U17356 ( .A0(n1509), .A1(n9293), .B0(n9294), .B1(n1020), .Y(
        top_core_EC_ss_sbox_out_r[71]) );
  OAI222XL U17357 ( .A0(n16356), .A1(n16357), .B0(n16358), .B1(n16359), .C0(
        n1509), .C1(n16360), .Y(top_core_EC_ss_sbox_out[71]) );
  AOI222X1 U17358 ( .A0(n2969), .A1(n9324), .B0(n9325), .B1(n9326), .C0(n5481), 
        .C1(n9327), .Y(n9293) );
  AOI22X1 U17359 ( .A0(top_core_EC_ss_sbox_out_r[40]), .A1(n2452), .B0(
        top_core_EC_ss_sbox_out[104]), .B1(n2535), .Y(top_core_EC_ss_n160) );
  OAI21XL U17360 ( .A0(n1515), .A1(n8684), .B0(n8685), .Y(
        top_core_EC_ss_sbox_out_r[40]) );
  OAI22X1 U17361 ( .A0(n18216), .A1(n950), .B0(n1530), .B1(n18217), .Y(
        top_core_EC_ss_sbox_out[104]) );
  AOI222X1 U17362 ( .A0(n3146), .A1(n8699), .B0(n8449), .B1(n8700), .C0(n5709), 
        .C1(n8701), .Y(n8684) );
  AOI22X1 U17363 ( .A0(top_core_EC_ss_sbox_out_r[41]), .A1(n2452), .B0(
        top_core_EC_ss_sbox_out[105]), .B1(n2535), .Y(top_core_EC_ss_n159) );
  OAI2BB2X1 U17364 ( .B0(n1530), .B1(n18188), .A0N(n1530), .A1N(n18189), .Y(
        top_core_EC_ss_sbox_out[105]) );
  OAI222XL U17365 ( .A0(n8659), .A1(n8630), .B0(n8660), .B1(n8632), .C0(n1515), 
        .C1(n8661), .Y(top_core_EC_ss_sbox_out_r[41]) );
  AOI222X1 U17366 ( .A0(n18204), .A1(n2667), .B0(n5055), .B1(n18205), .C0(
        n5056), .C1(n18206), .Y(n18188) );
  AOI22X1 U17367 ( .A0(top_core_EC_ss_sbox_out_r[42]), .A1(n2452), .B0(
        top_core_EC_ss_sbox_out[106]), .B1(n2371), .Y(top_core_EC_ss_n158) );
  OAI222XL U17368 ( .A0(n18155), .A1(n17932), .B0(n18156), .B1(n17934), .C0(
        n1530), .C1(n18157), .Y(top_core_EC_ss_sbox_out[106]) );
  OAI222XL U17369 ( .A0(n8629), .A1(n8630), .B0(n8631), .B1(n8632), .C0(n1515), 
        .C1(n8633), .Y(top_core_EC_ss_sbox_out_r[42]) );
  AOI221X1 U17370 ( .A0(n18128), .A1(n2703), .B0(n2682), .B1(n18173), .C0(
        n18174), .Y(n18156) );
  AOI22X1 U17371 ( .A0(top_core_EC_ss_sbox_out_r[43]), .A1(n2453), .B0(
        top_core_EC_ss_sbox_out[107]), .B1(n2375), .Y(top_core_EC_ss_n157) );
  OAI21XL U17372 ( .A0(n1530), .A1(n18121), .B0(n18122), .Y(
        top_core_EC_ss_sbox_out[107]) );
  OAI22X1 U17373 ( .A0(n8596), .A1(n1062), .B0(n1515), .B1(n8597), .Y(
        top_core_EC_ss_sbox_out_r[43]) );
  AOI211X1 U17374 ( .A0(n17996), .A1(n18141), .B0(n5054), .C0(n18142), .Y(
        n18121) );
  AOI22X1 U17375 ( .A0(top_core_EC_ss_sbox_out_r[45]), .A1(n2453), .B0(
        top_core_EC_ss_sbox_out[109]), .B1(n2500), .Y(top_core_EC_ss_n155) );
  OAI222XL U17376 ( .A0(n18047), .A1(n17934), .B0(n1530), .B1(n18048), .C0(
        n18049), .C1(n17932), .Y(top_core_EC_ss_sbox_out[109]) );
  OAI222XL U17377 ( .A0(n8517), .A1(n8472), .B0(n8518), .B1(n8474), .C0(n8519), 
        .C1(n1062), .Y(top_core_EC_ss_sbox_out_r[45]) );
  AOI222X1 U17378 ( .A0(n2681), .A1(n18050), .B0(n18051), .B1(n2683), .C0(
        n5060), .C1(n18052), .Y(n18049) );
  AOI22X1 U17379 ( .A0(top_core_EC_ss_sbox_out_r[46]), .A1(n2454), .B0(
        top_core_EC_ss_sbox_out[110]), .B1(n2499), .Y(top_core_EC_ss_n154) );
  OAI22X1 U17380 ( .A0(n1530), .A1(n17993), .B0(n17994), .B1(n950), .Y(
        top_core_EC_ss_sbox_out[110]) );
  OAI222XL U17381 ( .A0(n8471), .A1(n8472), .B0(n8473), .B1(n8474), .C0(n8475), 
        .C1(n1062), .Y(top_core_EC_ss_sbox_out_r[46]) );
  AOI211X1 U17382 ( .A0(n18023), .A1(n2669), .B0(n18024), .C0(n18025), .Y(
        n17993) );
  AOI22X1 U17383 ( .A0(top_core_EC_ss_sbox_out_r[47]), .A1(n2454), .B0(
        top_core_EC_ss_sbox_out[111]), .B1(n2498), .Y(top_core_EC_ss_n153) );
  OAI22X1 U17384 ( .A0(n1515), .A1(n8417), .B0(n8418), .B1(n1062), .Y(
        top_core_EC_ss_sbox_out_r[47]) );
  OAI222XL U17385 ( .A0(n17931), .A1(n17932), .B0(n17933), .B1(n17934), .C0(
        n1530), .C1(n17935), .Y(top_core_EC_ss_sbox_out[111]) );
  AOI222X1 U17386 ( .A0(n3146), .A1(n8448), .B0(n8449), .B1(n8450), .C0(n5709), 
        .C1(n8451), .Y(n8417) );
  AOI22X1 U17387 ( .A0(top_core_EC_ss_sbox_out_r[16]), .A1(n2455), .B0(
        top_core_EC_ss_sbox_out[16]), .B1(n2394), .Y(top_core_EC_ss_n151) );
  OAI21XL U17388 ( .A0(n1522), .A1(n7808), .B0(n7809), .Y(
        top_core_EC_ss_sbox_out_r[16]) );
  OAI22X1 U17389 ( .A0(n14751), .A1(n1104), .B0(n1522), .B1(n14752), .Y(
        top_core_EC_ss_sbox_out[16]) );
  AOI222X1 U17390 ( .A0(n3329), .A1(n7823), .B0(n7573), .B1(n7824), .C0(n5945), 
        .C1(n7825), .Y(n7808) );
  AOI22X1 U17391 ( .A0(top_core_EC_ss_sbox_out_r[17]), .A1(n2455), .B0(
        top_core_EC_ss_sbox_out[17]), .B1(n2394), .Y(top_core_EC_ss_n150) );
  OAI2BB2X1 U17392 ( .B0(n1522), .B1(n14723), .A0N(n1522), .A1N(n14724), .Y(
        top_core_EC_ss_sbox_out[17]) );
  OAI222XL U17393 ( .A0(n7783), .A1(n7754), .B0(n7784), .B1(n7756), .C0(n1522), 
        .C1(n7785), .Y(top_core_EC_ss_sbox_out_r[17]) );
  AOI222X1 U17394 ( .A0(n14739), .A1(n3330), .B0(n5949), .B1(n14740), .C0(
        n5950), .C1(n14741), .Y(n14723) );
  AOI22X1 U17395 ( .A0(top_core_EC_ss_sbox_out_r[18]), .A1(n2455), .B0(
        top_core_EC_ss_sbox_out[18]), .B1(n2394), .Y(top_core_EC_ss_n149) );
  OAI222XL U17396 ( .A0(n14690), .A1(n14467), .B0(n14691), .B1(n14469), .C0(
        n1522), .C1(n14692), .Y(top_core_EC_ss_sbox_out[18]) );
  OAI222XL U17397 ( .A0(n7753), .A1(n7754), .B0(n7755), .B1(n7756), .C0(n1522), 
        .C1(n7757), .Y(top_core_EC_ss_sbox_out_r[18]) );
  AOI221X1 U17398 ( .A0(n14663), .A1(n3366), .B0(n3345), .B1(n14708), .C0(
        n14709), .Y(n14691) );
  AOI22X1 U17399 ( .A0(top_core_EC_ss_sbox_out_r[19]), .A1(n2456), .B0(
        top_core_EC_ss_sbox_out[19]), .B1(n2394), .Y(top_core_EC_ss_n148) );
  OAI21XL U17400 ( .A0(n1522), .A1(n14656), .B0(n14657), .Y(
        top_core_EC_ss_sbox_out[19]) );
  OAI22X1 U17401 ( .A0(n7720), .A1(n1104), .B0(n1522), .B1(n7721), .Y(
        top_core_EC_ss_sbox_out_r[19]) );
  AOI211X1 U17402 ( .A0(n14531), .A1(n14676), .B0(n5948), .C0(n14677), .Y(
        n14656) );
  AOI22X1 U17403 ( .A0(top_core_EC_ss_sbox_out_r[21]), .A1(n2456), .B0(
        top_core_EC_ss_sbox_out[21]), .B1(n2394), .Y(top_core_EC_ss_n146) );
  OAI222XL U17404 ( .A0(n14582), .A1(n14469), .B0(n1522), .B1(n14583), .C0(
        n14584), .C1(n14467), .Y(top_core_EC_ss_sbox_out[21]) );
  OAI222XL U17405 ( .A0(n7641), .A1(n7596), .B0(n7642), .B1(n7598), .C0(n7643), 
        .C1(n1104), .Y(top_core_EC_ss_sbox_out_r[21]) );
  AOI222X1 U17406 ( .A0(n3343), .A1(n14585), .B0(n14586), .B1(n3347), .C0(
        n5954), .C1(n14587), .Y(n14584) );
  AOI22X1 U17407 ( .A0(top_core_EC_ss_sbox_out_r[22]), .A1(n2457), .B0(
        top_core_EC_ss_sbox_out[22]), .B1(n2394), .Y(top_core_EC_ss_n145) );
  OAI22X1 U17408 ( .A0(n1522), .A1(n14528), .B0(n14529), .B1(n1104), .Y(
        top_core_EC_ss_sbox_out[22]) );
  OAI222XL U17409 ( .A0(n7595), .A1(n7596), .B0(n7597), .B1(n7598), .C0(n7599), 
        .C1(n1104), .Y(top_core_EC_ss_sbox_out_r[22]) );
  AOI211X1 U17410 ( .A0(n14558), .A1(n3332), .B0(n14559), .C0(n14560), .Y(
        n14528) );
  AOI22X1 U17411 ( .A0(top_core_EC_ss_sbox_out_r[23]), .A1(n2457), .B0(
        top_core_EC_ss_sbox_out[23]), .B1(n2394), .Y(top_core_EC_ss_n144) );
  OAI22X1 U17412 ( .A0(n1522), .A1(n7541), .B0(n7542), .B1(n1104), .Y(
        top_core_EC_ss_sbox_out_r[23]) );
  OAI222XL U17413 ( .A0(n14466), .A1(n14467), .B0(n14468), .B1(n14469), .C0(
        n1522), .C1(n14470), .Y(top_core_EC_ss_sbox_out[23]) );
  AOI222X1 U17414 ( .A0(n3329), .A1(n7572), .B0(n7573), .B1(n7574), .C0(n5945), 
        .C1(n7575), .Y(n7541) );
  AOI22X1 U17415 ( .A0(top_core_EC_ss_sbox_out_r[120]), .A1(n2457), .B0(
        top_core_EC_ss_sbox_out[56]), .B1(n2394), .Y(top_core_EC_ss_n143) );
  OAI21XL U17416 ( .A0(n1525), .A1(n11604), .B0(n11605), .Y(
        top_core_EC_ss_sbox_out_r[120]) );
  OAI22X1 U17417 ( .A0(n16326), .A1(n1034), .B0(n1511), .B1(n16327), .Y(
        top_core_EC_ss_sbox_out[56]) );
  AOI222X1 U17418 ( .A0(n2544), .A1(n11619), .B0(n11369), .B1(n11620), .C0(
        n4851), .C1(n11621), .Y(n11604) );
  AOI22X1 U17419 ( .A0(top_core_EC_ss_sbox_out_r[121]), .A1(n2458), .B0(
        top_core_EC_ss_sbox_out[57]), .B1(n2394), .Y(top_core_EC_ss_n142) );
  OAI2BB2X1 U17420 ( .B0(n1511), .B1(n16298), .A0N(n1511), .A1N(n16299), .Y(
        top_core_EC_ss_sbox_out[57]) );
  OAI222XL U17421 ( .A0(n11579), .A1(n11550), .B0(n11580), .B1(n11552), .C0(
        n1525), .C1(n11581), .Y(top_core_EC_ss_sbox_out_r[121]) );
  AOI222X1 U17422 ( .A0(n16314), .A1(n3028), .B0(n5561), .B1(n16315), .C0(
        n5562), .C1(n16316), .Y(n16298) );
  AOI22X1 U17423 ( .A0(top_core_EC_ss_sbox_out_r[122]), .A1(n2458), .B0(
        top_core_EC_ss_sbox_out[58]), .B1(n2394), .Y(top_core_EC_ss_n140) );
  OAI222XL U17424 ( .A0(n16265), .A1(n16042), .B0(n16266), .B1(n16044), .C0(
        n1511), .C1(n16267), .Y(top_core_EC_ss_sbox_out[58]) );
  OAI222XL U17425 ( .A0(n11549), .A1(n11550), .B0(n11551), .B1(n11552), .C0(
        n1525), .C1(n11553), .Y(top_core_EC_ss_sbox_out_r[122]) );
  AOI221X1 U17426 ( .A0(n16238), .A1(n3065), .B0(n3043), .B1(n16283), .C0(
        n16284), .Y(n16266) );
  AOI22X1 U17427 ( .A0(top_core_EC_ss_sbox_out_r[123]), .A1(n2459), .B0(
        top_core_EC_ss_sbox_out[59]), .B1(n2394), .Y(top_core_EC_ss_n139) );
  OAI21XL U17428 ( .A0(n1511), .A1(n16231), .B0(n16232), .Y(
        top_core_EC_ss_sbox_out[59]) );
  OAI22X1 U17429 ( .A0(n11516), .A1(n922), .B0(n1525), .B1(n11517), .Y(
        top_core_EC_ss_sbox_out_r[123]) );
  AOI211X1 U17430 ( .A0(n16106), .A1(n16251), .B0(n5560), .C0(n16252), .Y(
        n16231) );
  AOI22X1 U17431 ( .A0(top_core_EC_ss_sbox_out_r[125]), .A1(n2459), .B0(
        top_core_EC_ss_sbox_out[61]), .B1(n2393), .Y(top_core_EC_ss_n137) );
  OAI222XL U17432 ( .A0(n16157), .A1(n16044), .B0(n1511), .B1(n16158), .C0(
        n16159), .C1(n16042), .Y(top_core_EC_ss_sbox_out[61]) );
  OAI222XL U17433 ( .A0(n11437), .A1(n11392), .B0(n11438), .B1(n11394), .C0(
        n11439), .C1(n922), .Y(top_core_EC_ss_sbox_out_r[125]) );
  AOI222X1 U17434 ( .A0(n3041), .A1(n16160), .B0(n16161), .B1(n3045), .C0(
        n5566), .C1(n16162), .Y(n16159) );
  AOI22X1 U17435 ( .A0(top_core_EC_ss_sbox_out_r[126]), .A1(n2460), .B0(
        top_core_EC_ss_sbox_out[62]), .B1(n2393), .Y(top_core_EC_ss_n136) );
  OAI22X1 U17436 ( .A0(n1511), .A1(n16103), .B0(n16104), .B1(n1034), .Y(
        top_core_EC_ss_sbox_out[62]) );
  OAI222XL U17437 ( .A0(n11391), .A1(n11392), .B0(n11393), .B1(n11394), .C0(
        n11395), .C1(n922), .Y(top_core_EC_ss_sbox_out_r[126]) );
  AOI211X1 U17438 ( .A0(n16133), .A1(n3030), .B0(n16134), .C0(n16135), .Y(
        n16103) );
  AOI22X1 U17439 ( .A0(top_core_EC_ss_sbox_out_r[127]), .A1(n2460), .B0(
        top_core_EC_ss_sbox_out[63]), .B1(n2393), .Y(top_core_EC_ss_n135) );
  OAI22X1 U17440 ( .A0(n1525), .A1(n11337), .B0(n11338), .B1(n922), .Y(
        top_core_EC_ss_sbox_out_r[127]) );
  OAI222XL U17441 ( .A0(n16041), .A1(n16042), .B0(n16043), .B1(n16044), .C0(
        n1511), .C1(n16045), .Y(top_core_EC_ss_sbox_out[63]) );
  AOI222X1 U17442 ( .A0(n2544), .A1(n11368), .B0(n11369), .B1(n11370), .C0(
        n4851), .C1(n11371), .Y(n11337) );
  AOI22X1 U17443 ( .A0(top_core_EC_ss_sbox_out_r[96]), .A1(n2460), .B0(
        top_core_EC_ss_sbox_out[96]), .B1(n2393), .Y(top_core_EC_ss_n134) );
  OAI21XL U17444 ( .A0(n1532), .A1(n10728), .B0(n10729), .Y(
        top_core_EC_ss_sbox_out_r[96]) );
  OAI22X1 U17445 ( .A0(n17901), .A1(n964), .B0(n1532), .B1(n17902), .Y(
        top_core_EC_ss_sbox_out[96]) );
  AOI222X1 U17446 ( .A0(n2726), .A1(n10743), .B0(n10493), .B1(n10744), .C0(
        n5159), .C1(n10745), .Y(n10728) );
  AOI22X1 U17447 ( .A0(top_core_EC_ss_sbox_out_r[97]), .A1(n2464), .B0(
        top_core_EC_ss_sbox_out[97]), .B1(n2384), .Y(top_core_EC_ss_n133) );
  OAI2BB2X1 U17448 ( .B0(n1532), .B1(n17873), .A0N(n1532), .A1N(n17874), .Y(
        top_core_EC_ss_sbox_out[97]) );
  OAI222XL U17449 ( .A0(n10703), .A1(n10674), .B0(n10704), .B1(n10676), .C0(
        n1532), .C1(n10705), .Y(top_core_EC_ss_sbox_out_r[97]) );
  AOI222X1 U17450 ( .A0(n17889), .A1(n2727), .B0(n5163), .B1(n17890), .C0(
        n5164), .C1(n17891), .Y(n17873) );
  AOI22X1 U17451 ( .A0(top_core_EC_ss_sbox_out_r[98]), .A1(n2461), .B0(
        top_core_EC_ss_sbox_out[98]), .B1(n2372), .Y(top_core_EC_ss_n132) );
  OAI222XL U17452 ( .A0(n17840), .A1(n17617), .B0(n17841), .B1(n17619), .C0(
        n1532), .C1(n17842), .Y(top_core_EC_ss_sbox_out[98]) );
  OAI222XL U17453 ( .A0(n10673), .A1(n10674), .B0(n10675), .B1(n10676), .C0(
        n1532), .C1(n10677), .Y(top_core_EC_ss_sbox_out_r[98]) );
  AOI221X1 U17454 ( .A0(n17813), .A1(n2763), .B0(n2742), .B1(n17858), .C0(
        n17859), .Y(n17841) );
  AOI22X1 U17455 ( .A0(top_core_EC_ss_sbox_out_r[99]), .A1(n2461), .B0(
        top_core_EC_ss_sbox_out[99]), .B1(n2538), .Y(top_core_EC_ss_n131) );
  OAI21XL U17456 ( .A0(n1532), .A1(n17806), .B0(n17807), .Y(
        top_core_EC_ss_sbox_out[99]) );
  OAI22X1 U17457 ( .A0(n10640), .A1(n964), .B0(n1532), .B1(n10641), .Y(
        top_core_EC_ss_sbox_out_r[99]) );
  AOI211X1 U17458 ( .A0(n17681), .A1(n17826), .B0(n5162), .C0(n17827), .Y(
        n17806) );
  AOI22X1 U17459 ( .A0(top_core_EC_ss_sbox_out_r[101]), .A1(n2475), .B0(
        top_core_EC_ss_sbox_out[101]), .B1(n2539), .Y(top_core_EC_ss_n255) );
  OAI222XL U17460 ( .A0(n17732), .A1(n17619), .B0(n1532), .B1(n17733), .C0(
        n17734), .C1(n17617), .Y(top_core_EC_ss_sbox_out[101]) );
  OAI222XL U17461 ( .A0(n10561), .A1(n10516), .B0(n10562), .B1(n10518), .C0(
        n10563), .C1(n964), .Y(top_core_EC_ss_sbox_out_r[101]) );
  AOI222X1 U17462 ( .A0(n2741), .A1(n17735), .B0(n17736), .B1(n2743), .C0(
        n5168), .C1(n17737), .Y(n17734) );
  AOI22X1 U17463 ( .A0(top_core_EC_ss_sbox_out_r[102]), .A1(n2475), .B0(
        top_core_EC_ss_sbox_out[102]), .B1(n2536), .Y(top_core_EC_ss_n254) );
  OAI22X1 U17464 ( .A0(n1532), .A1(n17678), .B0(n17679), .B1(n964), .Y(
        top_core_EC_ss_sbox_out[102]) );
  OAI222XL U17465 ( .A0(n10515), .A1(n10516), .B0(n10517), .B1(n10518), .C0(
        n10519), .C1(n964), .Y(top_core_EC_ss_sbox_out_r[102]) );
  AOI211X1 U17466 ( .A0(n17708), .A1(n2729), .B0(n17709), .C0(n17710), .Y(
        n17678) );
  AOI22X1 U17467 ( .A0(top_core_EC_ss_sbox_out_r[103]), .A1(n2474), .B0(
        top_core_EC_ss_sbox_out[103]), .B1(n2537), .Y(top_core_EC_ss_n253) );
  OAI22X1 U17468 ( .A0(n1532), .A1(n10461), .B0(n10462), .B1(n964), .Y(
        top_core_EC_ss_sbox_out_r[103]) );
  OAI222XL U17469 ( .A0(n17616), .A1(n17617), .B0(n17618), .B1(n17619), .C0(
        n1532), .C1(n17620), .Y(top_core_EC_ss_sbox_out[103]) );
  AOI222X1 U17470 ( .A0(n2726), .A1(n10492), .B0(n10493), .B1(n10494), .C0(
        n5159), .C1(n10495), .Y(n10461) );
  AOI22X1 U17471 ( .A0(top_core_EC_ss_sbox_out_r[72]), .A1(n2474), .B0(
        top_core_EC_ss_sbox_out[8]), .B1(n2376), .Y(top_core_EC_ss_n252) );
  OAI21XL U17472 ( .A0(n1507), .A1(n9852), .B0(n9853), .Y(
        top_core_EC_ss_sbox_out_r[72]) );
  OAI22X1 U17473 ( .A0(n14436), .A1(n1118), .B0(n1524), .B1(n14437), .Y(
        top_core_EC_ss_sbox_out[8]) );
  AOI222X1 U17474 ( .A0(n2908), .A1(n9867), .B0(n9617), .B1(n9868), .C0(n5405), 
        .C1(n9869), .Y(n9852) );
  AOI22X1 U17475 ( .A0(top_core_EC_ss_sbox_out_r[73]), .A1(n2474), .B0(
        top_core_EC_ss_sbox_out[9]), .B1(n2394), .Y(top_core_EC_ss_n251) );
  OAI2BB2X1 U17476 ( .B0(n1524), .B1(n14408), .A0N(n1524), .A1N(n14409), .Y(
        top_core_EC_ss_sbox_out[9]) );
  OAI222XL U17477 ( .A0(n9827), .A1(n9798), .B0(n9828), .B1(n9800), .C0(n1507), 
        .C1(n9829), .Y(top_core_EC_ss_sbox_out_r[73]) );
  AOI222X1 U17478 ( .A0(n14424), .A1(n3388), .B0(n6025), .B1(n14425), .C0(
        n6026), .C1(n14426), .Y(n14408) );
  AOI22X1 U17479 ( .A0(top_core_EC_ss_sbox_out_r[74]), .A1(n2473), .B0(
        top_core_EC_ss_sbox_out[10]), .B1(n2375), .Y(top_core_EC_ss_n250) );
  OAI222XL U17480 ( .A0(n14375), .A1(n14152), .B0(n14376), .B1(n14154), .C0(
        n1524), .C1(n14377), .Y(top_core_EC_ss_sbox_out[10]) );
  OAI222XL U17481 ( .A0(n9797), .A1(n9798), .B0(n9799), .B1(n9800), .C0(n1507), 
        .C1(n9801), .Y(top_core_EC_ss_sbox_out_r[74]) );
  AOI221X1 U17482 ( .A0(n14348), .A1(n3424), .B0(n3403), .B1(n14393), .C0(
        n14394), .Y(n14376) );
  AOI22X1 U17483 ( .A0(top_core_EC_ss_sbox_out_r[75]), .A1(n2473), .B0(
        top_core_EC_ss_sbox_out[11]), .B1(n2393), .Y(top_core_EC_ss_n249) );
  OAI21XL U17484 ( .A0(n1524), .A1(n14341), .B0(n14342), .Y(
        top_core_EC_ss_sbox_out[11]) );
  OAI22X1 U17485 ( .A0(n9764), .A1(n1006), .B0(n1507), .B1(n9765), .Y(
        top_core_EC_ss_sbox_out_r[75]) );
  AOI211X1 U17486 ( .A0(n14216), .A1(n14361), .B0(n6024), .C0(n14362), .Y(
        n14341) );
  AOI22X1 U17487 ( .A0(top_core_EC_ss_sbox_out_r[77]), .A1(n2472), .B0(
        top_core_EC_ss_sbox_out[13]), .B1(n2392), .Y(top_core_EC_ss_n247) );
  OAI222XL U17488 ( .A0(n14267), .A1(n14154), .B0(n1524), .B1(n14268), .C0(
        n14269), .C1(n14152), .Y(top_core_EC_ss_sbox_out[13]) );
  OAI222XL U17489 ( .A0(n9685), .A1(n9640), .B0(n9686), .B1(n9642), .C0(n9687), 
        .C1(n1006), .Y(top_core_EC_ss_sbox_out_r[77]) );
  AOI222X1 U17490 ( .A0(n3401), .A1(n14270), .B0(n14271), .B1(n3405), .C0(
        n6030), .C1(n14272), .Y(n14269) );
  AOI22X1 U17491 ( .A0(top_core_EC_ss_sbox_out_r[78]), .A1(n2472), .B0(
        top_core_EC_ss_sbox_out[14]), .B1(n2384), .Y(top_core_EC_ss_n245) );
  OAI22X1 U17492 ( .A0(n1524), .A1(n14213), .B0(n14214), .B1(n1118), .Y(
        top_core_EC_ss_sbox_out[14]) );
  OAI222XL U17493 ( .A0(n9639), .A1(n9640), .B0(n9641), .B1(n9642), .C0(n9643), 
        .C1(n1006), .Y(top_core_EC_ss_sbox_out_r[78]) );
  AOI211X1 U17494 ( .A0(n14243), .A1(n3390), .B0(n14244), .C0(n14245), .Y(
        n14213) );
  AOI22X1 U17495 ( .A0(top_core_EC_ss_sbox_out_r[79]), .A1(n2471), .B0(
        top_core_EC_ss_sbox_out[15]), .B1(n2376), .Y(top_core_EC_ss_n244) );
  OAI22X1 U17496 ( .A0(n1507), .A1(n9585), .B0(n9586), .B1(n1006), .Y(
        top_core_EC_ss_sbox_out_r[79]) );
  OAI222XL U17497 ( .A0(n14151), .A1(n14152), .B0(n14153), .B1(n14154), .C0(
        n1524), .C1(n14155), .Y(top_core_EC_ss_sbox_out[15]) );
  AOI222X1 U17498 ( .A0(n2908), .A1(n9616), .B0(n9617), .B1(n9618), .C0(n5405), 
        .C1(n9619), .Y(n9585) );
  AOI22X1 U17499 ( .A0(top_core_EC_ss_sbox_out_r[48]), .A1(n2471), .B0(
        top_core_EC_ss_sbox_out[48]), .B1(n2383), .Y(top_core_EC_ss_n243) );
  OAI21XL U17500 ( .A0(n1513), .A1(n8976), .B0(n8977), .Y(
        top_core_EC_ss_sbox_out_r[48]) );
  OAI22X1 U17501 ( .A0(n16011), .A1(n1048), .B0(n1513), .B1(n16012), .Y(
        top_core_EC_ss_sbox_out[48]) );
  AOI222X1 U17502 ( .A0(n3088), .A1(n8991), .B0(n8741), .B1(n8992), .C0(n5633), 
        .C1(n8993), .Y(n8976) );
  AOI22X1 U17503 ( .A0(top_core_EC_ss_sbox_out_r[49]), .A1(n2471), .B0(
        top_core_EC_ss_sbox_out[49]), .B1(n2381), .Y(top_core_EC_ss_n242) );
  OAI2BB2X1 U17504 ( .B0(n1513), .B1(n15983), .A0N(n1513), .A1N(n15984), .Y(
        top_core_EC_ss_sbox_out[49]) );
  OAI222XL U17505 ( .A0(n8951), .A1(n8922), .B0(n8952), .B1(n8924), .C0(n1513), 
        .C1(n8953), .Y(top_core_EC_ss_sbox_out_r[49]) );
  AOI222X1 U17506 ( .A0(n15999), .A1(n3089), .B0(n5637), .B1(n16000), .C0(
        n5638), .C1(n16001), .Y(n15983) );
  AOI22X1 U17507 ( .A0(top_core_EC_ss_sbox_out_r[50]), .A1(n2470), .B0(
        top_core_EC_ss_sbox_out[50]), .B1(n2382), .Y(top_core_EC_ss_n241) );
  OAI222XL U17508 ( .A0(n15950), .A1(n15727), .B0(n15951), .B1(n15729), .C0(
        n1513), .C1(n15952), .Y(top_core_EC_ss_sbox_out[50]) );
  OAI222XL U17509 ( .A0(n8921), .A1(n8922), .B0(n8923), .B1(n8924), .C0(n1513), 
        .C1(n8925), .Y(top_core_EC_ss_sbox_out_r[50]) );
  AOI221X1 U17510 ( .A0(n15923), .A1(n3125), .B0(n3104), .B1(n15968), .C0(
        n15969), .Y(n15951) );
  AOI22X1 U17511 ( .A0(top_core_EC_ss_sbox_out_r[51]), .A1(n2470), .B0(
        top_core_EC_ss_sbox_out[51]), .B1(n2380), .Y(top_core_EC_ss_n240) );
  OAI21XL U17512 ( .A0(n1513), .A1(n15916), .B0(n15917), .Y(
        top_core_EC_ss_sbox_out[51]) );
  OAI22X1 U17513 ( .A0(n8888), .A1(n1048), .B0(n1513), .B1(n8889), .Y(
        top_core_EC_ss_sbox_out_r[51]) );
  AOI211X1 U17514 ( .A0(n15791), .A1(n15936), .B0(n5636), .C0(n15937), .Y(
        n15916) );
  AOI22X1 U17515 ( .A0(top_core_EC_ss_sbox_out_r[53]), .A1(n2469), .B0(
        top_core_EC_ss_sbox_out[53]), .B1(n2378), .Y(top_core_EC_ss_n238) );
  OAI222XL U17516 ( .A0(n15842), .A1(n15729), .B0(n1513), .B1(n15843), .C0(
        n15844), .C1(n15727), .Y(top_core_EC_ss_sbox_out[53]) );
  OAI222XL U17517 ( .A0(n8809), .A1(n8764), .B0(n8810), .B1(n8766), .C0(n8811), 
        .C1(n1048), .Y(top_core_EC_ss_sbox_out_r[53]) );
  AOI222X1 U17518 ( .A0(n3103), .A1(n15845), .B0(n15846), .B1(n3105), .C0(
        n5642), .C1(n15847), .Y(n15844) );
  AOI22X1 U17519 ( .A0(top_core_EC_ss_sbox_out_r[54]), .A1(n2469), .B0(
        top_core_EC_ss_sbox_out[54]), .B1(n2379), .Y(top_core_EC_ss_n237) );
  OAI22X1 U17520 ( .A0(n1513), .A1(n15788), .B0(n15789), .B1(n1048), .Y(
        top_core_EC_ss_sbox_out[54]) );
  OAI222XL U17521 ( .A0(n8763), .A1(n8764), .B0(n8765), .B1(n8766), .C0(n8767), 
        .C1(n1048), .Y(top_core_EC_ss_sbox_out_r[54]) );
  AOI211X1 U17522 ( .A0(n15818), .A1(n3091), .B0(n15819), .C0(n15820), .Y(
        n15788) );
  AOI22X1 U17523 ( .A0(top_core_EC_ss_sbox_out_r[55]), .A1(n2469), .B0(
        top_core_EC_ss_sbox_out[55]), .B1(n2377), .Y(top_core_EC_ss_n236) );
  OAI22X1 U17524 ( .A0(n1513), .A1(n8709), .B0(n8710), .B1(n1048), .Y(
        top_core_EC_ss_sbox_out_r[55]) );
  OAI222XL U17525 ( .A0(n15726), .A1(n15727), .B0(n15728), .B1(n15729), .C0(
        n1513), .C1(n15730), .Y(top_core_EC_ss_sbox_out[55]) );
  AOI222X1 U17526 ( .A0(n3088), .A1(n8740), .B0(n8741), .B1(n8742), .C0(n5633), 
        .C1(n8743), .Y(n8709) );
  AOI22X1 U17527 ( .A0(top_core_EC_ss_sbox_out_r[24]), .A1(n2468), .B0(
        top_core_EC_ss_sbox_out[88]), .B1(n2499), .Y(top_core_EC_ss_n234) );
  OAI21XL U17528 ( .A0(n1520), .A1(n8100), .B0(n8101), .Y(
        top_core_EC_ss_sbox_out_r[24]) );
  OAI22X1 U17529 ( .A0(n17586), .A1(n978), .B0(n1502), .B1(n17587), .Y(
        top_core_EC_ss_sbox_out[88]) );
  AOI222X1 U17530 ( .A0(n3268), .A1(n8115), .B0(n7865), .B1(n8116), .C0(n5869), 
        .C1(n8117), .Y(n8100) );
  AOI22X1 U17531 ( .A0(top_core_EC_ss_sbox_out_r[25]), .A1(n2468), .B0(
        top_core_EC_ss_sbox_out[89]), .B1(n2498), .Y(top_core_EC_ss_n233) );
  OAI2BB2X1 U17532 ( .B0(n1502), .B1(n17558), .A0N(n1502), .A1N(n17559), .Y(
        top_core_EC_ss_sbox_out[89]) );
  OAI222XL U17533 ( .A0(n8075), .A1(n8046), .B0(n8076), .B1(n8048), .C0(n1520), 
        .C1(n8077), .Y(top_core_EC_ss_sbox_out_r[25]) );
  AOI222X1 U17534 ( .A0(n17574), .A1(n2788), .B0(n5241), .B1(n17575), .C0(
        n5242), .C1(n17576), .Y(n17558) );
  AOI22X1 U17535 ( .A0(top_core_EC_ss_sbox_out_r[26]), .A1(n2467), .B0(
        top_core_EC_ss_sbox_out[90]), .B1(n2497), .Y(top_core_EC_ss_n232) );
  OAI222XL U17536 ( .A0(n17525), .A1(n17302), .B0(n17526), .B1(n17304), .C0(
        n1502), .C1(n17527), .Y(top_core_EC_ss_sbox_out[90]) );
  OAI222XL U17537 ( .A0(n8045), .A1(n8046), .B0(n8047), .B1(n8048), .C0(n1520), 
        .C1(n8049), .Y(top_core_EC_ss_sbox_out_r[26]) );
  AOI221X1 U17538 ( .A0(n17498), .A1(n2825), .B0(n2803), .B1(n17543), .C0(
        n17544), .Y(n17526) );
  AOI22X1 U17539 ( .A0(top_core_EC_ss_sbox_out_r[27]), .A1(n2467), .B0(
        top_core_EC_ss_sbox_out[91]), .B1(n2374), .Y(top_core_EC_ss_n231) );
  OAI21XL U17540 ( .A0(n1502), .A1(n17491), .B0(n17492), .Y(
        top_core_EC_ss_sbox_out[91]) );
  OAI22X1 U17541 ( .A0(n8012), .A1(n1090), .B0(n1520), .B1(n8013), .Y(
        top_core_EC_ss_sbox_out_r[27]) );
  AOI211X1 U17542 ( .A0(n17366), .A1(n17511), .B0(n5240), .C0(n17512), .Y(
        n17491) );
  AOI22X1 U17543 ( .A0(top_core_EC_ss_sbox_out_r[29]), .A1(n2466), .B0(
        top_core_EC_ss_sbox_out[93]), .B1(n2383), .Y(top_core_EC_ss_n229) );
  OAI222XL U17544 ( .A0(n17417), .A1(n17304), .B0(n1502), .B1(n17418), .C0(
        n17419), .C1(n17302), .Y(top_core_EC_ss_sbox_out[93]) );
  OAI222XL U17545 ( .A0(n7933), .A1(n7888), .B0(n7934), .B1(n7890), .C0(n7935), 
        .C1(n1090), .Y(top_core_EC_ss_sbox_out_r[29]) );
  AOI222X1 U17546 ( .A0(n2801), .A1(n17420), .B0(n17421), .B1(n2804), .C0(
        n5246), .C1(n17422), .Y(n17419) );
  AOI22X1 U17547 ( .A0(top_core_EC_ss_sbox_out_r[30]), .A1(n2466), .B0(
        top_core_EC_ss_sbox_out[94]), .B1(n2378), .Y(top_core_EC_ss_n228) );
  OAI22X1 U17548 ( .A0(n1502), .A1(n17363), .B0(n17364), .B1(n978), .Y(
        top_core_EC_ss_sbox_out[94]) );
  OAI222XL U17549 ( .A0(n7887), .A1(n7888), .B0(n7889), .B1(n7890), .C0(n7891), 
        .C1(n1090), .Y(top_core_EC_ss_sbox_out_r[30]) );
  AOI211X1 U17550 ( .A0(n17393), .A1(n2790), .B0(n17394), .C0(n17395), .Y(
        n17363) );
  AOI22X1 U17551 ( .A0(top_core_EC_ss_sbox_out_r[31]), .A1(n2466), .B0(
        top_core_EC_ss_sbox_out[95]), .B1(n2496), .Y(top_core_EC_ss_n227) );
  OAI22X1 U17552 ( .A0(n1520), .A1(n7833), .B0(n7834), .B1(n1090), .Y(
        top_core_EC_ss_sbox_out_r[31]) );
  OAI222XL U17553 ( .A0(n17301), .A1(n17302), .B0(n17303), .B1(n17304), .C0(
        n1502), .C1(n17305), .Y(top_core_EC_ss_sbox_out[95]) );
  AOI222X1 U17554 ( .A0(n3268), .A1(n7864), .B0(n7865), .B1(n7866), .C0(n5869), 
        .C1(n7867), .Y(n7833) );
  INVX1 U17555 ( .A(top_core_KE_new_sboxw_15_), .Y(n6735) );
  INVX1 U17556 ( .A(top_core_KE_new_sboxw_13_), .Y(n6722) );
  INVX1 U17557 ( .A(top_core_KE_new_sboxw_10_), .Y(n6728) );
  INVX1 U17558 ( .A(top_core_KE_new_sboxw_7_), .Y(n6785) );
  INVX1 U17559 ( .A(top_core_KE_new_sboxw_5_), .Y(n6787) );
  INVX1 U17560 ( .A(top_core_KE_new_sboxw_2_), .Y(n6792) );
  INVX1 U17561 ( .A(top_core_KE_new_sboxw_31_), .Y(n6359) );
  INVX1 U17562 ( .A(top_core_KE_new_sboxw_29_), .Y(n6361) );
  INVX1 U17563 ( .A(top_core_KE_new_sboxw_26_), .Y(n6369) );
  NOR2X1 U17564 ( .A(n11674), .B(n11778), .Y(n11839) );
  NOR2X1 U17565 ( .A(top_core_KE_sb1_n99), .B(top_core_KE_sb1_n206), .Y(
        top_core_KE_sb1_n268) );
  NOR2X1 U17566 ( .A(n12305), .B(n12409), .Y(n12470) );
  NOR2X1 U17567 ( .A(n13251), .B(n13355), .Y(n13415) );
  NOR2X1 U17568 ( .A(n11990), .B(n12094), .Y(n12155) );
  NOR2X1 U17569 ( .A(n12621), .B(n12725), .Y(n12785) );
  NOR2X1 U17570 ( .A(n13566), .B(n13670), .Y(n13730) );
  NOR2X1 U17571 ( .A(n12936), .B(n13040), .Y(n13100) );
  NOR3XL U17572 ( .A(top_core_KE_n1865), .B(top_core_KE_N1), .C(
        top_core_KE_n2704), .Y(top_core_KE_n1870) );
  NOR2X1 U17573 ( .A(n685), .B(n1647), .Y(n13601) );
  OAI222XL U17574 ( .A0(n11718), .A1(n11717), .B0(n11852), .B1(n1815), .C0(
        n11779), .C1(n11651), .Y(n11850) );
  OAI222XL U17575 ( .A0(top_core_KE_sb1_n145), .A1(top_core_KE_sb1_n144), .B0(
        top_core_KE_sb1_n281), .B1(n1836), .C0(top_core_KE_sb1_n207), .C1(
        top_core_KE_sb1_n76), .Y(top_core_KE_sb1_n279) );
  OAI222XL U17576 ( .A0(n12349), .A1(n12348), .B0(n12483), .B1(n1771), .C0(
        n12410), .C1(n12283), .Y(n12481) );
  OAI222XL U17577 ( .A0(n13295), .A1(n13294), .B0(n13428), .B1(n1692), .C0(n3), 
        .C1(n13228), .Y(n13426) );
  OAI222XL U17578 ( .A0(n12034), .A1(n12033), .B0(n12168), .B1(n1794), .C0(
        n12095), .C1(n11967), .Y(n12166) );
  OAI222XL U17579 ( .A0(n12665), .A1(n12664), .B0(n12798), .B1(n1748), .C0(n4), 
        .C1(n12598), .Y(n12796) );
  OAI222XL U17580 ( .A0(n13610), .A1(n13609), .B0(n13743), .B1(n1662), .C0(n6), 
        .C1(n13543), .Y(n13741) );
  OAI222XL U17581 ( .A0(n12980), .A1(n12979), .B0(n13113), .B1(n1719), .C0(n5), 
        .C1(n12913), .Y(n13111) );
  NOR2X1 U17582 ( .A(top_core_KE_N1), .B(top_core_KE_N0), .Y(top_core_KE_n2704) );
  NOR3XL U17583 ( .A(n11735), .B(n1799), .C(n50), .Y(n11833) );
  NOR3XL U17584 ( .A(top_core_KE_sb1_n162), .B(n1820), .C(n51), .Y(
        top_core_KE_sb1_n262) );
  NOR3XL U17585 ( .A(n12366), .B(n1756), .C(n89), .Y(n12464) );
  NOR3XL U17586 ( .A(n12051), .B(n1778), .C(n53), .Y(n12149) );
  NOR3XL U17587 ( .A(n13627), .B(n1638), .C(n55), .Y(n13724) );
  NOR2X1 U17588 ( .A(n7007), .B(n7016), .Y(top_core_KE_n884) );
  OAI222XL U17589 ( .A0(n11812), .A1(n1796), .B0(n11813), .B1(n11679), .C0(
        top_core_KE_prev_key1_reg_13_), .C1(n11814), .Y(n11801) );
  AOI211X1 U17590 ( .A0(n6909), .A1(n1808), .B0(n11815), .C0(n11816), .Y(
        n11814) );
  AOI221X1 U17591 ( .A0(n6917), .A1(n689), .B0(n1221), .B1(n761), .C0(n11818), 
        .Y(n11812) );
  OAI222XL U17592 ( .A0(top_core_KE_sb1_n240), .A1(n1817), .B0(
        top_core_KE_sb1_n241), .B1(top_core_KE_sb1_n104), .C0(
        top_core_KE_prev_key1_reg_5_), .C1(top_core_KE_sb1_n242), .Y(
        top_core_KE_sb1_n229) );
  AOI211X1 U17593 ( .A0(n6863), .A1(n1829), .B0(top_core_KE_sb1_n243), .C0(
        top_core_KE_sb1_n244), .Y(top_core_KE_sb1_n242) );
  AOI221X1 U17594 ( .A0(n6871), .A1(n690), .B0(n1215), .B1(n762), .C0(
        top_core_KE_sb1_n246), .Y(top_core_KE_sb1_n240) );
  OAI222XL U17595 ( .A0(n12443), .A1(n1753), .B0(n12444), .B1(n12310), .C0(
        n1757), .C1(n12445), .Y(n12432) );
  AOI211X1 U17596 ( .A0(n6616), .A1(n1766), .B0(n12446), .C0(n12447), .Y(
        n12445) );
  AOI221X1 U17597 ( .A0(n6624), .A1(n691), .B0(n1183), .B1(n760), .C0(n12449), 
        .Y(n12443) );
  OAI222XL U17598 ( .A0(n12128), .A1(n1775), .B0(n12129), .B1(n11995), .C0(
        top_core_KE_prev_key1_reg_21_), .C1(n12130), .Y(n12117) );
  AOI211X1 U17599 ( .A0(n6569), .A1(n1787), .B0(n12131), .C0(n12132), .Y(
        n12130) );
  AOI221X1 U17600 ( .A0(n6577), .A1(n693), .B0(n1175), .B1(n763), .C0(n12134), 
        .Y(n12128) );
  OAI222XL U17601 ( .A0(n13703), .A1(n1635), .B0(n13704), .B1(n13571), .C0(
        n1639), .C1(n13705), .Y(n13692) );
  AOI211X1 U17602 ( .A0(n6592), .A1(n1657), .B0(n13706), .C0(n13707), .Y(
        n13705) );
  AOI221X1 U17603 ( .A0(n6600), .A1(n695), .B0(n1180), .B1(n759), .C0(n13709), 
        .Y(n13703) );
  NOR2X1 U17604 ( .A(n681), .B(n1798), .Y(n11654) );
  NOR2X1 U17605 ( .A(n682), .B(n1819), .Y(top_core_KE_sb1_n79) );
  NOR2X1 U17606 ( .A(n683), .B(top_core_KE_prev_key1_reg_29_), .Y(n12286) );
  NOR2X1 U17607 ( .A(n684), .B(n1777), .Y(n11970) );
  NOR2X1 U17608 ( .A(n669), .B(n1640), .Y(n13546) );
  OAI221XL U17609 ( .A0(n11778), .A1(n11651), .B0(n1810), .B1(n50), .C0(n11773), .Y(n11942) );
  OAI221XL U17610 ( .A0(top_core_KE_sb1_n206), .A1(top_core_KE_sb1_n76), .B0(
        n1831), .B1(n51), .C0(top_core_KE_sb1_n201), .Y(top_core_KE_sb1_n372)
         );
  OAI221XL U17611 ( .A0(n12409), .A1(n12283), .B0(n1768), .B1(n89), .C0(n12404), .Y(n12573) );
  OAI221XL U17612 ( .A0(n12094), .A1(n11967), .B0(n1789), .B1(n53), .C0(n12089), .Y(n12258) );
  OAI222XL U17613 ( .A0(n11674), .A1(n11672), .B0(n1800), .B1(n11686), .C0(
        n11687), .C1(n1795), .Y(n11682) );
  AND3X2 U17614 ( .A(n11688), .B(n11689), .C(n11690), .Y(n11687) );
  OAI222XL U17615 ( .A0(top_core_KE_sb1_n99), .A1(top_core_KE_sb1_n97), .B0(
        n1821), .B1(top_core_KE_sb1_n111), .C0(top_core_KE_sb1_n112), .C1(
        n1816), .Y(top_core_KE_sb1_n107) );
  AND3X2 U17616 ( .A(top_core_KE_sb1_n113), .B(top_core_KE_sb1_n114), .C(
        top_core_KE_sb1_n115), .Y(top_core_KE_sb1_n112) );
  OAI222XL U17617 ( .A0(n12305), .A1(n12303), .B0(n1757), .B1(n12317), .C0(
        n12318), .C1(n1752), .Y(n12313) );
  AND3X2 U17618 ( .A(n12319), .B(n12320), .C(n12321), .Y(n12318) );
  OAI222XL U17619 ( .A0(n13251), .A1(n13249), .B0(n1667), .B1(n13263), .C0(
        n13264), .C1(n1672), .Y(n13259) );
  AND3X2 U17620 ( .A(n13265), .B(n13266), .C(n13267), .Y(n13264) );
  OAI222XL U17621 ( .A0(n11990), .A1(n11988), .B0(n1779), .B1(n12002), .C0(
        n12003), .C1(n1774), .Y(n11998) );
  AND3X2 U17622 ( .A(n12004), .B(n12005), .C(n12006), .Y(n12003) );
  OAI222XL U17623 ( .A0(n12936), .A1(n12934), .B0(n1696), .B1(n12948), .C0(
        n12949), .C1(n1701), .Y(n12944) );
  AND3X2 U17624 ( .A(n12950), .B(n12951), .C(n12952), .Y(n12949) );
  OAI222XL U17625 ( .A0(n13566), .A1(n13564), .B0(n1640), .B1(n13578), .C0(
        n13579), .C1(n1635), .Y(n13574) );
  AND3X2 U17626 ( .A(n13580), .B(n13581), .C(n13582), .Y(n13579) );
  OAI222XL U17627 ( .A0(n12621), .A1(n12619), .B0(n1725), .B1(n12633), .C0(
        n12634), .C1(n1730), .Y(n12629) );
  AND3X2 U17628 ( .A(n12635), .B(n12636), .C(n12637), .Y(n12634) );
  NOR2XL U17629 ( .A(n11779), .B(n577), .Y(n11764) );
  NOR2XL U17630 ( .A(top_core_KE_sb1_n207), .B(n578), .Y(top_core_KE_sb1_n192)
         );
  NOR2XL U17631 ( .A(n12410), .B(n579), .Y(n12395) );
  NOR2XL U17632 ( .A(n12095), .B(n581), .Y(n12080) );
  NAND2X1 U17633 ( .A(n6622), .B(n1171), .Y(n12290) );
  AOI32XL U17634 ( .A0(n13355), .A1(n1679), .A2(n686), .B0(n13373), .B1(n1172), 
        .Y(n13445) );
  NAND2X1 U17635 ( .A(n3447), .B(n1506), .Y(n13837) );
  NAND2X1 U17636 ( .A(n2846), .B(n1504), .Y(n16987) );
  NAND2X1 U17637 ( .A(n2604), .B(n1528), .Y(n18247) );
  NAND2X1 U17638 ( .A(n3206), .B(n1518), .Y(n15097) );
  NAND2X1 U17639 ( .A(n3145), .B(n1515), .Y(n15412) );
  NAND2X1 U17640 ( .A(n2907), .B(n1507), .Y(n16672) );
  NAND2X1 U17641 ( .A(n2543), .B(n1525), .Y(n18562) );
  NAND2X1 U17642 ( .A(n3267), .B(n1520), .Y(n14782) );
  NAND2X1 U17643 ( .A(n2968), .B(n1509), .Y(n16357) );
  NAND2X1 U17644 ( .A(n2665), .B(n1530), .Y(n17932) );
  NAND2X1 U17645 ( .A(n3328), .B(n1522), .Y(n14467) );
  NAND2X1 U17646 ( .A(n3026), .B(n1511), .Y(n16042) );
  NAND2X1 U17647 ( .A(n2725), .B(n1532), .Y(n17617) );
  NAND2X1 U17648 ( .A(n3386), .B(n1524), .Y(n14152) );
  NAND2X1 U17649 ( .A(n3087), .B(n1513), .Y(n15727) );
  NAND2X1 U17650 ( .A(n2786), .B(n1502), .Y(n17302) );
  NAND2X1 U17651 ( .A(n752), .B(n1171), .Y(n12437) );
  OAI221XL U17652 ( .A0(n1799), .A1(n11940), .B0(n11691), .B1(n11852), .C0(
        n11941), .Y(n11932) );
  AOI21X1 U17653 ( .A0(n6826), .A1(n11942), .B0(n11943), .Y(n11941) );
  OAI32X1 U17654 ( .A0(n1211), .A1(n11944), .A2(n1796), .B0(n1221), .B1(n11675), .Y(n11943) );
  OAI221XL U17655 ( .A0(n1820), .A1(top_core_KE_sb1_n370), .B0(
        top_core_KE_sb1_n116), .B1(top_core_KE_sb1_n281), .C0(
        top_core_KE_sb1_n371), .Y(top_core_KE_sb1_n361) );
  AOI21X1 U17656 ( .A0(n6804), .A1(top_core_KE_sb1_n372), .B0(
        top_core_KE_sb1_n373), .Y(top_core_KE_sb1_n371) );
  OAI32X1 U17657 ( .A0(n1210), .A1(top_core_KE_sb1_n374), .A2(n1817), .B0(
        n1215), .B1(top_core_KE_sb1_n100), .Y(top_core_KE_sb1_n373) );
  OAI221XL U17658 ( .A0(n1757), .A1(n12571), .B0(n12322), .B1(n12483), .C0(
        n12572), .Y(n12563) );
  AOI21X1 U17659 ( .A0(n6530), .A1(n12573), .B0(n12574), .Y(n12572) );
  OAI32X1 U17660 ( .A0(n1171), .A1(n12575), .A2(n1753), .B0(n1183), .B1(n12306), .Y(n12574) );
  OAI221XL U17661 ( .A0(n1778), .A1(n12256), .B0(n12007), .B1(n12168), .C0(
        n12257), .Y(n12248) );
  AOI21X1 U17662 ( .A0(n6507), .A1(n12258), .B0(n12259), .Y(n12257) );
  OAI32X1 U17663 ( .A0(n1170), .A1(n12260), .A2(n1775), .B0(n1175), .B1(n11991), .Y(n12259) );
  OAI221XL U17664 ( .A0(n1639), .A1(n13831), .B0(n13583), .B1(n13743), .C0(
        n13832), .Y(n13823) );
  AOI21X1 U17665 ( .A0(n6519), .A1(n13833), .B0(n13834), .Y(n13832) );
  OAI32X1 U17666 ( .A0(n1644), .A1(n13835), .A2(n1636), .B0(n1180), .B1(n13567), .Y(n13834) );
  OAI211X1 U17667 ( .A0(n1222), .A1(n11919), .B0(n11920), .C0(n11921), .Y(
        n11918) );
  AOI31XL U17668 ( .A0(n1222), .A1(n11769), .A2(n11652), .B0(n6828), .Y(n11920) );
  NAND4X1 U17669 ( .A(n11884), .B(n11808), .C(n11923), .D(n11924), .Y(n11922)
         );
  OAI211X1 U17670 ( .A0(n1216), .A1(top_core_KE_sb1_n348), .B0(
        top_core_KE_sb1_n349), .C0(top_core_KE_sb1_n350), .Y(
        top_core_KE_sb1_n347) );
  AOI31XL U17671 ( .A0(n1216), .A1(top_core_KE_sb1_n197), .A2(
        top_core_KE_sb1_n77), .B0(n6806), .Y(top_core_KE_sb1_n349) );
  NAND4X1 U17672 ( .A(top_core_KE_sb1_n313), .B(top_core_KE_sb1_n236), .C(
        top_core_KE_sb1_n352), .D(top_core_KE_sb1_n353), .Y(
        top_core_KE_sb1_n351) );
  OAI211X1 U17673 ( .A0(n1181), .A1(n12550), .B0(n12551), .C0(n12552), .Y(
        n12549) );
  AOI31XL U17674 ( .A0(n1181), .A1(n12400), .A2(n12284), .B0(n6532), .Y(n12551) );
  NAND4X1 U17675 ( .A(n12515), .B(n12439), .C(n12554), .D(n12555), .Y(n12553)
         );
  OAI211X1 U17676 ( .A0(n1176), .A1(n12235), .B0(n12236), .C0(n12237), .Y(
        n12234) );
  AOI31XL U17677 ( .A0(n1176), .A1(n12085), .A2(n11968), .B0(n6509), .Y(n12236) );
  NAND4X1 U17678 ( .A(n12200), .B(n12124), .C(n12239), .D(n12240), .Y(n12238)
         );
  OAI211X1 U17679 ( .A0(n1178), .A1(n13810), .B0(n13811), .C0(n13812), .Y(
        n13809) );
  AOI31XL U17680 ( .A0(n1178), .A1(n13661), .A2(n13544), .B0(n6521), .Y(n13811) );
  NAND4X1 U17681 ( .A(n13775), .B(n13699), .C(n13814), .D(n13815), .Y(n13813)
         );
  NOR2X1 U17682 ( .A(n1845), .B(n7019), .Y(top_core_KE_n2506) );
  NAND2X1 U17683 ( .A(n1506), .B(n3451), .Y(n13839) );
  NAND2X1 U17684 ( .A(n1504), .B(n2850), .Y(n16989) );
  NAND2X1 U17685 ( .A(n1528), .B(n2608), .Y(n18249) );
  NAND2X1 U17686 ( .A(n1518), .B(n3210), .Y(n15099) );
  NAND2X1 U17687 ( .A(n1515), .B(n3149), .Y(n15414) );
  NAND2X1 U17688 ( .A(n1507), .B(n2911), .Y(n16674) );
  NAND2X1 U17689 ( .A(n1525), .B(n2547), .Y(n18564) );
  NAND2X1 U17690 ( .A(n1520), .B(n3271), .Y(n14784) );
  NAND2X1 U17691 ( .A(n1509), .B(n2972), .Y(n16359) );
  NAND2X1 U17692 ( .A(n1530), .B(n2669), .Y(n17934) );
  NAND2X1 U17693 ( .A(n1522), .B(n3332), .Y(n14469) );
  NAND2X1 U17694 ( .A(n1511), .B(n3030), .Y(n16044) );
  NAND2X1 U17695 ( .A(n1532), .B(n2729), .Y(n17619) );
  NAND2X1 U17696 ( .A(n1524), .B(n3390), .Y(n14154) );
  NAND2X1 U17697 ( .A(n1513), .B(n3091), .Y(n15729) );
  NAND2X1 U17698 ( .A(n1502), .B(n2790), .Y(n17304) );
  NAND2X1 U17699 ( .A(n151), .B(n1500), .Y(top_core_KE_n2710) );
  AOI31X1 U17700 ( .A0(n11669), .A1(n11670), .A2(n11671), .B0(n1801), .Y(
        n11668) );
  AOI31X1 U17701 ( .A0(top_core_KE_sb1_n94), .A1(top_core_KE_sb1_n95), .A2(
        top_core_KE_sb1_n96), .B0(n1822), .Y(top_core_KE_sb1_n93) );
  AOI31X1 U17702 ( .A0(n12300), .A1(n12301), .A2(n12302), .B0(n1754), .Y(
        n12299) );
  AOI31X1 U17703 ( .A0(n11985), .A1(n11986), .A2(n11987), .B0(n1780), .Y(
        n11984) );
  OAI221XL U17704 ( .A0(n513), .A1(n2870), .B0(n2867), .B1(n2893), .C0(n1505), 
        .Y(n17107) );
  OAI221XL U17705 ( .A0(n514), .A1(n3471), .B0(n3468), .B1(n3494), .C0(n1517), 
        .Y(n13957) );
  OAI221XL U17706 ( .A0(n515), .A1(n2628), .B0(n2625), .B1(n2650), .C0(n1529), 
        .Y(n18367) );
  OAI221XL U17707 ( .A0(n516), .A1(n3230), .B0(n3227), .B1(n3253), .C0(n1519), 
        .Y(n15217) );
  OAI221XL U17708 ( .A0(n517), .A1(n3169), .B0(n3166), .B1(n3192), .C0(n1516), 
        .Y(n15532) );
  OAI221XL U17709 ( .A0(n518), .A1(n2567), .B0(n2564), .B1(n2590), .C0(n1526), 
        .Y(n18682) );
  OAI221XL U17710 ( .A0(n519), .A1(n2931), .B0(n2928), .B1(n2954), .C0(n1508), 
        .Y(n16792) );
  OAI221XL U17711 ( .A0(n520), .A1(n3291), .B0(n3288), .B1(n3314), .C0(n1521), 
        .Y(n14902) );
  OAI221XL U17712 ( .A0(n521), .A1(n2992), .B0(n2989), .B1(n3015), .C0(n1510), 
        .Y(n16477) );
  OAI221XL U17713 ( .A0(n522), .A1(n2689), .B0(n2686), .B1(n2711), .C0(n1531), 
        .Y(n18052) );
  OAI221XL U17714 ( .A0(n523), .A1(n3352), .B0(n3349), .B1(n3375), .C0(n1523), 
        .Y(n14587) );
  OAI221XL U17715 ( .A0(n524), .A1(n3050), .B0(n3047), .B1(n3072), .C0(n1512), 
        .Y(n16162) );
  OAI221XL U17716 ( .A0(n525), .A1(n2747), .B0(n2746), .B1(n2772), .C0(n1501), 
        .Y(n17737) );
  OAI221XL U17717 ( .A0(n526), .A1(n3410), .B0(n3407), .B1(n3433), .C0(n1527), 
        .Y(n14272) );
  OAI221XL U17718 ( .A0(n527), .A1(n3111), .B0(n3108), .B1(n3134), .C0(n1514), 
        .Y(n15847) );
  OAI221XL U17719 ( .A0(n528), .A1(n2810), .B0(n2807), .B1(n2833), .C0(n1503), 
        .Y(n17422) );
  OAI221XL U17720 ( .A0(n6540), .A1(n1665), .B0(n1667), .B1(n13287), .C0(
        n13288), .Y(n13271) );
  INVX1 U17721 ( .A(n13296), .Y(n6540) );
  AOI22X1 U17722 ( .A0(n6476), .A1(n1174), .B0(n677), .B1(n13289), .Y(n13288)
         );
  OAI221XL U17723 ( .A0(n6835), .A1(n1723), .B0(n1725), .B1(n12657), .C0(
        n12658), .Y(n12641) );
  INVX1 U17724 ( .A(n12666), .Y(n6835) );
  AOI22X1 U17725 ( .A0(n6779), .A1(n1214), .B0(n678), .B1(n12659), .Y(n12658)
         );
  OAI221XL U17726 ( .A0(n6881), .A1(n1694), .B0(n1696), .B1(n12972), .C0(
        n12973), .Y(n12956) );
  INVX1 U17727 ( .A(n12981), .Y(n6881) );
  AOI22X1 U17728 ( .A0(n6818), .A1(n1220), .B0(n680), .B1(n12974), .Y(n12973)
         );
  OAI221XL U17729 ( .A0(n6905), .A1(n1796), .B0(n1799), .B1(n11710), .C0(
        n11711), .Y(n11694) );
  INVX1 U17730 ( .A(n11719), .Y(n6905) );
  AOI22X1 U17731 ( .A0(n6829), .A1(n613), .B0(n673), .B1(n11712), .Y(n11711)
         );
  OAI221XL U17732 ( .A0(n6859), .A1(n1817), .B0(n1820), .B1(
        top_core_KE_sb1_n136), .C0(top_core_KE_sb1_n137), .Y(
        top_core_KE_sb1_n119) );
  INVX1 U17733 ( .A(top_core_KE_sb1_n146), .Y(n6859) );
  AOI22X1 U17734 ( .A0(n6808), .A1(n614), .B0(n674), .B1(top_core_KE_sb1_n138), 
        .Y(top_core_KE_sb1_n137) );
  OAI221XL U17735 ( .A0(n6612), .A1(n1753), .B0(n1754), .B1(n12341), .C0(
        n12342), .Y(n12325) );
  INVX1 U17736 ( .A(n12350), .Y(n6612) );
  AOI22X1 U17737 ( .A0(n6533), .A1(n601), .B0(n675), .B1(n12343), .Y(n12342)
         );
  OAI221XL U17738 ( .A0(n6565), .A1(n1775), .B0(n1778), .B1(n12026), .C0(
        n12027), .Y(n12010) );
  INVX1 U17739 ( .A(n12035), .Y(n6565) );
  AOI22X1 U17740 ( .A0(n6511), .A1(n615), .B0(n676), .B1(n12028), .Y(n12027)
         );
  OAI221XL U17741 ( .A0(n6588), .A1(n1636), .B0(n1640), .B1(n13602), .C0(
        n13603), .Y(n13586) );
  INVX1 U17742 ( .A(n13611), .Y(n6588) );
  AOI22X1 U17743 ( .A0(n6522), .A1(n1179), .B0(n679), .B1(n13604), .Y(n13603)
         );
  OAI22XL U17744 ( .A0(n1209), .A1(n1804), .B0(n1802), .B1(n11778), .Y(n11798)
         );
  OAI22XL U17745 ( .A0(n1207), .A1(n1825), .B0(n1823), .B1(
        top_core_KE_sb1_n206), .Y(top_core_KE_sb1_n226) );
  OAI22XL U17746 ( .A0(n1169), .A1(n1765), .B0(n1760), .B1(n12409), .Y(n12429)
         );
  OAI22XL U17747 ( .A0(n1167), .A1(n1783), .B0(n1781), .B1(n12094), .Y(n12114)
         );
  OAI22XL U17748 ( .A0(n1168), .A1(n1656), .B0(n1651), .B1(n13670), .Y(n13689)
         );
  OAI22XL U17749 ( .A0(n1166), .A1(n1686), .B0(n1680), .B1(n13355), .Y(n13374)
         );
  OAI22XL U17750 ( .A0(n1206), .A1(n1744), .B0(n1738), .B1(n12725), .Y(n12744)
         );
  OAI22XL U17751 ( .A0(n1208), .A1(n1715), .B0(n1709), .B1(n13040), .Y(n13059)
         );
  AOI21X1 U17752 ( .A0(n6587), .A1(n631), .B0(n13696), .Y(n13695) );
  AOI31X1 U17753 ( .A0(n6826), .A1(n1209), .A2(n665), .B0(n6825), .Y(n11936)
         );
  AOI31X1 U17754 ( .A0(n6804), .A1(n1207), .A2(n666), .B0(n6803), .Y(
        top_core_KE_sb1_n365) );
  AOI31X1 U17755 ( .A0(n6530), .A1(n1169), .A2(n667), .B0(n6529), .Y(n12567)
         );
  AOI31X1 U17756 ( .A0(n6507), .A1(n1167), .A2(n668), .B0(n6506), .Y(n12252)
         );
  AOI31X1 U17757 ( .A0(n6775), .A1(n1206), .A2(n688), .B0(n6774), .Y(n12882)
         );
  AOI31X1 U17758 ( .A0(n6519), .A1(n1168), .A2(n685), .B0(n6518), .Y(n13827)
         );
  AOI31X1 U17759 ( .A0(n6815), .A1(n1208), .A2(n687), .B0(n6814), .Y(n13197)
         );
  NOR4BX1 U17760 ( .AN(n11937), .B(n11938), .C(n6920), .D(n11681), .Y(n11935)
         );
  OAI221XL U17761 ( .A0(n1221), .A1(n11852), .B0(n1815), .B1(n80), .C0(n11939), 
        .Y(n11938) );
  AOI22X1 U17762 ( .A0(n689), .A1(n745), .B0(n6914), .B1(n1804), .Y(n11939) );
  NOR4BX1 U17763 ( .AN(top_core_KE_sb1_n366), .B(top_core_KE_sb1_n367), .C(
        n6874), .D(top_core_KE_sb1_n106), .Y(top_core_KE_sb1_n364) );
  OAI221XL U17764 ( .A0(n1215), .A1(top_core_KE_sb1_n281), .B0(n1836), .B1(n81), .C0(top_core_KE_sb1_n368), .Y(top_core_KE_sb1_n367) );
  AOI22X1 U17765 ( .A0(n690), .A1(n746), .B0(n6868), .B1(n1825), .Y(
        top_core_KE_sb1_n368) );
  NOR4BX1 U17766 ( .AN(n12568), .B(n12569), .C(n6627), .D(n12312), .Y(n12566)
         );
  OAI221XL U17767 ( .A0(n1183), .A1(n12483), .B0(n1770), .B1(n82), .C0(n12570), 
        .Y(n12569) );
  AOI22X1 U17768 ( .A0(n691), .A1(n744), .B0(n6621), .B1(n1763), .Y(n12570) );
  NOR4BX1 U17769 ( .AN(n12253), .B(n12254), .C(n6580), .D(n11997), .Y(n12251)
         );
  OAI221XL U17770 ( .A0(n1175), .A1(n12168), .B0(n1794), .B1(n83), .C0(n12255), 
        .Y(n12254) );
  AOI22X1 U17771 ( .A0(n693), .A1(n747), .B0(n6574), .B1(n1783), .Y(n12255) );
  INVX1 U17772 ( .A(top_core_KE_new_sboxw_14_), .Y(n6721) );
  INVX1 U17773 ( .A(top_core_KE_new_sboxw_8_), .Y(n6739) );
  INVX1 U17774 ( .A(top_core_KE_new_sboxw_6_), .Y(n6786) );
  INVX1 U17775 ( .A(top_core_KE_new_sboxw_0_), .Y(n6797) );
  INVX1 U17776 ( .A(top_core_KE_new_sboxw_30_), .Y(n6347) );
  INVX1 U17777 ( .A(top_core_KE_new_sboxw_24_), .Y(n6355) );
  INVX1 U17778 ( .A(top_core_KE_new_sboxw_9_), .Y(n6736) );
  INVX1 U17779 ( .A(top_core_KE_new_sboxw_1_), .Y(n6795) );
  INVX1 U17780 ( .A(top_core_KE_new_sboxw_25_), .Y(n6374) );
  INVX1 U17781 ( .A(top_core_KE_new_sboxw_12_), .Y(n6725) );
  INVX1 U17782 ( .A(top_core_KE_new_sboxw_11_), .Y(n6732) );
  INVX1 U17783 ( .A(top_core_KE_new_sboxw_4_), .Y(n6788) );
  INVX1 U17784 ( .A(top_core_KE_new_sboxw_3_), .Y(n6790) );
  AOI31XL U17785 ( .A0(n11742), .A1(n185), .A2(n11686), .B0(n11679), .Y(n11761) );
  AOI31XL U17786 ( .A0(top_core_KE_sb1_n169), .A1(n186), .A2(
        top_core_KE_sb1_n111), .B0(top_core_KE_sb1_n104), .Y(
        top_core_KE_sb1_n189) );
  AOI31XL U17787 ( .A0(n12373), .A1(n46), .A2(n12317), .B0(n12310), .Y(n12392)
         );
  AOI31XL U17788 ( .A0(n13319), .A1(n187), .A2(n13263), .B0(n13256), .Y(n13338) );
  AOI31XL U17789 ( .A0(n12058), .A1(n188), .A2(n12002), .B0(n11995), .Y(n12077) );
  AOI31XL U17790 ( .A0(n12689), .A1(n189), .A2(n12633), .B0(n12626), .Y(n12708) );
  AOI31XL U17791 ( .A0(n13634), .A1(n190), .A2(n13578), .B0(n13571), .Y(n13653) );
  AOI31XL U17792 ( .A0(n13004), .A1(n191), .A2(n12948), .B0(n12941), .Y(n13023) );
  INVX1 U17793 ( .A(top_core_KE_new_sboxw_28_), .Y(n6351) );
  INVX1 U17794 ( .A(top_core_KE_new_sboxw_27_), .Y(n6365) );
  INVX1 U17795 ( .A(top_core_KE_n2517), .Y(n6485) );
  INVX1 U17796 ( .A(top_core_KE_n2526), .Y(n6492) );
  INVX1 U17797 ( .A(top_core_KE_n2514), .Y(n6484) );
  INVX1 U17798 ( .A(top_core_KE_n2532), .Y(n6499) );
  INVX1 U17799 ( .A(top_core_KE_n2520), .Y(n6486) );
  INVX1 U17800 ( .A(top_core_KE_n2523), .Y(n6489) );
  INVX1 U17801 ( .A(top_core_KE_n2529), .Y(n6496) );
  NOR2XL U17802 ( .A(n77), .B(n1809), .Y(n11879) );
  NOR2XL U17803 ( .A(n78), .B(n1830), .Y(top_core_KE_sb1_n308) );
  NOR2XL U17804 ( .A(n184), .B(n1767), .Y(n12510) );
  NOR2XL U17805 ( .A(n79), .B(n1788), .Y(n12195) );
  NAND2X1 U17806 ( .A(n1144), .B(n1517), .Y(n13949) );
  NAND2X1 U17807 ( .A(n1005), .B(n1505), .Y(n17099) );
  NAND2X1 U17808 ( .A(n1089), .B(n1519), .Y(n15209) );
  NAND2X1 U17809 ( .A(n949), .B(n1529), .Y(n18359) );
  NAND2X1 U17810 ( .A(n1075), .B(n1516), .Y(n15524) );
  NAND2X1 U17811 ( .A(n935), .B(n1526), .Y(n18674) );
  NAND2X1 U17812 ( .A(n1019), .B(n1508), .Y(n16784) );
  NAND2X1 U17813 ( .A(n1103), .B(n1521), .Y(n14894) );
  NAND2X1 U17814 ( .A(n1033), .B(n1510), .Y(n16469) );
  NAND2X1 U17815 ( .A(n963), .B(n1531), .Y(n18044) );
  NAND2X1 U17816 ( .A(n1117), .B(n1523), .Y(n14579) );
  NAND2X1 U17817 ( .A(n1047), .B(n1512), .Y(n16154) );
  NAND2X1 U17818 ( .A(n977), .B(n1501), .Y(n17729) );
  NAND2X1 U17819 ( .A(n1131), .B(n1527), .Y(n14264) );
  NAND2X1 U17820 ( .A(n1061), .B(n1514), .Y(n15839) );
  NAND2X1 U17821 ( .A(n991), .B(n1503), .Y(n17414) );
  AOI211X1 U17822 ( .A0(n17008), .A1(n17096), .B0(n17097), .C0(n17098), .Y(
        n17095) );
  AOI22X1 U17823 ( .A0(n2854), .A1(n17100), .B0(n17101), .B1(n2851), .Y(n17094) );
  OAI21XL U17824 ( .A0(n2866), .A1(n450), .B0(n1505), .Y(n17096) );
  AOI211X1 U17825 ( .A0(n13858), .A1(n13946), .B0(n13947), .C0(n13948), .Y(
        n13945) );
  AOI22X1 U17826 ( .A0(n3455), .A1(n13950), .B0(n13951), .B1(n3452), .Y(n13944) );
  OAI21XL U17827 ( .A0(n3467), .A1(n449), .B0(n1517), .Y(n13946) );
  AOI211X1 U17828 ( .A0(n18268), .A1(n18356), .B0(n18357), .C0(n18358), .Y(
        n18355) );
  AOI22X1 U17829 ( .A0(n2612), .A1(n18360), .B0(n18361), .B1(n2609), .Y(n18354) );
  OAI21XL U17830 ( .A0(n2624), .A1(n451), .B0(n1529), .Y(n18356) );
  AOI211X1 U17831 ( .A0(n15118), .A1(n15206), .B0(n15207), .C0(n15208), .Y(
        n15205) );
  AOI22X1 U17832 ( .A0(n3214), .A1(n15210), .B0(n15211), .B1(n3211), .Y(n15204) );
  OAI21XL U17833 ( .A0(n3226), .A1(n452), .B0(n1519), .Y(n15206) );
  AOI211X1 U17834 ( .A0(n15433), .A1(n15521), .B0(n15522), .C0(n15523), .Y(
        n15520) );
  AOI22X1 U17835 ( .A0(n3153), .A1(n15525), .B0(n15526), .B1(n3150), .Y(n15519) );
  OAI21XL U17836 ( .A0(n3165), .A1(n453), .B0(n1516), .Y(n15521) );
  AOI211X1 U17837 ( .A0(n18583), .A1(n18671), .B0(n18672), .C0(n18673), .Y(
        n18670) );
  AOI22X1 U17838 ( .A0(n2551), .A1(n18675), .B0(n18676), .B1(n2548), .Y(n18669) );
  OAI21XL U17839 ( .A0(n2563), .A1(n454), .B0(n1526), .Y(n18671) );
  AOI211X1 U17840 ( .A0(n16693), .A1(n16781), .B0(n16782), .C0(n16783), .Y(
        n16780) );
  AOI22X1 U17841 ( .A0(n2915), .A1(n16785), .B0(n16786), .B1(n2912), .Y(n16779) );
  OAI21XL U17842 ( .A0(n2927), .A1(n455), .B0(n1508), .Y(n16781) );
  AOI211X1 U17843 ( .A0(n14803), .A1(n14891), .B0(n14892), .C0(n14893), .Y(
        n14890) );
  AOI22X1 U17844 ( .A0(n3275), .A1(n14895), .B0(n14896), .B1(n3272), .Y(n14889) );
  OAI21XL U17845 ( .A0(n3287), .A1(n456), .B0(n1521), .Y(n14891) );
  AOI211X1 U17846 ( .A0(n16378), .A1(n16466), .B0(n16467), .C0(n16468), .Y(
        n16465) );
  AOI22X1 U17847 ( .A0(n2976), .A1(n16470), .B0(n16471), .B1(n2973), .Y(n16464) );
  OAI21XL U17848 ( .A0(n2988), .A1(n457), .B0(n1510), .Y(n16466) );
  AOI211X1 U17849 ( .A0(n17953), .A1(n18041), .B0(n18042), .C0(n18043), .Y(
        n18040) );
  AOI22X1 U17850 ( .A0(n2673), .A1(n18045), .B0(n18046), .B1(n2670), .Y(n18039) );
  OAI21XL U17851 ( .A0(n2685), .A1(n458), .B0(n1531), .Y(n18041) );
  AOI211X1 U17852 ( .A0(n14488), .A1(n14576), .B0(n14577), .C0(n14578), .Y(
        n14575) );
  AOI22X1 U17853 ( .A0(n3336), .A1(n14580), .B0(n14581), .B1(n3333), .Y(n14574) );
  OAI21XL U17854 ( .A0(n3348), .A1(n459), .B0(n1523), .Y(n14576) );
  AOI211X1 U17855 ( .A0(n16063), .A1(n16151), .B0(n16152), .C0(n16153), .Y(
        n16150) );
  AOI22X1 U17856 ( .A0(n3034), .A1(n16155), .B0(n16156), .B1(n3031), .Y(n16149) );
  OAI21XL U17857 ( .A0(n3046), .A1(n460), .B0(n1512), .Y(n16151) );
  AOI211X1 U17858 ( .A0(n17638), .A1(n17726), .B0(n17727), .C0(n17728), .Y(
        n17725) );
  AOI22X1 U17859 ( .A0(n2733), .A1(n17730), .B0(n17731), .B1(n2730), .Y(n17724) );
  OAI21XL U17860 ( .A0(n2745), .A1(n461), .B0(n1501), .Y(n17726) );
  AOI211X1 U17861 ( .A0(n14173), .A1(n14261), .B0(n14262), .C0(n14263), .Y(
        n14260) );
  AOI22X1 U17862 ( .A0(n3394), .A1(n14265), .B0(n14266), .B1(n3391), .Y(n14259) );
  OAI21XL U17863 ( .A0(n3406), .A1(n462), .B0(n1527), .Y(n14261) );
  AOI211X1 U17864 ( .A0(n15748), .A1(n15836), .B0(n15837), .C0(n15838), .Y(
        n15835) );
  AOI22X1 U17865 ( .A0(n3095), .A1(n15840), .B0(n15841), .B1(n3092), .Y(n15834) );
  OAI21XL U17866 ( .A0(n3107), .A1(n463), .B0(n1514), .Y(n15836) );
  AOI211X1 U17867 ( .A0(n17323), .A1(n17411), .B0(n17412), .C0(n17413), .Y(
        n17410) );
  AOI22X1 U17868 ( .A0(n2794), .A1(n17415), .B0(n17416), .B1(n2791), .Y(n17409) );
  OAI21XL U17869 ( .A0(n2806), .A1(n464), .B0(n1503), .Y(n17411) );
  OAI211XL U17870 ( .A0(n1803), .A1(n11779), .B0(n11734), .C0(n11864), .Y(
        n11880) );
  OAI211XL U17871 ( .A0(n1824), .A1(top_core_KE_sb1_n207), .B0(
        top_core_KE_sb1_n161), .C0(top_core_KE_sb1_n293), .Y(
        top_core_KE_sb1_n309) );
  OAI211XL U17872 ( .A0(n1761), .A1(n12410), .B0(n12365), .C0(n12495), .Y(
        n12511) );
  OAI211XL U17873 ( .A0(n1782), .A1(n12095), .B0(n12050), .C0(n12180), .Y(
        n12196) );
  OAI211XL U17874 ( .A0(n11929), .A1(n185), .B0(n11680), .C0(n11670), .Y(
        n11928) );
  OAI211XL U17875 ( .A0(top_core_KE_sb1_n358), .A1(n186), .B0(
        top_core_KE_sb1_n105), .C0(top_core_KE_sb1_n95), .Y(
        top_core_KE_sb1_n357) );
  OAI211XL U17876 ( .A0(n12560), .A1(n46), .B0(n12311), .C0(n12301), .Y(n12559) );
  OAI211XL U17877 ( .A0(n13505), .A1(n187), .B0(n13257), .C0(n13247), .Y(
        n13504) );
  OAI211XL U17878 ( .A0(n12245), .A1(n188), .B0(n11996), .C0(n11986), .Y(
        n12244) );
  OAI211XL U17879 ( .A0(n12875), .A1(n189), .B0(n12627), .C0(n12617), .Y(
        n12874) );
  OAI211XL U17880 ( .A0(n13820), .A1(n190), .B0(n13572), .C0(n13562), .Y(
        n13819) );
  OAI211XL U17881 ( .A0(n13190), .A1(n191), .B0(n12942), .C0(n12932), .Y(
        n13189) );
  OAI211XL U17882 ( .A0(n11651), .A1(n80), .B0(n11689), .C0(n11877), .Y(n11872) );
  NOR3X1 U17883 ( .A(n1204), .B(n613), .C(n11849), .Y(n11878) );
  OAI211XL U17884 ( .A0(top_core_KE_sb1_n76), .A1(n81), .B0(
        top_core_KE_sb1_n114), .C0(top_core_KE_sb1_n306), .Y(
        top_core_KE_sb1_n301) );
  NOR3X1 U17885 ( .A(n1195), .B(n614), .C(top_core_KE_sb1_n278), .Y(
        top_core_KE_sb1_n307) );
  OAI211XL U17886 ( .A0(n12283), .A1(n82), .B0(n12320), .C0(n12508), .Y(n12503) );
  NOR3X1 U17887 ( .A(n1164), .B(n601), .C(n12480), .Y(n12509) );
  NOR3X1 U17888 ( .A(n1150), .B(n1174), .C(n13425), .Y(n13454) );
  OAI211XL U17889 ( .A0(n11967), .A1(n83), .B0(n12005), .C0(n12193), .Y(n12188) );
  NOR3X1 U17890 ( .A(n1155), .B(n615), .C(n12165), .Y(n12194) );
  NOR3X1 U17891 ( .A(n1190), .B(n1214), .C(n12795), .Y(n12824) );
  NOR3X1 U17892 ( .A(n1159), .B(n1179), .C(n13740), .Y(n13769) );
  NOR3X1 U17893 ( .A(n1199), .B(n1220), .C(n13110), .Y(n13139) );
  NAND2X1 U17894 ( .A(n1635), .B(n1146), .Y(n13592) );
  NAND2X1 U17895 ( .A(n1795), .B(n1187), .Y(n11700) );
  NAND2X1 U17896 ( .A(n1816), .B(n1224), .Y(top_core_KE_sb1_n125) );
  NAND2X1 U17897 ( .A(n1670), .B(n1185), .Y(n13277) );
  NAND2X1 U17898 ( .A(n1774), .B(n1184), .Y(n12016) );
  NAND2X1 U17899 ( .A(n1728), .B(n1225), .Y(n12647) );
  NAND2X1 U17900 ( .A(n1699), .B(n1186), .Y(n12962) );
  NAND2X1 U17901 ( .A(n1752), .B(n1147), .Y(n12331) );
  NAND2X1 U17902 ( .A(n1506), .B(n3447), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n276) );
  NAND2X1 U17903 ( .A(n1504), .B(n2846), .Y(n10090) );
  NAND2X1 U17904 ( .A(n1528), .B(n2604), .Y(n11258) );
  NAND2X1 U17905 ( .A(n1518), .B(n3206), .Y(n8338) );
  NAND2X1 U17906 ( .A(n1530), .B(n2665), .Y(n10966) );
  NAND2X1 U17907 ( .A(n1511), .B(n3026), .Y(n9214) );
  NAND2X1 U17908 ( .A(n1524), .B(n3386), .Y(n7462) );
  NAND2X1 U17909 ( .A(n1502), .B(n2786), .Y(n10382) );
  NAND2X1 U17910 ( .A(n1509), .B(n2968), .Y(n9506) );
  NAND2X1 U17911 ( .A(n1515), .B(n3145), .Y(n8630) );
  NAND2X1 U17912 ( .A(n1522), .B(n3328), .Y(n7754) );
  NAND2X1 U17913 ( .A(n1525), .B(n2543), .Y(n11550) );
  NAND2X1 U17914 ( .A(n1532), .B(n2725), .Y(n10674) );
  NAND2X1 U17915 ( .A(n1507), .B(n2907), .Y(n9798) );
  NAND2X1 U17916 ( .A(n1513), .B(n3087), .Y(n8922) );
  NAND2X1 U17917 ( .A(n1520), .B(n3267), .Y(n8046) );
  NAND2X1 U17918 ( .A(n1506), .B(n3450), .Y(
        top_core_EC_ss_gen_tbox_0__sboxs_r_n278) );
  NAND2X1 U17919 ( .A(n1504), .B(n2849), .Y(n10092) );
  NAND2X1 U17920 ( .A(n1528), .B(n2607), .Y(n11260) );
  NAND2X1 U17921 ( .A(n1518), .B(n3209), .Y(n8340) );
  NAND2X1 U17922 ( .A(n1530), .B(n2668), .Y(n10968) );
  NAND2X1 U17923 ( .A(n1511), .B(n3029), .Y(n9216) );
  NAND2X1 U17924 ( .A(n1524), .B(n3389), .Y(n7464) );
  NAND2X1 U17925 ( .A(n1502), .B(n2789), .Y(n10384) );
  NAND2X1 U17926 ( .A(n1509), .B(n2971), .Y(n9508) );
  NAND2X1 U17927 ( .A(n1515), .B(n3148), .Y(n8632) );
  NAND2X1 U17928 ( .A(n1522), .B(n3331), .Y(n7756) );
  NAND2X1 U17929 ( .A(n1525), .B(n2546), .Y(n11552) );
  NAND2X1 U17930 ( .A(n1532), .B(n2728), .Y(n10676) );
  NAND2X1 U17931 ( .A(n1507), .B(n2910), .Y(n9800) );
  NAND2X1 U17932 ( .A(n1513), .B(n3090), .Y(n8924) );
  NAND2X1 U17933 ( .A(n1520), .B(n3270), .Y(n8048) );
  NOR4BX1 U17934 ( .AN(n11795), .B(n11702), .C(n11796), .D(n6917), .Y(n11794)
         );
  AOI222X1 U17935 ( .A0(n1810), .A1(n6904), .B0(n665), .B1(n11797), .C0(n753), 
        .C1(n689), .Y(n11795) );
  AOI2BB1X1 U17936 ( .A0N(n761), .A1N(n11704), .B0(n613), .Y(n11796) );
  NOR4BX1 U17937 ( .AN(top_core_KE_sb1_n223), .B(top_core_KE_sb1_n127), .C(
        top_core_KE_sb1_n224), .D(n6871), .Y(top_core_KE_sb1_n222) );
  AOI222X1 U17938 ( .A0(n1831), .A1(n6858), .B0(n666), .B1(
        top_core_KE_sb1_n225), .C0(n754), .C1(n690), .Y(top_core_KE_sb1_n223)
         );
  AOI2BB1X1 U17939 ( .A0N(n762), .A1N(top_core_KE_sb1_n129), .B0(n614), .Y(
        top_core_KE_sb1_n224) );
  NOR4BX1 U17940 ( .AN(n12426), .B(n12333), .C(n12427), .D(n6624), .Y(n12425)
         );
  AOI222X1 U17941 ( .A0(n1768), .A1(n6611), .B0(n667), .B1(n12428), .C0(n752), 
        .C1(n691), .Y(n12426) );
  AOI2BB1X1 U17942 ( .A0N(n760), .A1N(n12335), .B0(n601), .Y(n12427) );
  NOR4BX1 U17943 ( .AN(n13371), .B(n13279), .C(n13372), .D(n6552), .Y(n13370)
         );
  AOI222X1 U17944 ( .A0(n1688), .A1(n6539), .B0(n670), .B1(n13373), .C0(n748), 
        .C1(n692), .Y(n13371) );
  AOI2BB1X1 U17945 ( .A0N(n756), .A1N(n13281), .B0(n1174), .Y(n13372) );
  NOR4BX1 U17946 ( .AN(n12111), .B(n12018), .C(n12112), .D(n6577), .Y(n12110)
         );
  AOI222X1 U17947 ( .A0(n1789), .A1(n6564), .B0(n668), .B1(n12113), .C0(n755), 
        .C1(n693), .Y(n12111) );
  AOI2BB1X1 U17948 ( .A0N(n763), .A1N(n12020), .B0(n615), .Y(n12112) );
  NOR4BX1 U17949 ( .AN(n12741), .B(n12649), .C(n12742), .D(n6847), .Y(n12740)
         );
  AOI222X1 U17950 ( .A0(n1746), .A1(n6834), .B0(n671), .B1(n12743), .C0(n749), 
        .C1(n694), .Y(n12741) );
  AOI2BB1X1 U17951 ( .A0N(n757), .A1N(n12651), .B0(n1214), .Y(n12742) );
  NOR4BX1 U17952 ( .AN(n13686), .B(n13594), .C(n13687), .D(n6600), .Y(n13685)
         );
  AOI222X1 U17953 ( .A0(n1659), .A1(n6587), .B0(n669), .B1(n13688), .C0(n751), 
        .C1(n695), .Y(n13686) );
  AOI2BB1X1 U17954 ( .A0N(n759), .A1N(n13596), .B0(n1179), .Y(n13687) );
  NOR4BX1 U17955 ( .AN(n13056), .B(n12964), .C(n13057), .D(n6893), .Y(n13055)
         );
  AOI222X1 U17956 ( .A0(n1717), .A1(n6880), .B0(n672), .B1(n13058), .C0(n750), 
        .C1(n696), .Y(n13056) );
  AOI2BB1X1 U17957 ( .A0N(n758), .A1N(n12966), .B0(n1220), .Y(n13057) );
  NOR2X1 U17958 ( .A(n12340), .B(n691), .Y(n12366) );
  NOR2X1 U17959 ( .A(n11709), .B(n689), .Y(n11735) );
  NOR2X1 U17960 ( .A(top_core_KE_sb1_n134), .B(n690), .Y(top_core_KE_sb1_n162)
         );
  NOR2X1 U17961 ( .A(n12025), .B(n693), .Y(n12051) );
  NAND3XL U17962 ( .A(n12278), .B(n1171), .C(n12400), .Y(n12515) );
  AOI31X1 U17963 ( .A0(n13301), .A1(n13302), .A2(n6543), .B0(n13217), .Y(
        n13300) );
  INVX1 U17964 ( .A(n13303), .Y(n6543) );
  OAI21XL U17965 ( .A0(n187), .A1(n13294), .B0(n13304), .Y(n13303) );
  AOI31X1 U17966 ( .A0(n12671), .A1(n12672), .A2(n6838), .B0(n12587), .Y(
        n12670) );
  INVX1 U17967 ( .A(n12673), .Y(n6838) );
  OAI21XL U17968 ( .A0(n189), .A1(n12664), .B0(n12674), .Y(n12673) );
  AOI31X1 U17969 ( .A0(n12986), .A1(n12987), .A2(n6884), .B0(n12902), .Y(
        n12985) );
  INVX1 U17970 ( .A(n12988), .Y(n6884) );
  OAI21XL U17971 ( .A0(n191), .A1(n12979), .B0(n12989), .Y(n12988) );
  AOI31X1 U17972 ( .A0(n12355), .A1(n12356), .A2(n6615), .B0(n12272), .Y(
        n12354) );
  INVX1 U17973 ( .A(n12357), .Y(n6615) );
  OAI21XL U17974 ( .A0(n46), .A1(n12348), .B0(n12358), .Y(n12357) );
  AOI31X1 U17975 ( .A0(n13616), .A1(n13617), .A2(n6591), .B0(n13532), .Y(
        n13615) );
  INVX1 U17976 ( .A(n13618), .Y(n6591) );
  OAI21XL U17977 ( .A0(n190), .A1(n13609), .B0(n13619), .Y(n13618) );
  AOI31X1 U17978 ( .A0(n11724), .A1(n11725), .A2(n6908), .B0(n11640), .Y(
        n11723) );
  INVX1 U17979 ( .A(n11726), .Y(n6908) );
  OAI21XL U17980 ( .A0(n185), .A1(n11717), .B0(n11727), .Y(n11726) );
  AOI31X1 U17981 ( .A0(top_core_KE_sb1_n151), .A1(top_core_KE_sb1_n152), .A2(
        n6862), .B0(top_core_KE_sb1_n65), .Y(top_core_KE_sb1_n150) );
  INVX1 U17982 ( .A(top_core_KE_sb1_n153), .Y(n6862) );
  OAI21XL U17983 ( .A0(n186), .A1(top_core_KE_sb1_n144), .B0(
        top_core_KE_sb1_n154), .Y(top_core_KE_sb1_n153) );
  AOI31X1 U17984 ( .A0(n12040), .A1(n12041), .A2(n6568), .B0(n11956), .Y(
        n12039) );
  INVX1 U17985 ( .A(n12042), .Y(n6568) );
  OAI21XL U17986 ( .A0(n188), .A1(n12033), .B0(n12043), .Y(n12042) );
  AOI31X1 U17987 ( .A0(n13733), .A1(n13734), .A2(n13735), .B0(n13592), .Y(
        n13732) );
  AOI222X1 U17988 ( .A0(n13628), .A1(n751), .B0(n1157), .B1(n1663), .C0(n679), 
        .C1(n1161), .Y(n13735) );
  AOI22X1 U17989 ( .A0(n6592), .A1(n1658), .B0(n6587), .B1(n1179), .Y(n13733)
         );
  AOI31X1 U17990 ( .A0(n11842), .A1(n11843), .A2(n11844), .B0(n11700), .Y(
        n11841) );
  AOI222X1 U17991 ( .A0(n11736), .A1(n753), .B0(n1202), .B1(n1814), .C0(n673), 
        .C1(n1205), .Y(n11844) );
  AOI22X1 U17992 ( .A0(n6909), .A1(n1809), .B0(n6904), .B1(n605), .Y(n11842)
         );
  AOI31X1 U17993 ( .A0(top_core_KE_sb1_n271), .A1(top_core_KE_sb1_n272), .A2(
        top_core_KE_sb1_n273), .B0(top_core_KE_sb1_n125), .Y(
        top_core_KE_sb1_n270) );
  AOI222X1 U17994 ( .A0(top_core_KE_sb1_n163), .A1(n754), .B0(n1193), .B1(
        n1835), .C0(n674), .C1(n1196), .Y(top_core_KE_sb1_n273) );
  AOI22X1 U17995 ( .A0(n6863), .A1(n1830), .B0(n6858), .B1(n606), .Y(
        top_core_KE_sb1_n271) );
  AOI31X1 U17996 ( .A0(n12473), .A1(n12474), .A2(n12475), .B0(n12331), .Y(
        n12472) );
  AOI222X1 U17997 ( .A0(n12367), .A1(n752), .B0(n1162), .B1(n1773), .C0(n675), 
        .C1(n1165), .Y(n12475) );
  AOI22X1 U17998 ( .A0(n6616), .A1(n1767), .B0(n6611), .B1(n607), .Y(n12473)
         );
  AOI31X1 U17999 ( .A0(n12158), .A1(n12159), .A2(n12160), .B0(n12016), .Y(
        n12157) );
  AOI222X1 U18000 ( .A0(n12052), .A1(n755), .B0(n1153), .B1(n1793), .C0(n676), 
        .C1(n1156), .Y(n12160) );
  AOI22X1 U18001 ( .A0(n6569), .A1(n1788), .B0(n6564), .B1(n608), .Y(n12158)
         );
  NOR2XL U18002 ( .A(n7008), .B(top_core_KE_n1865), .Y(top_core_KE_n2703) );
  INVX1 U18003 ( .A(top_core_KE_n2183), .Y(n6483) );
  NOR2XL U18004 ( .A(n80), .B(n1797), .Y(n11656) );
  NOR2XL U18005 ( .A(n81), .B(n1818), .Y(top_core_KE_sb1_n81) );
  NOR2XL U18006 ( .A(n82), .B(n1754), .Y(n12288) );
  NOR2XL U18007 ( .A(n83), .B(n1776), .Y(n11972) );
  NOR2XL U18008 ( .A(n76), .B(top_core_KE_prev_key1_reg_93_), .Y(n13548) );
  NOR2X1 U18009 ( .A(n697), .B(n627), .Y(n12560) );
  XNOR2X1 U18010 ( .A(n1171), .B(n1767), .Y(n697) );
  NAND2X1 U18011 ( .A(n6306), .B(top_core_EC_n943), .Y(top_core_EC_n870) );
  NAND2X1 U18012 ( .A(top_core_KE_n1864), .B(n2142), .Y(top_core_KE_n2695) );
  NAND2X1 U18013 ( .A(n13373), .B(n1688), .Y(n13444) );
  NAND2X1 U18014 ( .A(n11797), .B(n1809), .Y(n11868) );
  NAND2X1 U18015 ( .A(top_core_KE_sb1_n225), .B(n1830), .Y(
        top_core_KE_sb1_n297) );
  NAND2X1 U18016 ( .A(n12428), .B(n1767), .Y(n12499) );
  NAND2X1 U18017 ( .A(n12113), .B(n1788), .Y(n12184) );
  NAND2X1 U18018 ( .A(n12743), .B(n1746), .Y(n12814) );
  NAND2X1 U18019 ( .A(n13688), .B(n1658), .Y(n13759) );
  NAND2X1 U18020 ( .A(n13058), .B(n1717), .Y(n13129) );
  OAI22XL U18021 ( .A0(n1505), .A1(n433), .B0(n17093), .B1(n17075), .Y(n17101)
         );
  OAI22XL U18022 ( .A0(n1517), .A1(n434), .B0(n13943), .B1(n13925), .Y(n13951)
         );
  OAI22XL U18023 ( .A0(n1529), .A1(n435), .B0(n18353), .B1(n18335), .Y(n18361)
         );
  OAI22XL U18024 ( .A0(n1519), .A1(n436), .B0(n15203), .B1(n15185), .Y(n15211)
         );
  OAI22XL U18025 ( .A0(n1516), .A1(n437), .B0(n15518), .B1(n15500), .Y(n15526)
         );
  OAI22XL U18026 ( .A0(n1526), .A1(n439), .B0(n18668), .B1(n18650), .Y(n18676)
         );
  OAI22XL U18027 ( .A0(n1508), .A1(n438), .B0(n16778), .B1(n16760), .Y(n16786)
         );
  OAI22XL U18028 ( .A0(n1521), .A1(n440), .B0(n14888), .B1(n14870), .Y(n14896)
         );
  OAI22XL U18029 ( .A0(n1510), .A1(n441), .B0(n16463), .B1(n16445), .Y(n16471)
         );
  OAI22XL U18030 ( .A0(n1531), .A1(n442), .B0(n18038), .B1(n18020), .Y(n18046)
         );
  OAI22XL U18031 ( .A0(n1523), .A1(n443), .B0(n14573), .B1(n14555), .Y(n14581)
         );
  OAI22XL U18032 ( .A0(n1512), .A1(n444), .B0(n16148), .B1(n16130), .Y(n16156)
         );
  OAI22XL U18033 ( .A0(n1501), .A1(n445), .B0(n17723), .B1(n17705), .Y(n17731)
         );
  OAI22XL U18034 ( .A0(n1527), .A1(n446), .B0(n14258), .B1(n14240), .Y(n14266)
         );
  OAI22XL U18035 ( .A0(n1514), .A1(n447), .B0(n15833), .B1(n15815), .Y(n15841)
         );
  OAI22XL U18036 ( .A0(n1503), .A1(n448), .B0(n17408), .B1(n17390), .Y(n17416)
         );
  CLKINVX3 U18037 ( .A(n11716), .Y(n6914) );
  CLKINVX3 U18038 ( .A(top_core_KE_sb1_n143), .Y(n6868) );
  CLKINVX3 U18039 ( .A(n12347), .Y(n6621) );
  CLKINVX3 U18040 ( .A(n12032), .Y(n6574) );
  INVX1 U18041 ( .A(top_core_KE_n896), .Y(n7021) );
  NAND2X1 U18042 ( .A(n13240), .B(n1172), .Y(n13330) );
  NAND2X1 U18043 ( .A(n12610), .B(n1212), .Y(n12700) );
  NAND2X1 U18044 ( .A(n12925), .B(n1218), .Y(n13015) );
  NAND2X1 U18045 ( .A(n13555), .B(n1180), .Y(n13645) );
  NAND2X1 U18046 ( .A(n12294), .B(n1183), .Y(n12384) );
  NAND2X1 U18047 ( .A(n11663), .B(n1221), .Y(n11753) );
  NAND2X1 U18048 ( .A(top_core_KE_sb1_n88), .B(n1215), .Y(top_core_KE_sb1_n181) );
  NAND2X1 U18049 ( .A(n11979), .B(n1175), .Y(n12069) );
  NAND2X1 U18050 ( .A(n13593), .B(n1635), .Y(n13765) );
  NAND2X1 U18051 ( .A(n11701), .B(n1795), .Y(n11874) );
  NAND2X1 U18052 ( .A(top_core_KE_sb1_n126), .B(n1816), .Y(
        top_core_KE_sb1_n303) );
  NAND2X1 U18053 ( .A(n12017), .B(n1774), .Y(n12190) );
  NAND2X1 U18054 ( .A(n12332), .B(n1752), .Y(n12505) );
  AOI22X1 U18055 ( .A0(n6745), .A1(n11846), .B0(n6746), .B1(n11847), .Y(n11845) );
  NAND4XL U18056 ( .A(n11807), .B(n11718), .C(n11724), .D(n11848), .Y(n11847)
         );
  NAND4BXL U18057 ( .AN(n11850), .B(n11671), .C(n11787), .D(n11851), .Y(n11846) );
  AOI22X1 U18058 ( .A0(n6807), .A1(top_core_KE_sb1_n275), .B0(n6801), .B1(
        top_core_KE_sb1_n276), .Y(top_core_KE_sb1_n274) );
  NAND4XL U18059 ( .A(top_core_KE_sb1_n235), .B(top_core_KE_sb1_n145), .C(
        top_core_KE_sb1_n151), .D(top_core_KE_sb1_n277), .Y(
        top_core_KE_sb1_n276) );
  NAND4BXL U18060 ( .AN(top_core_KE_sb1_n279), .B(top_core_KE_sb1_n96), .C(
        top_core_KE_sb1_n215), .D(top_core_KE_sb1_n280), .Y(
        top_core_KE_sb1_n275) );
  AOI22X1 U18061 ( .A0(n6442), .A1(n12477), .B0(n6443), .B1(n12478), .Y(n12476) );
  NAND4XL U18062 ( .A(n12438), .B(n12349), .C(n12355), .D(n12479), .Y(n12478)
         );
  NAND4BXL U18063 ( .AN(n12481), .B(n12302), .C(n12418), .D(n12482), .Y(n12477) );
  AOI22X1 U18064 ( .A0(n6510), .A1(n12162), .B0(n6504), .B1(n12163), .Y(n12161) );
  NAND4XL U18065 ( .A(n12123), .B(n12034), .C(n12040), .D(n12164), .Y(n12163)
         );
  NAND4BXL U18066 ( .AN(n12166), .B(n11987), .C(n12103), .D(n12167), .Y(n12162) );
  AOI22X1 U18067 ( .A0(n6778), .A1(n12792), .B0(n6772), .B1(n12793), .Y(n12791) );
  NAND4XL U18068 ( .A(n12753), .B(n12665), .C(n12671), .D(n12794), .Y(n12793)
         );
  NAND4BXL U18069 ( .AN(n12796), .B(n12618), .C(n12733), .D(n12797), .Y(n12792) );
  AOI22X1 U18070 ( .A0(n6433), .A1(n13737), .B0(n6434), .B1(n13738), .Y(n13736) );
  NAND4XL U18071 ( .A(n13698), .B(n13610), .C(n13616), .D(n13739), .Y(n13738)
         );
  NAND4BXL U18072 ( .AN(n13741), .B(n13563), .C(n13678), .D(n13742), .Y(n13737) );
  AOI22X1 U18073 ( .A0(n6714), .A1(n13107), .B0(n6715), .B1(n13108), .Y(n13106) );
  NAND4XL U18074 ( .A(n13068), .B(n12980), .C(n12986), .D(n13109), .Y(n13108)
         );
  NAND4BXL U18075 ( .AN(n13111), .B(n12933), .C(n13048), .D(n13112), .Y(n13107) );
  NAND2X1 U18076 ( .A(n13278), .B(n1671), .Y(n13450) );
  NAND2X1 U18077 ( .A(n12648), .B(n1726), .Y(n12820) );
  NAND2X1 U18078 ( .A(n12963), .B(n1697), .Y(n13135) );
  AOI22X1 U18079 ( .A0(n13373), .A1(n580), .B0(n6636), .B1(n1673), .Y(n13446)
         );
  NAND2X1 U18080 ( .A(top_core_KE_n2704), .B(n743), .Y(top_core_KE_n2701) );
  INVX1 U18081 ( .A(n13532), .Y(n6434) );
  INVX1 U18082 ( .A(n11640), .Y(n6746) );
  INVX1 U18083 ( .A(top_core_KE_sb1_n65), .Y(n6801) );
  INVX1 U18084 ( .A(n12272), .Y(n6443) );
  INVX1 U18085 ( .A(n11956), .Y(n6504) );
  INVX1 U18086 ( .A(n13217), .Y(n6469) );
  INVX1 U18087 ( .A(n12587), .Y(n6772) );
  INVX1 U18088 ( .A(n12902), .Y(n6715) );
  NAND2XL U18089 ( .A(n82), .B(n12437), .Y(n12273) );
  NAND2XL U18090 ( .A(n80), .B(n11806), .Y(n11641) );
  NAND2XL U18091 ( .A(n81), .B(top_core_KE_sb1_n234), .Y(top_core_KE_sb1_n66)
         );
  NAND2XL U18092 ( .A(n83), .B(n12122), .Y(n11957) );
  NAND4X1 U18093 ( .A(n6922), .B(n11716), .C(n11884), .D(n11885), .Y(n11881)
         );
  AOI221X1 U18094 ( .A0(n6920), .A1(n1222), .B0(n11819), .B1(n1221), .C0(
        n11886), .Y(n11885) );
  AOI21XL U18095 ( .A0(n50), .A1(n11733), .B0(n1806), .Y(n11886) );
  NAND4X1 U18096 ( .A(n6876), .B(top_core_KE_sb1_n143), .C(
        top_core_KE_sb1_n313), .D(top_core_KE_sb1_n314), .Y(
        top_core_KE_sb1_n310) );
  AOI221X1 U18097 ( .A0(n6874), .A1(n1216), .B0(top_core_KE_sb1_n247), .B1(
        n1215), .C0(top_core_KE_sb1_n315), .Y(top_core_KE_sb1_n314) );
  AOI21XL U18098 ( .A0(n51), .A1(top_core_KE_sb1_n160), .B0(n1827), .Y(
        top_core_KE_sb1_n315) );
  NAND4X1 U18099 ( .A(n6629), .B(n12347), .C(n12515), .D(n12516), .Y(n12512)
         );
  AOI221X1 U18100 ( .A0(n6627), .A1(n1181), .B0(n12450), .B1(n1183), .C0(
        n12517), .Y(n12516) );
  AOI21XL U18101 ( .A0(n89), .A1(n12364), .B0(n1764), .Y(n12517) );
  NAND4X1 U18102 ( .A(n6558), .B(n13293), .C(n13460), .D(n13461), .Y(n13457)
         );
  AOI221X1 U18103 ( .A0(n6556), .A1(n1173), .B0(n13395), .B1(n1172), .C0(
        n13462), .Y(n13461) );
  AOI21XL U18104 ( .A0(n52), .A1(n13310), .B0(n1682), .Y(n13462) );
  NAND4X1 U18105 ( .A(n6582), .B(n12032), .C(n12200), .D(n12201), .Y(n12197)
         );
  AOI221X1 U18106 ( .A0(n6580), .A1(n1176), .B0(n12135), .B1(n1175), .C0(
        n12202), .Y(n12201) );
  AOI21XL U18107 ( .A0(n53), .A1(n12049), .B0(n1785), .Y(n12202) );
  NAND4X1 U18108 ( .A(n6853), .B(n12663), .C(n12830), .D(n12831), .Y(n12827)
         );
  AOI221X1 U18109 ( .A0(n6851), .A1(n1213), .B0(n12765), .B1(n1212), .C0(
        n12832), .Y(n12831) );
  AOI21XL U18110 ( .A0(n54), .A1(n12680), .B0(n1740), .Y(n12832) );
  NAND4X1 U18111 ( .A(n6606), .B(n13608), .C(n13775), .D(n13776), .Y(n13772)
         );
  AOI221X1 U18112 ( .A0(n6604), .A1(n1178), .B0(n13710), .B1(n1180), .C0(
        n13777), .Y(n13776) );
  AOI21XL U18113 ( .A0(n55), .A1(n13625), .B0(n1655), .Y(n13777) );
  NAND4X1 U18114 ( .A(n6899), .B(n12978), .C(n13145), .D(n13146), .Y(n13142)
         );
  AOI221X1 U18115 ( .A0(n6897), .A1(n1219), .B0(n13080), .B1(n1218), .C0(
        n13147), .Y(n13146) );
  AOI21XL U18116 ( .A0(n56), .A1(n12995), .B0(n1711), .Y(n13147) );
  XNOR2X1 U18117 ( .A(top_core_KE_new_sboxw_15_), .B(top_core_KE_n2030), .Y(
        top_core_KE_n1485) );
  XNOR2X1 U18118 ( .A(top_core_KE_new_sboxw_13_), .B(top_core_KE_n2036), .Y(
        top_core_KE_n1501) );
  XNOR2X1 U18119 ( .A(top_core_KE_new_sboxw_10_), .B(top_core_KE_n2045), .Y(
        top_core_KE_n1525) );
  XNOR2X1 U18120 ( .A(top_core_KE_new_sboxw_7_), .B(top_core_KE_n2054), .Y(
        top_core_KE_n1549) );
  XNOR2X1 U18121 ( .A(top_core_KE_new_sboxw_5_), .B(top_core_KE_n2060), .Y(
        top_core_KE_n1565) );
  XNOR2X1 U18122 ( .A(top_core_KE_new_sboxw_2_), .B(top_core_KE_n2069), .Y(
        top_core_KE_n1589) );
  XNOR2X1 U18123 ( .A(top_core_KE_new_sboxw_29_), .B(top_core_KE_n1983), .Y(
        top_core_KE_n1373) );
  XNOR2X1 U18124 ( .A(top_core_KE_new_sboxw_26_), .B(top_core_KE_n1995), .Y(
        top_core_KE_n1397) );
  XNOR2X1 U18125 ( .A(top_core_KE_new_sboxw_31_), .B(top_core_KE_n1975), .Y(
        top_core_KE_n1358) );
  INVX1 U18126 ( .A(n13307), .Y(n6475) );
  INVX1 U18127 ( .A(n12992), .Y(n6714) );
  INVX1 U18128 ( .A(n12677), .Y(n6778) );
  INVX1 U18129 ( .A(n11730), .Y(n6745) );
  INVX1 U18130 ( .A(top_core_KE_sb1_n157), .Y(n6807) );
  INVX1 U18131 ( .A(n12361), .Y(n6442) );
  INVX1 U18132 ( .A(n12046), .Y(n6510) );
  INVX1 U18133 ( .A(n13622), .Y(n6433) );
  XOR2X1 U18134 ( .A(n6483), .B(top_core_KE_n1975), .Y(top_core_KE_n1359) );
  AOI21X1 U18135 ( .A0(n11742), .A1(n11650), .B0(n11679), .Y(n11740) );
  AOI21X1 U18136 ( .A0(top_core_KE_sb1_n169), .A1(top_core_KE_sb1_n75), .B0(
        top_core_KE_sb1_n104), .Y(top_core_KE_sb1_n167) );
  AOI21X1 U18137 ( .A0(n12373), .A1(n12282), .B0(n12310), .Y(n12371) );
  AOI21X1 U18138 ( .A0(n13319), .A1(n13227), .B0(n13256), .Y(n13317) );
  AOI21X1 U18139 ( .A0(n12058), .A1(n11966), .B0(n11995), .Y(n12056) );
  AOI21X1 U18140 ( .A0(n12689), .A1(n12597), .B0(n12626), .Y(n12687) );
  AOI21X1 U18141 ( .A0(n13004), .A1(n12912), .B0(n12941), .Y(n13002) );
  AOI21X1 U18142 ( .A0(n13634), .A1(n13542), .B0(n13571), .Y(n13632) );
  XNOR2X1 U18143 ( .A(top_core_KE_new_sboxw_23_), .B(top_core_KE_n2006), .Y(
        top_core_KE_n1421) );
  XNOR2X1 U18144 ( .A(top_core_KE_new_sboxw_21_), .B(top_core_KE_n2012), .Y(
        top_core_KE_n1437) );
  XNOR2X1 U18145 ( .A(top_core_KE_new_sboxw_18_), .B(top_core_KE_n2021), .Y(
        top_core_KE_n1461) );
  OAI21XL U18146 ( .A0(n1802), .A1(n80), .B0(n11669), .Y(n11743) );
  OAI21XL U18147 ( .A0(n1823), .A1(n81), .B0(top_core_KE_sb1_n94), .Y(
        top_core_KE_sb1_n170) );
  OAI21XL U18148 ( .A0(n1760), .A1(n82), .B0(n12300), .Y(n12374) );
  OAI21XL U18149 ( .A0(n1781), .A1(n83), .B0(n11985), .Y(n12059) );
  AOI22X1 U18150 ( .A0(n629), .A1(n13289), .B0(n6462), .B1(n13362), .Y(n13361)
         );
  NAND4X1 U18151 ( .A(n13363), .B(n6558), .C(n13364), .D(n13365), .Y(n13362)
         );
  NAND3XL U18152 ( .A(n13346), .B(n13282), .C(n1674), .Y(n13364) );
  AOI22X1 U18153 ( .A0(n630), .A1(n12659), .B0(n6763), .B1(n12732), .Y(n12731)
         );
  NAND4X1 U18154 ( .A(n12733), .B(n6853), .C(n12734), .D(n12735), .Y(n12732)
         );
  NAND3XL U18155 ( .A(n12716), .B(n12652), .C(n1732), .Y(n12734) );
  AOI22X1 U18156 ( .A0(n631), .A1(n13604), .B0(n6419), .B1(n13677), .Y(n13676)
         );
  NAND4X1 U18157 ( .A(n13678), .B(n6606), .C(n13679), .D(n13680), .Y(n13677)
         );
  NAND3XL U18158 ( .A(n13661), .B(n13597), .C(n1645), .Y(n13679) );
  AOI22X1 U18159 ( .A0(n632), .A1(n12974), .B0(n6706), .B1(n13047), .Y(n13046)
         );
  NAND4X1 U18160 ( .A(n13048), .B(n6899), .C(n13049), .D(n13050), .Y(n13047)
         );
  NAND3XL U18161 ( .A(n13031), .B(n12967), .C(n1703), .Y(n13049) );
  XNOR2X1 U18162 ( .A(top_core_KE_new_sboxw_14_), .B(top_core_KE_n2033), .Y(
        top_core_KE_n1493) );
  XNOR2X1 U18163 ( .A(top_core_KE_new_sboxw_8_), .B(top_core_KE_n2051), .Y(
        top_core_KE_n1541) );
  XNOR2X1 U18164 ( .A(top_core_KE_new_sboxw_6_), .B(top_core_KE_n2057), .Y(
        top_core_KE_n1557) );
  XNOR2X1 U18165 ( .A(top_core_KE_new_sboxw_0_), .B(top_core_KE_n2075), .Y(
        top_core_KE_n1605) );
  XNOR2X1 U18166 ( .A(top_core_KE_new_sboxw_30_), .B(top_core_KE_n1979), .Y(
        top_core_KE_n1365) );
  XNOR2X1 U18167 ( .A(top_core_KE_new_sboxw_24_), .B(top_core_KE_n2003), .Y(
        top_core_KE_n1413) );
  XNOR2X1 U18168 ( .A(top_core_KE_new_sboxw_9_), .B(top_core_KE_n2048), .Y(
        top_core_KE_n1533) );
  XNOR2X1 U18169 ( .A(top_core_KE_new_sboxw_1_), .B(top_core_KE_n2072), .Y(
        top_core_KE_n1597) );
  XNOR2X1 U18170 ( .A(top_core_KE_new_sboxw_25_), .B(top_core_KE_n1999), .Y(
        top_core_KE_n1405) );
  XNOR2X1 U18171 ( .A(top_core_KE_new_sboxw_12_), .B(top_core_KE_n2039), .Y(
        top_core_KE_n1509) );
  XNOR2X1 U18172 ( .A(top_core_KE_new_sboxw_11_), .B(top_core_KE_n2042), .Y(
        top_core_KE_n1517) );
  XNOR2X1 U18173 ( .A(top_core_KE_new_sboxw_4_), .B(top_core_KE_n2063), .Y(
        top_core_KE_n1573) );
  XNOR2X1 U18174 ( .A(top_core_KE_new_sboxw_3_), .B(top_core_KE_n2066), .Y(
        top_core_KE_n1581) );
  XNOR2X1 U18175 ( .A(top_core_KE_new_sboxw_28_), .B(top_core_KE_n1987), .Y(
        top_core_KE_n1381) );
  XNOR2X1 U18176 ( .A(top_core_KE_new_sboxw_27_), .B(top_core_KE_n1991), .Y(
        top_core_KE_n1389) );
  AOI21XL U18177 ( .A0(n11709), .A1(n11769), .B0(n6952), .Y(n11930) );
  INVX1 U18178 ( .A(n11868), .Y(n6952) );
  AOI21XL U18179 ( .A0(top_core_KE_sb1_n134), .A1(top_core_KE_sb1_n197), .B0(
        n6937), .Y(top_core_KE_sb1_n359) );
  INVX1 U18180 ( .A(top_core_KE_sb1_n297), .Y(n6937) );
  AOI21XL U18181 ( .A0(n12340), .A1(n12400), .B0(n6662), .Y(n12561) );
  INVX1 U18182 ( .A(n12499), .Y(n6662) );
  AOI21XL U18183 ( .A0(n12025), .A1(n12085), .B0(n6646), .Y(n12246) );
  INVX1 U18184 ( .A(n12184), .Y(n6646) );
  XNOR2X1 U18185 ( .A(n6735), .B(top_core_KE_n2006), .Y(top_core_KE_n1423) );
  XNOR2X1 U18186 ( .A(n6722), .B(top_core_KE_n2012), .Y(top_core_KE_n1439) );
  XNOR2X1 U18187 ( .A(n6728), .B(top_core_KE_n2021), .Y(top_core_KE_n1463) );
  XNOR2X1 U18188 ( .A(n6785), .B(top_core_KE_n2030), .Y(top_core_KE_n1487) );
  XNOR2X1 U18189 ( .A(n6787), .B(top_core_KE_n2036), .Y(top_core_KE_n1503) );
  XNOR2X1 U18190 ( .A(n6792), .B(top_core_KE_n2045), .Y(top_core_KE_n1527) );
  XNOR2X1 U18191 ( .A(n6359), .B(top_core_KE_n2054), .Y(top_core_KE_n1551) );
  XNOR2X1 U18192 ( .A(n6361), .B(top_core_KE_n2060), .Y(top_core_KE_n1567) );
  XNOR2X1 U18193 ( .A(n6369), .B(top_core_KE_n2069), .Y(top_core_KE_n1591) );
  XNOR2X1 U18194 ( .A(top_core_KE_n2517), .B(top_core_KE_n1983), .Y(
        top_core_KE_n1375) );
  XNOR2X1 U18195 ( .A(top_core_KE_n2526), .B(top_core_KE_n1995), .Y(
        top_core_KE_n1399) );
  XNOR2X1 U18196 ( .A(top_core_KE_n2514), .B(top_core_KE_n1979), .Y(
        top_core_KE_n1367) );
  XNOR2X1 U18197 ( .A(top_core_KE_n2520), .B(top_core_KE_n1987), .Y(
        top_core_KE_n1383) );
  XNOR2X1 U18198 ( .A(top_core_KE_n2523), .B(top_core_KE_n1991), .Y(
        top_core_KE_n1391) );
  XNOR2X1 U18199 ( .A(top_core_KE_n2529), .B(top_core_KE_n1999), .Y(
        top_core_KE_n1407) );
  XNOR2X1 U18200 ( .A(top_core_KE_n2532), .B(top_core_KE_n2003), .Y(
        top_core_KE_n1415) );
  XNOR2X1 U18201 ( .A(n6721), .B(top_core_KE_n2009), .Y(top_core_KE_n1431) );
  XNOR2X1 U18202 ( .A(n6739), .B(top_core_KE_n2027), .Y(top_core_KE_n1479) );
  XNOR2X1 U18203 ( .A(n6786), .B(top_core_KE_n2033), .Y(top_core_KE_n1495) );
  XNOR2X1 U18204 ( .A(n6797), .B(top_core_KE_n2051), .Y(top_core_KE_n1543) );
  XNOR2X1 U18205 ( .A(n6347), .B(top_core_KE_n2057), .Y(top_core_KE_n1559) );
  XNOR2X1 U18206 ( .A(n6355), .B(top_core_KE_n2075), .Y(top_core_KE_n1607) );
  XNOR2X1 U18207 ( .A(n6725), .B(top_core_KE_n2015), .Y(top_core_KE_n1447) );
  XNOR2X1 U18208 ( .A(n6732), .B(top_core_KE_n2018), .Y(top_core_KE_n1455) );
  XNOR2X1 U18209 ( .A(n6736), .B(top_core_KE_n2024), .Y(top_core_KE_n1471) );
  XNOR2X1 U18210 ( .A(n6788), .B(top_core_KE_n2039), .Y(top_core_KE_n1511) );
  XNOR2X1 U18211 ( .A(n6790), .B(top_core_KE_n2042), .Y(top_core_KE_n1519) );
  XNOR2X1 U18212 ( .A(n6795), .B(top_core_KE_n2048), .Y(top_core_KE_n1535) );
  XNOR2X1 U18213 ( .A(n6351), .B(top_core_KE_n2063), .Y(top_core_KE_n1575) );
  XNOR2X1 U18214 ( .A(n6365), .B(top_core_KE_n2066), .Y(top_core_KE_n1583) );
  XNOR2X1 U18215 ( .A(n6374), .B(top_core_KE_n2072), .Y(top_core_KE_n1599) );
  OAI21XL U18216 ( .A0(n631), .A1(n1168), .B0(n1276), .Y(n13657) );
  OAI21XL U18217 ( .A0(n625), .A1(n1209), .B0(n1257), .Y(n11765) );
  OAI21XL U18218 ( .A0(n626), .A1(n1207), .B0(n1329), .Y(top_core_KE_sb1_n193)
         );
  OAI21XL U18219 ( .A0(n629), .A1(n1166), .B0(n1273), .Y(n13342) );
  OAI21XL U18220 ( .A0(n628), .A1(n1167), .B0(n1260), .Y(n12081) );
  OAI21XL U18221 ( .A0(n630), .A1(n1206), .B0(n1267), .Y(n12712) );
  OAI21XL U18222 ( .A0(n632), .A1(n1208), .B0(n1270), .Y(n13027) );
  AOI2BB2X1 U18223 ( .B0(n6826), .B1(n11798), .A0N(n50), .A1N(n11662), .Y(
        n11910) );
  AOI2BB2X1 U18224 ( .B0(n6804), .B1(top_core_KE_sb1_n226), .A0N(n51), .A1N(
        top_core_KE_sb1_n87), .Y(top_core_KE_sb1_n339) );
  AOI2BB2X1 U18225 ( .B0(n6530), .B1(n12429), .A0N(n89), .A1N(n12293), .Y(
        n12541) );
  AOI2BB2X1 U18226 ( .B0(n6507), .B1(n12114), .A0N(n53), .A1N(n11978), .Y(
        n12226) );
  AOI2BB2X1 U18227 ( .B0(n6519), .B1(n13689), .A0N(n55), .A1N(n13554), .Y(
        n13801) );
  XNOR2X1 U18228 ( .A(top_core_KE_new_sboxw_22_), .B(top_core_KE_n2009), .Y(
        top_core_KE_n1429) );
  XNOR2X1 U18229 ( .A(top_core_KE_new_sboxw_16_), .B(top_core_KE_n2027), .Y(
        top_core_KE_n1477) );
  XNOR2X1 U18230 ( .A(n6995), .B(top_core_KE_n1081), .Y(top_core_KE_n1305) );
  XNOR2X1 U18231 ( .A(n6994), .B(top_core_KE_n1025), .Y(top_core_KE_n1249) );
  XNOR2X1 U18232 ( .A(n6990), .B(top_core_KE_n969), .Y(top_core_KE_n1193) );
  XNOR2X1 U18233 ( .A(n1705), .B(top_core_KE_n1060), .Y(top_core_KE_n1284) );
  XNOR2X1 U18234 ( .A(n1734), .B(top_core_KE_n1116), .Y(top_core_KE_n1340) );
  XNOR2X1 U18235 ( .A(n1699), .B(top_core_KE_n1039), .Y(top_core_KE_n1263) );
  XNOR2X1 U18236 ( .A(n1728), .B(top_core_KE_n1095), .Y(top_core_KE_n1319) );
  XNOR2X1 U18237 ( .A(n1677), .B(top_core_KE_n1004), .Y(top_core_KE_n1228) );
  XNOR2X1 U18238 ( .A(n1670), .B(top_core_KE_n983), .Y(top_core_KE_n1207) );
  XNOR2X1 U18239 ( .A(n1225), .B(top_core_KE_n1088), .Y(top_core_KE_n1312) );
  XNOR2X1 U18240 ( .A(n1722), .B(top_core_KE_n1074), .Y(top_core_KE_n1298) );
  XNOR2X1 U18241 ( .A(n1751), .B(top_core_KE_n1130), .Y(top_core_KE_n1354) );
  XNOR2X1 U18242 ( .A(n1712), .B(top_core_KE_n1067), .Y(top_core_KE_n1291) );
  XNOR2X1 U18243 ( .A(n1741), .B(top_core_KE_n1123), .Y(top_core_KE_n1347) );
  XNOR2X1 U18244 ( .A(n1208), .B(top_core_KE_n1053), .Y(top_core_KE_n1277) );
  XNOR2X1 U18245 ( .A(n1206), .B(top_core_KE_n1109), .Y(top_core_KE_n1333) );
  XNOR2X1 U18246 ( .A(n1199), .B(top_core_KE_n1046), .Y(top_core_KE_n1270) );
  XNOR2X1 U18247 ( .A(n1190), .B(top_core_KE_n1102), .Y(top_core_KE_n1326) );
  XNOR2X1 U18248 ( .A(n1186), .B(top_core_KE_n1032), .Y(top_core_KE_n1256) );
  XNOR2X1 U18249 ( .A(n1185), .B(top_core_KE_n976), .Y(top_core_KE_n1200) );
  XNOR2X1 U18250 ( .A(n1693), .B(top_core_KE_n1018), .Y(top_core_KE_n1242) );
  XNOR2X1 U18251 ( .A(n1683), .B(top_core_KE_n1011), .Y(top_core_KE_n1235) );
  XNOR2X1 U18252 ( .A(n1166), .B(top_core_KE_n997), .Y(top_core_KE_n1221) );
  XNOR2X1 U18253 ( .A(n1150), .B(top_core_KE_n990), .Y(top_core_KE_n1214) );
  OAI21XL U18254 ( .A0(n627), .A1(n1169), .B0(n1264), .Y(n12396) );
  XNOR2X1 U18255 ( .A(top_core_KE_new_sboxw_17_), .B(top_core_KE_n2024), .Y(
        top_core_KE_n1469) );
  XNOR2X1 U18256 ( .A(top_core_KE_new_sboxw_20_), .B(top_core_KE_n2015), .Y(
        top_core_KE_n1445) );
  XNOR2X1 U18257 ( .A(top_core_KE_new_sboxw_19_), .B(top_core_KE_n2018), .Y(
        top_core_KE_n1453) );
  AOI2BB2X1 U18258 ( .B0(n1798), .B1(n11914), .A0N(n11675), .A1N(n689), .Y(
        n11912) );
  OAI22XL U18259 ( .A0(n613), .A1(n77), .B0(n1811), .B1(n11779), .Y(n11914) );
  AOI2BB2X1 U18260 ( .B0(n1819), .B1(top_core_KE_sb1_n343), .A0N(
        top_core_KE_sb1_n100), .A1N(n690), .Y(top_core_KE_sb1_n341) );
  OAI22XL U18261 ( .A0(n614), .A1(n78), .B0(n1832), .B1(top_core_KE_sb1_n207), 
        .Y(top_core_KE_sb1_n343) );
  AOI2BB2X1 U18262 ( .B0(n1755), .B1(n12545), .A0N(n12306), .A1N(n691), .Y(
        n12543) );
  OAI22XL U18263 ( .A0(n601), .A1(n184), .B0(n1770), .B1(n12410), .Y(n12545)
         );
  AOI2BB2X1 U18264 ( .B0(n1777), .B1(n12230), .A0N(n11991), .A1N(n693), .Y(
        n12228) );
  OAI22XL U18265 ( .A0(n615), .A1(n79), .B0(n1790), .B1(n12095), .Y(n12230) );
  AOI2BB2X1 U18266 ( .B0(n1639), .B1(n13805), .A0N(n13567), .A1N(n695), .Y(
        n13803) );
  OAI22XL U18267 ( .A0(n1179), .A1(n183), .B0(n1660), .B1(n6), .Y(n13805) );
  CLKINVX3 U18268 ( .A(n1638), .Y(n1635) );
  INVX1 U18269 ( .A(top_core_KE_n883), .Y(n7013) );
  CLKINVX3 U18270 ( .A(n1649), .Y(n1643) );
  NAND4X1 U18271 ( .A(n12387), .B(n12388), .C(n12389), .D(n12390), .Y(n12386)
         );
  AOI21X1 U18272 ( .A0(n6530), .A1(n12396), .B0(n6528), .Y(n12389) );
  OAI22X1 U18273 ( .A0(n12393), .A1(n1752), .B0(n1754), .B1(n12394), .Y(n12391) );
  NAND4X1 U18274 ( .A(n13333), .B(n13334), .C(n13335), .D(n13336), .Y(n13332)
         );
  AOI21X1 U18275 ( .A0(n6472), .A1(n13342), .B0(n6470), .Y(n13335) );
  OAI22X1 U18276 ( .A0(n13339), .A1(n1668), .B0(n1666), .B1(n13340), .Y(n13337) );
  NAND4X1 U18277 ( .A(n12703), .B(n12704), .C(n12705), .D(n12706), .Y(n12702)
         );
  AOI21X1 U18278 ( .A0(n6775), .A1(n12712), .B0(n6773), .Y(n12705) );
  OAI22X1 U18279 ( .A0(n12709), .A1(n1726), .B0(n1724), .B1(n12710), .Y(n12707) );
  NAND4X1 U18280 ( .A(n13648), .B(n13649), .C(n13650), .D(n13651), .Y(n13647)
         );
  AOI21X1 U18281 ( .A0(n6519), .A1(n13657), .B0(n6517), .Y(n13650) );
  OAI22X1 U18282 ( .A0(n13654), .A1(n1635), .B0(n1637), .B1(n13655), .Y(n13652) );
  NAND4X1 U18283 ( .A(n13018), .B(n13019), .C(n13020), .D(n13021), .Y(n13017)
         );
  AOI21X1 U18284 ( .A0(n6815), .A1(n13027), .B0(n6813), .Y(n13020) );
  OAI22X1 U18285 ( .A0(n13024), .A1(n1697), .B0(n1695), .B1(n13025), .Y(n13022) );
  OAI2BB2X1 U18286 ( .B0(n607), .B1(n12437), .A0N(n1265), .A1N(n12442), .Y(
        n12447) );
  OAI2BB2X1 U18287 ( .B0(n605), .B1(n11806), .A0N(n1258), .A1N(n11811), .Y(
        n11816) );
  OAI2BB2X1 U18288 ( .B0(n606), .B1(top_core_KE_sb1_n234), .A0N(n1330), .A1N(
        top_core_KE_sb1_n239), .Y(top_core_KE_sb1_n244) );
  OAI2BB2X1 U18289 ( .B0(n608), .B1(n12122), .A0N(n1261), .A1N(n12127), .Y(
        n12132) );
  INVX1 U18290 ( .A(n1505), .Y(n5386) );
  INVX1 U18291 ( .A(n1529), .Y(n5032) );
  INVX1 U18292 ( .A(n1519), .Y(n5858) );
  INVX1 U18293 ( .A(n1517), .Y(n6170) );
  INVX1 U18294 ( .A(n1531), .Y(n5116) );
  INVX1 U18295 ( .A(n1527), .Y(n6086) );
  INVX1 U18296 ( .A(n1512), .Y(n5622) );
  INVX1 U18297 ( .A(n1503), .Y(n5302) );
  INVX1 U18298 ( .A(n1510), .Y(n5546) );
  INVX1 U18299 ( .A(n1516), .Y(n5774) );
  INVX1 U18300 ( .A(n1523), .Y(n6010) );
  INVX1 U18301 ( .A(n1526), .Y(n4916) );
  INVX1 U18302 ( .A(n1501), .Y(n5224) );
  INVX1 U18303 ( .A(n1508), .Y(n5470) );
  INVX1 U18304 ( .A(n1514), .Y(n5698) );
  INVX1 U18305 ( .A(n1521), .Y(n5934) );
  OAI2BB2X1 U18306 ( .B0(n12806), .B1(n12677), .A0N(n12807), .A1N(n6763), .Y(
        n12805) );
  AOI211X1 U18307 ( .A0(n6851), .A1(n1740), .B0(n12811), .C0(n12812), .Y(
        n12806) );
  NAND4BXL U18308 ( .AN(n12808), .B(n12809), .C(n12754), .D(n12733), .Y(n12807) );
  OAI21XL U18309 ( .A0(n12813), .A1(n12638), .B0(n12814), .Y(n12812) );
  OAI2BB2X1 U18310 ( .B0(n13121), .B1(n12992), .A0N(n13122), .A1N(n6706), .Y(
        n13120) );
  AOI211X1 U18311 ( .A0(n6897), .A1(n1711), .B0(n13126), .C0(n13127), .Y(
        n13121) );
  NAND4BXL U18312 ( .AN(n13123), .B(n13124), .C(n13069), .D(n13048), .Y(n13122) );
  OAI21XL U18313 ( .A0(n13128), .A1(n12953), .B0(n13129), .Y(n13127) );
  OAI2BB2X1 U18314 ( .B0(n13751), .B1(n13622), .A0N(n13752), .A1N(n6419), .Y(
        n13750) );
  AOI211X1 U18315 ( .A0(n6604), .A1(n1654), .B0(n13756), .C0(n13757), .Y(
        n13751) );
  NAND4BXL U18316 ( .AN(n13753), .B(n13754), .C(n13699), .D(n13678), .Y(n13752) );
  OAI21XL U18317 ( .A0(n13758), .A1(n13583), .B0(n13759), .Y(n13757) );
  OAI2BB2X1 U18318 ( .B0(n12491), .B1(n12361), .A0N(n12492), .A1N(n6439), .Y(
        n12490) );
  AOI211X1 U18319 ( .A0(n6627), .A1(n1765), .B0(n12496), .C0(n12497), .Y(
        n12491) );
  NAND4BXL U18320 ( .AN(n12493), .B(n12494), .C(n12439), .D(n12418), .Y(n12492) );
  OAI21XL U18321 ( .A0(n12498), .A1(n12322), .B0(n12499), .Y(n12497) );
  OAI2BB2X1 U18322 ( .B0(n11860), .B1(n11730), .A0N(n11861), .A1N(n6731), .Y(
        n11859) );
  AOI211X1 U18323 ( .A0(n6920), .A1(n1808), .B0(n11865), .C0(n11866), .Y(
        n11860) );
  NAND4BXL U18324 ( .AN(n11862), .B(n11863), .C(n11808), .D(n11787), .Y(n11861) );
  OAI21XL U18325 ( .A0(n11867), .A1(n11691), .B0(n11868), .Y(n11866) );
  OAI2BB2X1 U18326 ( .B0(top_core_KE_sb1_n289), .B1(top_core_KE_sb1_n157), 
        .A0N(top_core_KE_sb1_n290), .A1N(n6794), .Y(top_core_KE_sb1_n288) );
  AOI211X1 U18327 ( .A0(n6874), .A1(n1829), .B0(top_core_KE_sb1_n294), .C0(
        top_core_KE_sb1_n295), .Y(top_core_KE_sb1_n289) );
  NAND4BXL U18328 ( .AN(top_core_KE_sb1_n291), .B(top_core_KE_sb1_n292), .C(
        top_core_KE_sb1_n236), .D(top_core_KE_sb1_n215), .Y(
        top_core_KE_sb1_n290) );
  OAI21XL U18329 ( .A0(top_core_KE_sb1_n296), .A1(top_core_KE_sb1_n116), .B0(
        top_core_KE_sb1_n297), .Y(top_core_KE_sb1_n295) );
  OAI2BB2X1 U18330 ( .B0(n12176), .B1(n12046), .A0N(n12177), .A1N(n6495), .Y(
        n12175) );
  AOI211X1 U18331 ( .A0(n6580), .A1(n1787), .B0(n12181), .C0(n12182), .Y(
        n12176) );
  NAND4BXL U18332 ( .AN(n12178), .B(n12179), .C(n12124), .D(n12103), .Y(n12177) );
  OAI21XL U18333 ( .A0(n12183), .A1(n12007), .B0(n12184), .Y(n12182) );
  NAND4X1 U18334 ( .A(n13383), .B(n13384), .C(n13385), .D(n13386), .Y(n13378)
         );
  NAND4X1 U18335 ( .A(n11657), .B(n11706), .C(n11707), .D(n11708), .Y(n11696)
         );
  AOI22XL U18336 ( .A0(n11709), .A1(n50), .B0(n6909), .B1(n673), .Y(n11707) );
  NAND4X1 U18337 ( .A(top_core_KE_sb1_n82), .B(top_core_KE_sb1_n131), .C(
        top_core_KE_sb1_n132), .D(top_core_KE_sb1_n133), .Y(
        top_core_KE_sb1_n121) );
  AOI22XL U18338 ( .A0(top_core_KE_sb1_n134), .A1(n51), .B0(n6863), .B1(n674), 
        .Y(top_core_KE_sb1_n132) );
  NAND4X1 U18339 ( .A(n12289), .B(n12337), .C(n12338), .D(n12339), .Y(n12327)
         );
  AOI22XL U18340 ( .A0(n12340), .A1(n89), .B0(n6616), .B1(n675), .Y(n12338) );
  NAND4X1 U18341 ( .A(n11973), .B(n12022), .C(n12023), .D(n12024), .Y(n12012)
         );
  AOI22XL U18342 ( .A0(n12025), .A1(n53), .B0(n6569), .B1(n676), .Y(n12023) );
  AOI21XL U18343 ( .A0(n77), .A1(n11673), .B0(n1800), .Y(n11829) );
  AOI21XL U18344 ( .A0(n78), .A1(top_core_KE_sb1_n98), .B0(n1821), .Y(
        top_core_KE_sb1_n258) );
  AOI21XL U18345 ( .A0(n184), .A1(n12304), .B0(n1755), .Y(n12460) );
  AOI21XL U18346 ( .A0(n79), .A1(n11989), .B0(n1779), .Y(n12145) );
  AOI21XL U18347 ( .A0(n183), .A1(n13565), .B0(n1637), .Y(n13720) );
  AOI21X1 U18348 ( .A0(n13590), .A1(n13591), .B0(n13592), .Y(n13589) );
  AOI211X1 U18349 ( .A0(n13593), .A1(n1662), .B0(n13594), .C0(n13595), .Y(
        n13591) );
  AOI21X1 U18350 ( .A0(n11698), .A1(n11699), .B0(n11700), .Y(n11697) );
  AOI211X1 U18351 ( .A0(n11701), .A1(n1812), .B0(n11702), .C0(n11703), .Y(
        n11699) );
  AOI21X1 U18352 ( .A0(top_core_KE_sb1_n123), .A1(top_core_KE_sb1_n124), .B0(
        top_core_KE_sb1_n125), .Y(top_core_KE_sb1_n122) );
  AOI211X1 U18353 ( .A0(top_core_KE_sb1_n126), .A1(n1833), .B0(
        top_core_KE_sb1_n127), .C0(top_core_KE_sb1_n128), .Y(
        top_core_KE_sb1_n124) );
  AOI21X1 U18354 ( .A0(n12329), .A1(n12330), .B0(n12331), .Y(n12328) );
  AOI211X1 U18355 ( .A0(n12332), .A1(n1772), .B0(n12333), .C0(n12334), .Y(
        n12330) );
  AOI21X1 U18356 ( .A0(n12014), .A1(n12015), .B0(n12016), .Y(n12013) );
  AOI211X1 U18357 ( .A0(n12017), .A1(n1791), .B0(n12018), .C0(n12019), .Y(
        n12015) );
  AOI21X1 U18358 ( .A0(n13275), .A1(n13276), .B0(n13277), .Y(n13274) );
  AOI211X1 U18359 ( .A0(n13278), .A1(n1693), .B0(n13279), .C0(n13280), .Y(
        n13276) );
  AOI21X1 U18360 ( .A0(n12645), .A1(n12646), .B0(n12647), .Y(n12644) );
  AOI211X1 U18361 ( .A0(n12648), .A1(n1751), .B0(n12649), .C0(n12650), .Y(
        n12646) );
  AOI21X1 U18362 ( .A0(n12960), .A1(n12961), .B0(n12962), .Y(n12959) );
  AOI211X1 U18363 ( .A0(n12963), .A1(n1722), .B0(n12964), .C0(n12965), .Y(
        n12961) );
  OAI21XL U18364 ( .A0(n13511), .A1(n1669), .B0(n13512), .Y(n13510) );
  NOR4BX1 U18365 ( .AN(n13513), .B(n13514), .C(n6556), .D(n13258), .Y(n13511)
         );
  AOI31X1 U18366 ( .A0(n6472), .A1(n1166), .A2(n670), .B0(n6471), .Y(n13512)
         );
  CLKINVX3 U18367 ( .A(n2336), .Y(n2330) );
  CLKINVX3 U18368 ( .A(top_core_KE_prev_key1_reg_13_), .Y(n1795) );
  CLKINVX3 U18369 ( .A(top_core_KE_prev_key1_reg_5_), .Y(n1816) );
  CLKINVX3 U18370 ( .A(top_core_KE_prev_key1_reg_21_), .Y(n1774) );
  CLKINVX3 U18371 ( .A(n2336), .Y(n2333) );
  CLKINVX3 U18372 ( .A(n2335), .Y(n2332) );
  CLKINVX3 U18373 ( .A(n2335), .Y(n2331) );
  CLKINVX3 U18374 ( .A(n1758), .Y(n1752) );
  AOI21X1 U18375 ( .A0(n11830), .A1(n11831), .B0(n1795), .Y(n11828) );
  AOI211X1 U18376 ( .A0(n6909), .A1(n1803), .B0(n11741), .C0(n11832), .Y(
        n11831) );
  AOI21X1 U18377 ( .A0(n11716), .A1(n11706), .B0(n577), .Y(n11832) );
  AOI21X1 U18378 ( .A0(top_core_KE_sb1_n259), .A1(top_core_KE_sb1_n260), .B0(
        n1816), .Y(top_core_KE_sb1_n257) );
  AOI211X1 U18379 ( .A0(n6863), .A1(n1824), .B0(top_core_KE_sb1_n168), .C0(
        top_core_KE_sb1_n261), .Y(top_core_KE_sb1_n260) );
  AOI21X1 U18380 ( .A0(top_core_KE_sb1_n143), .A1(top_core_KE_sb1_n131), .B0(
        n578), .Y(top_core_KE_sb1_n261) );
  AOI21X1 U18381 ( .A0(n12146), .A1(n12147), .B0(n1774), .Y(n12144) );
  AOI211X1 U18382 ( .A0(n6569), .A1(n1782), .B0(n12057), .C0(n12148), .Y(
        n12147) );
  AOI21X1 U18383 ( .A0(n12032), .A1(n12022), .B0(n581), .Y(n12148) );
  AOI21X1 U18384 ( .A0(n12461), .A1(n12462), .B0(n1752), .Y(n12459) );
  AOI211X1 U18385 ( .A0(n6616), .A1(n1761), .B0(n12372), .C0(n12463), .Y(
        n12462) );
  AOI21X1 U18386 ( .A0(n12347), .A1(n12337), .B0(n579), .Y(n12463) );
  NAND4X1 U18387 ( .A(n11734), .B(n11787), .C(n11657), .D(n11869), .Y(n11858)
         );
  AOI32XL U18388 ( .A0(n11778), .A1(n1211), .A2(n681), .B0(n11797), .B1(n1221), 
        .Y(n11869) );
  NAND4X1 U18389 ( .A(top_core_KE_sb1_n161), .B(top_core_KE_sb1_n215), .C(
        top_core_KE_sb1_n82), .D(top_core_KE_sb1_n298), .Y(
        top_core_KE_sb1_n287) );
  AOI32XL U18390 ( .A0(top_core_KE_sb1_n206), .A1(n1210), .A2(n682), .B0(
        top_core_KE_sb1_n225), .B1(n1215), .Y(top_core_KE_sb1_n298) );
  NAND4X1 U18391 ( .A(n12365), .B(n12418), .C(n12289), .D(n12500), .Y(n12489)
         );
  AOI32XL U18392 ( .A0(n12409), .A1(n1171), .A2(n683), .B0(n12428), .B1(n1183), 
        .Y(n12500) );
  NAND4X1 U18393 ( .A(n12050), .B(n12103), .C(n11973), .D(n12185), .Y(n12174)
         );
  AOI32XL U18394 ( .A0(n12094), .A1(n1170), .A2(n684), .B0(n12113), .B1(n1175), 
        .Y(n12185) );
  NAND4X1 U18395 ( .A(n12681), .B(n12733), .C(n12604), .D(n12815), .Y(n12804)
         );
  AOI32XL U18396 ( .A0(n12725), .A1(n1737), .A2(n671), .B0(n12743), .B1(n1212), 
        .Y(n12815) );
  NAND4X1 U18397 ( .A(n13626), .B(n13678), .C(n13549), .D(n13760), .Y(n13749)
         );
  AOI32XL U18398 ( .A0(n13670), .A1(n1644), .A2(n669), .B0(n13688), .B1(n1180), 
        .Y(n13760) );
  NAND4X1 U18399 ( .A(n12996), .B(n13048), .C(n12919), .D(n13130), .Y(n13119)
         );
  AOI32XL U18400 ( .A0(n13040), .A1(n1708), .A2(n672), .B0(n13058), .B1(n1218), 
        .Y(n13130) );
  CLKINVX3 U18401 ( .A(n3705), .Y(n3688) );
  CLKINVX3 U18402 ( .A(n896), .Y(n3526) );
  NAND4BXL U18403 ( .AN(n12650), .B(n12681), .C(n12816), .D(n12817), .Y(n12803) );
  AOI22X1 U18404 ( .A0(n12743), .A1(n584), .B0(n6928), .B1(n1731), .Y(n12816)
         );
  NAND4BXL U18405 ( .AN(n13595), .B(n13626), .C(n13761), .D(n13762), .Y(n13748) );
  AOI22X1 U18406 ( .A0(n13688), .A1(n583), .B0(n6653), .B1(n1645), .Y(n13761)
         );
  NAND4BXL U18407 ( .AN(n12965), .B(n12996), .C(n13131), .D(n13132), .Y(n13118) );
  AOI22X1 U18408 ( .A0(n13058), .A1(n582), .B0(n6943), .B1(n1702), .Y(n13131)
         );
  NAND4X1 U18409 ( .A(n12289), .B(n12290), .C(n12291), .D(n12292), .Y(n12266)
         );
  AOI21X1 U18410 ( .A0(n12294), .A1(n1767), .B0(n12295), .Y(n12291) );
  NAND4X1 U18411 ( .A(n13549), .B(n13550), .C(n13551), .D(n13552), .Y(n13526)
         );
  AOI21X1 U18412 ( .A0(n13555), .A1(n1658), .B0(n13556), .Y(n13551) );
  NAND4X1 U18413 ( .A(n11657), .B(n11658), .C(n11659), .D(n11660), .Y(n11634)
         );
  AOI21X1 U18414 ( .A0(n11663), .A1(n1809), .B0(n11664), .Y(n11659) );
  NAND4X1 U18415 ( .A(top_core_KE_sb1_n82), .B(top_core_KE_sb1_n83), .C(
        top_core_KE_sb1_n84), .D(top_core_KE_sb1_n85), .Y(top_core_KE_sb1_n59)
         );
  AOI21X1 U18416 ( .A0(top_core_KE_sb1_n88), .A1(n1830), .B0(
        top_core_KE_sb1_n89), .Y(top_core_KE_sb1_n84) );
  NAND4X1 U18417 ( .A(n11973), .B(n11974), .C(n11975), .D(n11976), .Y(n11950)
         );
  AOI21X1 U18418 ( .A0(n11979), .A1(n1788), .B0(n11980), .Y(n11975) );
  CLKINVX3 U18419 ( .A(n2336), .Y(n2329) );
  CLKINVX3 U18420 ( .A(n2336), .Y(n2328) );
  CLKINVX3 U18421 ( .A(n2336), .Y(n2327) );
  INVX1 U18422 ( .A(top_core_EC_n950), .Y(n3577) );
  CLKINVX3 U18423 ( .A(n3558), .Y(n3554) );
  CLKINVX3 U18424 ( .A(n3558), .Y(n3555) );
  CLKINVX3 U18425 ( .A(n3558), .Y(n3556) );
  CLKINVX3 U18426 ( .A(n3558), .Y(n3557) );
  NAND4X1 U18427 ( .A(n13234), .B(n13235), .C(n13236), .D(n13237), .Y(n13211)
         );
  AOI21X1 U18428 ( .A0(n13240), .A1(n1687), .B0(n13241), .Y(n13236) );
  NAND4X1 U18429 ( .A(n12919), .B(n12920), .C(n12921), .D(n12922), .Y(n12896)
         );
  AOI21X1 U18430 ( .A0(n12925), .A1(n1716), .B0(n12926), .Y(n12921) );
  NAND4X1 U18431 ( .A(n12604), .B(n12605), .C(n12606), .D(n12607), .Y(n12581)
         );
  AOI21X1 U18432 ( .A0(n12610), .A1(n1745), .B0(n12611), .Y(n12606) );
  INVX1 U18433 ( .A(top_core_EC_n951), .Y(n3581) );
  AOI222X1 U18434 ( .A0(n1149), .A1(n1173), .B0(n6554), .B1(n677), .C0(n610), 
        .C1(n1151), .Y(n13483) );
  AOI222X1 U18435 ( .A0(n1189), .A1(n1213), .B0(n6849), .B1(n678), .C0(n611), 
        .C1(n1191), .Y(n12853) );
  NAND4X1 U18436 ( .A(n11756), .B(n11669), .C(n11906), .D(n11907), .Y(n11905)
         );
  AOI222X1 U18437 ( .A0(n1203), .A1(n1222), .B0(n6919), .B1(n673), .C0(n1223), 
        .C1(n745), .Y(n11907) );
  NAND4X1 U18438 ( .A(top_core_KE_sb1_n184), .B(top_core_KE_sb1_n94), .C(
        top_core_KE_sb1_n335), .D(top_core_KE_sb1_n336), .Y(
        top_core_KE_sb1_n334) );
  AOI222X1 U18439 ( .A0(n1194), .A1(n1216), .B0(n6873), .B1(n674), .C0(n1217), 
        .C1(n746), .Y(top_core_KE_sb1_n336) );
  NAND4X1 U18440 ( .A(n12387), .B(n12300), .C(n12537), .D(n12538), .Y(n12536)
         );
  AOI222X1 U18441 ( .A0(n1163), .A1(n1181), .B0(n6626), .B1(n675), .C0(n1182), 
        .C1(n744), .Y(n12538) );
  AOI222X1 U18442 ( .A0(n1158), .A1(n1178), .B0(n6602), .B1(n679), .C0(n616), 
        .C1(n1160), .Y(n13798) );
  AOI222X1 U18443 ( .A0(n1198), .A1(n1219), .B0(n6895), .B1(n680), .C0(n612), 
        .C1(n1200), .Y(n13168) );
  NAND4X1 U18444 ( .A(n12072), .B(n11985), .C(n12222), .D(n12223), .Y(n12221)
         );
  AOI222X1 U18445 ( .A0(n1154), .A1(n1176), .B0(n6579), .B1(n676), .C0(n1177), 
        .C1(n747), .Y(n12223) );
  CLKINVX3 U18446 ( .A(n3706), .Y(n3687) );
  NAND4BXL U18447 ( .AN(n11664), .B(n11680), .C(n6922), .D(n11751), .Y(n11748)
         );
  AOI211X1 U18448 ( .A0(n6904), .A1(n1223), .B0(n6950), .C0(n11752), .Y(n11751) );
  INVX1 U18449 ( .A(n11753), .Y(n6950) );
  AOI21XL U18450 ( .A0(n80), .A1(n11706), .B0(n1259), .Y(n11752) );
  NAND4BXL U18451 ( .AN(top_core_KE_sb1_n89), .B(top_core_KE_sb1_n105), .C(
        n6876), .D(top_core_KE_sb1_n179), .Y(top_core_KE_sb1_n176) );
  AOI211X1 U18452 ( .A0(n6858), .A1(n1217), .B0(n6935), .C0(
        top_core_KE_sb1_n180), .Y(top_core_KE_sb1_n179) );
  INVX1 U18453 ( .A(top_core_KE_sb1_n181), .Y(n6935) );
  AOI21XL U18454 ( .A0(n81), .A1(top_core_KE_sb1_n131), .B0(n1331), .Y(
        top_core_KE_sb1_n180) );
  NAND4BXL U18455 ( .AN(n12295), .B(n12311), .C(n6629), .D(n12382), .Y(n12379)
         );
  AOI211X1 U18456 ( .A0(n6611), .A1(n1182), .B0(n6660), .C0(n12383), .Y(n12382) );
  INVX1 U18457 ( .A(n12384), .Y(n6660) );
  AOI21XL U18458 ( .A0(n82), .A1(n12337), .B0(n1266), .Y(n12383) );
  NAND4BXL U18459 ( .AN(n11980), .B(n11996), .C(n6582), .D(n12067), .Y(n12064)
         );
  AOI211X1 U18460 ( .A0(n6564), .A1(n1177), .B0(n6644), .C0(n12068), .Y(n12067) );
  INVX1 U18461 ( .A(n12069), .Y(n6644) );
  AOI21XL U18462 ( .A0(n83), .A1(n12022), .B0(n1262), .Y(n12068) );
  CLKINVX3 U18463 ( .A(n1799), .Y(n1796) );
  CLKINVX3 U18464 ( .A(n1820), .Y(n1817) );
  CLKINVX3 U18465 ( .A(n1778), .Y(n1775) );
  NAND3X1 U18466 ( .A(n11874), .B(n11875), .C(n11876), .Y(n11873) );
  NAND3XL U18467 ( .A(n1259), .B(n11778), .C(n6826), .Y(n11876) );
  NAND3X1 U18468 ( .A(top_core_KE_sb1_n303), .B(top_core_KE_sb1_n304), .C(
        top_core_KE_sb1_n305), .Y(top_core_KE_sb1_n302) );
  NAND3XL U18469 ( .A(n1331), .B(top_core_KE_sb1_n206), .C(n6804), .Y(
        top_core_KE_sb1_n305) );
  NAND3X1 U18470 ( .A(n12505), .B(n12506), .C(n12507), .Y(n12504) );
  NAND3XL U18471 ( .A(n1266), .B(n12409), .C(n6530), .Y(n12507) );
  NAND3X1 U18472 ( .A(n13450), .B(n13451), .C(n13452), .Y(n13449) );
  NAND3XL U18473 ( .A(n13282), .B(n13355), .C(n6472), .Y(n13452) );
  NAND3X1 U18474 ( .A(n12190), .B(n12191), .C(n12192), .Y(n12189) );
  NAND3XL U18475 ( .A(n1262), .B(n12094), .C(n6507), .Y(n12192) );
  NAND3X1 U18476 ( .A(n12820), .B(n12821), .C(n12822), .Y(n12819) );
  NAND3XL U18477 ( .A(n12652), .B(n12725), .C(n6775), .Y(n12822) );
  NAND3X1 U18478 ( .A(n13765), .B(n13766), .C(n13767), .Y(n13764) );
  NAND3XL U18479 ( .A(n13597), .B(n13670), .C(n6519), .Y(n13767) );
  NAND3X1 U18480 ( .A(n13135), .B(n13136), .C(n13137), .Y(n13134) );
  NAND3XL U18481 ( .A(n12967), .B(n13040), .C(n6815), .Y(n13137) );
  BUFX3 U18482 ( .A(n6906), .Y(n1202) );
  INVXL U18483 ( .A(n80), .Y(n6906) );
  BUFX3 U18484 ( .A(n6860), .Y(n1193) );
  INVXL U18485 ( .A(n81), .Y(n6860) );
  BUFX3 U18486 ( .A(n6613), .Y(n1162) );
  INVXL U18487 ( .A(n82), .Y(n6613) );
  BUFX3 U18488 ( .A(n6566), .Y(n1153) );
  INVXL U18489 ( .A(n83), .Y(n6566) );
  BUFX3 U18490 ( .A(n6907), .Y(n1203) );
  INVXL U18491 ( .A(n185), .Y(n6907) );
  BUFX3 U18492 ( .A(n6861), .Y(n1194) );
  INVXL U18493 ( .A(n186), .Y(n6861) );
  BUFX3 U18494 ( .A(n6614), .Y(n1163) );
  INVXL U18495 ( .A(n46), .Y(n6614) );
  BUFX3 U18496 ( .A(n6542), .Y(n1149) );
  INVXL U18497 ( .A(n187), .Y(n6542) );
  BUFX3 U18498 ( .A(n6567), .Y(n1154) );
  INVXL U18499 ( .A(n188), .Y(n6567) );
  BUFX3 U18500 ( .A(n6837), .Y(n1189) );
  INVXL U18501 ( .A(n189), .Y(n6837) );
  BUFX3 U18502 ( .A(n6590), .Y(n1158) );
  INVXL U18503 ( .A(n190), .Y(n6590) );
  BUFX3 U18504 ( .A(n6883), .Y(n1198) );
  INVXL U18505 ( .A(n191), .Y(n6883) );
  CLKINVX3 U18506 ( .A(n3568), .Y(n3564) );
  INVX1 U18507 ( .A(top_core_EC_n947), .Y(n3568) );
  CLKINVX3 U18508 ( .A(n2253), .Y(n2244) );
  BUFX3 U18509 ( .A(top_core_EC_mc_mix_in_4_56_), .Y(n1540) );
  OAI22X1 U18510 ( .A0(n2399), .A1(top_core_EC_ss_n171), .B0(n2372), .B1(n195), 
        .Y(top_core_EC_mc_mix_in_4_56_) );
  BUFX3 U18511 ( .A(top_core_EC_mc_mix_in_4_88_), .Y(n1534) );
  OAI22X1 U18512 ( .A0(n2534), .A1(top_core_EC_ss_n136), .B0(n2374), .B1(n215), 
        .Y(top_core_EC_mc_mix_in_4_88_) );
  BUFX3 U18513 ( .A(top_core_EC_mc_mix_in_8[120]), .Y(n1553) );
  OAI22X1 U18514 ( .A0(n2524), .A1(top_core_EC_ss_n229), .B0(n2368), .B1(n234), 
        .Y(top_core_EC_mc_mix_in_8[120]) );
  BUFX3 U18515 ( .A(top_core_EC_mc_mix_in_4_120_), .Y(n1552) );
  OAI22X1 U18516 ( .A0(n2412), .A1(top_core_EC_ss_n228), .B0(n2368), .B1(n235), 
        .Y(top_core_EC_mc_mix_in_4_120_) );
  BUFX3 U18517 ( .A(top_core_EC_mc_mix_in_8[56]), .Y(n1541) );
  OAI22X1 U18518 ( .A0(n2398), .A1(top_core_EC_ss_n172), .B0(n2372), .B1(n194), 
        .Y(top_core_EC_mc_mix_in_8[56]) );
  BUFX3 U18519 ( .A(top_core_EC_mc_mix_in_8[88]), .Y(n1535) );
  OAI22X1 U18520 ( .A0(n2420), .A1(top_core_EC_ss_n137), .B0(n2374), .B1(n214), 
        .Y(top_core_EC_mc_mix_in_8[88]) );
  BUFX3 U18521 ( .A(n6921), .Y(n1205) );
  INVXL U18522 ( .A(n77), .Y(n6921) );
  BUFX3 U18523 ( .A(n6875), .Y(n1196) );
  INVXL U18524 ( .A(n78), .Y(n6875) );
  BUFX3 U18525 ( .A(n6628), .Y(n1165) );
  INVXL U18526 ( .A(n184), .Y(n6628) );
  BUFX3 U18527 ( .A(n6581), .Y(n1156) );
  INVXL U18528 ( .A(n79), .Y(n6581) );
  CLKINVX3 U18529 ( .A(n1756), .Y(n1753) );
  BUFX3 U18530 ( .A(n6099), .Y(n1132) );
  INVX1 U18531 ( .A(n1506), .Y(n6099) );
  BUFX3 U18532 ( .A(n5315), .Y(n992) );
  INVX1 U18533 ( .A(n1504), .Y(n5315) );
  BUFX3 U18534 ( .A(n4961), .Y(n936) );
  INVX1 U18535 ( .A(n1528), .Y(n4961) );
  BUFX3 U18536 ( .A(n5787), .Y(n1076) );
  INVX1 U18537 ( .A(n1518), .Y(n5787) );
  BUFX3 U18538 ( .A(n5477), .Y(n1020) );
  INVX1 U18539 ( .A(n1509), .Y(n5477) );
  BUFX3 U18540 ( .A(n5044), .Y(n950) );
  INVX1 U18541 ( .A(n1530), .Y(n5044) );
  BUFX3 U18542 ( .A(n5705), .Y(n1062) );
  INVX1 U18543 ( .A(n1515), .Y(n5705) );
  BUFX3 U18544 ( .A(n5941), .Y(n1104) );
  INVX1 U18545 ( .A(n1522), .Y(n5941) );
  BUFX3 U18546 ( .A(n5553), .Y(n1034) );
  INVX1 U18547 ( .A(n1511), .Y(n5553) );
  BUFX3 U18548 ( .A(n4842), .Y(n922) );
  INVX1 U18549 ( .A(n1525), .Y(n4842) );
  BUFX3 U18550 ( .A(n5155), .Y(n964) );
  INVX1 U18551 ( .A(n1532), .Y(n5155) );
  BUFX3 U18552 ( .A(n6017), .Y(n1118) );
  INVX1 U18553 ( .A(n1524), .Y(n6017) );
  BUFX3 U18554 ( .A(n5396), .Y(n1006) );
  INVX1 U18555 ( .A(n1507), .Y(n5396) );
  BUFX3 U18556 ( .A(n5629), .Y(n1048) );
  INVX1 U18557 ( .A(n1513), .Y(n5629) );
  BUFX3 U18558 ( .A(n5231), .Y(n978) );
  INVX1 U18559 ( .A(n1502), .Y(n5231) );
  BUFX3 U18560 ( .A(n5865), .Y(n1090) );
  INVX1 U18561 ( .A(n1520), .Y(n5865) );
  BUFX3 U18562 ( .A(top_core_EC_mc_mix_in_4_72_), .Y(n1537) );
  OAI22X1 U18563 ( .A0(n2492), .A1(top_core_EC_ss_n154), .B0(n2373), .B1(n205), 
        .Y(top_core_EC_mc_mix_in_4_72_) );
  BUFX3 U18564 ( .A(top_core_EC_mc_mix_in_4_104_), .Y(n1555) );
  OAI22X1 U18565 ( .A0(n2426), .A1(top_core_EC_ss_n245), .B0(n2367), .B1(n225), 
        .Y(top_core_EC_mc_mix_in_4_104_) );
  BUFX3 U18566 ( .A(top_core_EC_mc_mix_in_8[104]), .Y(n1556) );
  OAI22X1 U18567 ( .A0(n2436), .A1(top_core_EC_ss_n247), .B0(n2367), .B1(n224), 
        .Y(top_core_EC_mc_mix_in_8[104]) );
  BUFX3 U18568 ( .A(top_core_EC_mc_mix_in_8[72]), .Y(n1538) );
  OAI22X1 U18569 ( .A0(n2491), .A1(top_core_EC_ss_n155), .B0(n2373), .B1(n204), 
        .Y(top_core_EC_mc_mix_in_8[72]) );
  BUFX3 U18570 ( .A(n6964), .Y(n1211) );
  BUFX3 U18571 ( .A(n6958), .Y(n1210) );
  BUFX3 U18572 ( .A(n6670), .Y(n1170) );
  XNOR2X1 U18573 ( .A(top_core_KE_new_sboxw_192_2_), .B(top_core_KE_n2288), 
        .Y(top_core_KE_n2287) );
  XNOR2X1 U18574 ( .A(top_core_KE_new_sboxw_192_26_), .B(top_core_KE_n2328), 
        .Y(top_core_KE_n2327) );
  XNOR2X1 U18575 ( .A(top_core_KE_new_sboxw_192_5_), .B(top_core_KE_n2273), 
        .Y(top_core_KE_n2272) );
  XNOR2X1 U18576 ( .A(top_core_KE_new_sboxw_192_29_), .B(top_core_KE_n2313), 
        .Y(top_core_KE_n2312) );
  XNOR2X1 U18577 ( .A(top_core_KE_new_sboxw_192_10_), .B(top_core_KE_n2248), 
        .Y(top_core_KE_n2247) );
  XNOR2X1 U18578 ( .A(top_core_KE_new_sboxw_192_13_), .B(top_core_KE_n2233), 
        .Y(top_core_KE_n2232) );
  XNOR2X1 U18579 ( .A(top_core_KE_new_sboxw_192_15_), .B(top_core_KE_n2223), 
        .Y(top_core_KE_n2222) );
  XNOR2X1 U18580 ( .A(top_core_KE_new_sboxw_192_31_), .B(top_core_KE_n2303), 
        .Y(top_core_KE_n2302) );
  XNOR2X1 U18581 ( .A(top_core_KE_new_sboxw_192_7_), .B(top_core_KE_n2263), 
        .Y(top_core_KE_n2262) );
  INVX1 U18582 ( .A(top_core_KE_n2509), .Y(n7015) );
  BUFX3 U18583 ( .A(top_core_EC_mc_mix_in_2_56_), .Y(n1539) );
  OAI22X1 U18584 ( .A0(n2523), .A1(top_core_EC_ss_n170), .B0(n2372), .B1(n196), 
        .Y(top_core_EC_mc_mix_in_2_56_) );
  BUFX3 U18585 ( .A(top_core_EC_mc_mix_in_2_88_), .Y(n1533) );
  OAI22X1 U18586 ( .A0(n2523), .A1(top_core_EC_ss_n135), .B0(n2374), .B1(n216), 
        .Y(top_core_EC_mc_mix_in_2_88_) );
  BUFX3 U18587 ( .A(top_core_EC_mc_mix_in_2_120_), .Y(n1551) );
  OAI22X1 U18588 ( .A0(n2413), .A1(top_core_EC_ss_n227), .B0(n2368), .B1(n236), 
        .Y(top_core_EC_mc_mix_in_2_120_) );
  INVX1 U18589 ( .A(top_core_KE_n907), .Y(n2170) );
  INVX1 U18590 ( .A(n13319), .Y(n6636) );
  INVX1 U18591 ( .A(n12689), .Y(n6928) );
  INVX1 U18592 ( .A(n13004), .Y(n6943) );
  INVX1 U18593 ( .A(n13634), .Y(n6653) );
  INVX1 U18594 ( .A(n12373), .Y(n6661) );
  INVX1 U18595 ( .A(n11742), .Y(n6951) );
  INVX1 U18596 ( .A(top_core_KE_sb1_n169), .Y(n6936) );
  INVX1 U18597 ( .A(n12058), .Y(n6645) );
  CLKINVX3 U18598 ( .A(n2263), .Y(n2254) );
  CLKINVX3 U18599 ( .A(n2189), .Y(n2180) );
  INVX1 U18600 ( .A(top_core_KE_n910), .Y(n2189) );
  CLKINVX3 U18601 ( .A(n2283), .Y(n2274) );
  INVX1 U18602 ( .A(top_core_KE_n1877), .Y(n2283) );
  INVX1 U18603 ( .A(top_core_EC_add_out_r_1_), .Y(n6102) );
  INVX1 U18604 ( .A(top_core_EC_add_out_r_18_), .Y(n5316) );
  INVX1 U18605 ( .A(top_core_EC_add_out_r_2_), .Y(n6100) );
  INVX1 U18606 ( .A(top_core_EC_add_out_r_34_), .Y(n5788) );
  INVX1 U18607 ( .A(top_core_EC_add_out_r_50_), .Y(n4962) );
  INVX1 U18608 ( .A(top_core_EC_add_out_r_16_), .Y(n5314) );
  INVX1 U18609 ( .A(top_core_EC_add_out_r_0_), .Y(n6095) );
  INVX1 U18610 ( .A(top_core_EC_add_out_r_19_), .Y(n5313) );
  INVX1 U18611 ( .A(top_core_EC_add_out_r_7_), .Y(n6096) );
  INVX1 U18612 ( .A(top_core_EC_add_out_r_3_), .Y(n6098) );
  INVX1 U18613 ( .A(top_core_EC_add_out_r_32_), .Y(n5786) );
  INVX1 U18614 ( .A(top_core_EC_add_out_r_48_), .Y(n4960) );
  INVX1 U18615 ( .A(top_core_EC_add_out_r_51_), .Y(n4959) );
  INVX1 U18616 ( .A(top_core_EC_add_out_r_35_), .Y(n5785) );
  INVX1 U18617 ( .A(top_core_EC_add_out_r_17_), .Y(n5317) );
  INVX1 U18618 ( .A(top_core_EC_add_out_r_10_), .Y(n5045) );
  INVX1 U18619 ( .A(top_core_EC_add_out_r_11_), .Y(n5043) );
  INVX1 U18620 ( .A(top_core_EC_add_out_r_20_), .Y(n5312) );
  INVX1 U18621 ( .A(top_core_EC_add_out_r_4_), .Y(n6094) );
  INVX1 U18622 ( .A(top_core_EC_add_out_r_21_), .Y(n5311) );
  INVX1 U18623 ( .A(top_core_EC_add_out_r_5_), .Y(n6097) );
  INVX1 U18624 ( .A(top_core_EC_add_out_r_22_), .Y(n5310) );
  INVX1 U18625 ( .A(top_core_EC_add_out_r_6_), .Y(n6093) );
  INVX1 U18626 ( .A(top_core_EC_add_out_r_23_), .Y(n5309) );
  INVX1 U18627 ( .A(top_core_EC_add_out_r_49_), .Y(n4963) );
  INVX1 U18628 ( .A(top_core_EC_add_out_r_33_), .Y(n5789) );
  INVX1 U18629 ( .A(top_core_EC_add_out_r_52_), .Y(n4958) );
  INVX1 U18630 ( .A(top_core_EC_add_out_r_53_), .Y(n4957) );
  INVX1 U18631 ( .A(top_core_EC_add_out_r_36_), .Y(n5784) );
  INVX1 U18632 ( .A(top_core_EC_add_out_r_54_), .Y(n4955) );
  INVX1 U18633 ( .A(top_core_EC_add_out_r_37_), .Y(n5783) );
  INVX1 U18634 ( .A(top_core_EC_add_out_r_55_), .Y(n4950) );
  INVX1 U18635 ( .A(top_core_EC_add_out_r_39_), .Y(n5781) );
  INVX1 U18636 ( .A(top_core_EC_add_out_r_38_), .Y(n5782) );
  INVX1 U18637 ( .A(top_core_EC_add_out_r_15_), .Y(n5039) );
  INVX1 U18638 ( .A(top_core_EC_add_out_r_8_), .Y(n5047) );
  INVX1 U18639 ( .A(top_core_EC_add_out_r_13_), .Y(n5041) );
  INVX1 U18640 ( .A(top_core_EC_add_out_r_14_), .Y(n5040) );
  INVX1 U18641 ( .A(top_core_EC_add_out_r_31_), .Y(n4845) );
  INVX1 U18642 ( .A(top_core_EC_add_out_r_29_), .Y(n4846) );
  INVX1 U18643 ( .A(top_core_EC_add_out_r_30_), .Y(n4832) );
  INVX1 U18644 ( .A(top_core_EC_add_out_r_47_), .Y(n5399) );
  INVX1 U18645 ( .A(top_core_EC_add_out_r_40_), .Y(n5395) );
  INVX1 U18646 ( .A(top_core_EC_add_out_r_42_), .Y(n5402) );
  INVX1 U18647 ( .A(top_core_EC_add_out_r_43_), .Y(n5401) );
  INVX1 U18648 ( .A(top_core_EC_add_out_r_45_), .Y(n5400) );
  INVX1 U18649 ( .A(top_core_EC_add_out_r_46_), .Y(n5393) );
  INVX1 U18650 ( .A(top_core_EC_add_out_r_24_), .Y(n4841) );
  INVX1 U18651 ( .A(top_core_EC_add_out_r_26_), .Y(n4848) );
  INVX1 U18652 ( .A(top_core_EC_add_out_r_27_), .Y(n4847) );
  INVX1 U18653 ( .A(top_core_EC_add_out_r_9_), .Y(n5046) );
  INVX1 U18654 ( .A(top_core_EC_add_out_r_12_), .Y(n5042) );
  INVX1 U18655 ( .A(top_core_EC_add_out_r_25_), .Y(n4850) );
  INVX1 U18656 ( .A(top_core_EC_add_out_r_28_), .Y(n4836) );
  INVX1 U18657 ( .A(top_core_EC_add_out_r_56_), .Y(n5233) );
  INVX1 U18658 ( .A(top_core_EC_add_out_r_41_), .Y(n5404) );
  INVX1 U18659 ( .A(top_core_EC_add_out_r_44_), .Y(n5394) );
  INVX1 U18660 ( .A(top_core_EC_add_out_r_57_), .Y(n5232) );
  CLKINVX3 U18661 ( .A(n1639), .Y(n1636) );
  BUFX3 U18662 ( .A(top_core_KE_n2707), .Y(n1500) );
  AOI21X1 U18663 ( .A0(n2140), .A1(n2198), .B0(top_core_KE_n2696), .Y(
        top_core_KE_n2707) );
  BUFX3 U18664 ( .A(top_core_EC_mc_mix_in_2_72_), .Y(n1536) );
  OAI22X1 U18665 ( .A0(n2487), .A1(top_core_EC_ss_n153), .B0(n2373), .B1(n206), 
        .Y(top_core_EC_mc_mix_in_2_72_) );
  BUFX3 U18666 ( .A(top_core_EC_mc_mix_in_2_104_), .Y(n1554) );
  OAI22X1 U18667 ( .A0(n2426), .A1(top_core_EC_ss_n244), .B0(n2370), .B1(n226), 
        .Y(top_core_EC_mc_mix_in_2_104_) );
  XNOR2X1 U18668 ( .A(top_core_KE_new_sboxw_192_0_), .B(top_core_KE_n2298), 
        .Y(top_core_KE_n2297) );
  XNOR2X1 U18669 ( .A(top_core_KE_new_sboxw_192_24_), .B(top_core_KE_n2338), 
        .Y(top_core_KE_n2337) );
  XNOR2X1 U18670 ( .A(top_core_KE_new_sboxw_192_6_), .B(top_core_KE_n2268), 
        .Y(top_core_KE_n2267) );
  XNOR2X1 U18671 ( .A(top_core_KE_new_sboxw_192_8_), .B(top_core_KE_n2258), 
        .Y(top_core_KE_n2257) );
  XNOR2X1 U18672 ( .A(top_core_KE_new_sboxw_192_14_), .B(top_core_KE_n2228), 
        .Y(top_core_KE_n2227) );
  XNOR2X1 U18673 ( .A(top_core_KE_new_sboxw_192_30_), .B(top_core_KE_n2308), 
        .Y(top_core_KE_n2307) );
  XNOR2X1 U18674 ( .A(top_core_KE_new_sboxw_192_1_), .B(top_core_KE_n2293), 
        .Y(top_core_KE_n2292) );
  XNOR2X1 U18675 ( .A(top_core_KE_new_sboxw_192_25_), .B(top_core_KE_n2333), 
        .Y(top_core_KE_n2332) );
  XNOR2X1 U18676 ( .A(top_core_KE_new_sboxw_192_9_), .B(top_core_KE_n2253), 
        .Y(top_core_KE_n2252) );
  XNOR2X1 U18677 ( .A(top_core_KE_new_sboxw_192_3_), .B(top_core_KE_n2283), 
        .Y(top_core_KE_n2282) );
  XNOR2X1 U18678 ( .A(top_core_KE_new_sboxw_192_27_), .B(top_core_KE_n2323), 
        .Y(top_core_KE_n2322) );
  XNOR2X1 U18679 ( .A(top_core_KE_new_sboxw_192_4_), .B(top_core_KE_n2278), 
        .Y(top_core_KE_n2277) );
  XNOR2X1 U18680 ( .A(top_core_KE_new_sboxw_192_28_), .B(top_core_KE_n2318), 
        .Y(top_core_KE_n2317) );
  XNOR2X1 U18681 ( .A(top_core_KE_new_sboxw_192_11_), .B(top_core_KE_n2243), 
        .Y(top_core_KE_n2242) );
  XNOR2X1 U18682 ( .A(top_core_KE_new_sboxw_192_12_), .B(top_core_KE_n2238), 
        .Y(top_core_KE_n2237) );
  XOR2X1 U18683 ( .A(top_core_KE_n2298), .B(top_core_KE_n2466), .Y(
        top_core_KE_n2465) );
  XNOR2X1 U18684 ( .A(top_core_KE_new_sboxw_192_0_), .B(n1716), .Y(
        top_core_KE_n2466) );
  XOR2X1 U18685 ( .A(top_core_KE_n2338), .B(top_core_KE_n2508), .Y(
        top_core_KE_n2507) );
  XNOR2X1 U18686 ( .A(top_core_KE_new_sboxw_192_24_), .B(n1745), .Y(
        top_core_KE_n2508) );
  XOR2X1 U18687 ( .A(top_core_KE_n2293), .B(top_core_KE_n2461), .Y(
        top_core_KE_n2460) );
  XNOR2X1 U18688 ( .A(top_core_KE_new_sboxw_192_1_), .B(n1709), .Y(
        top_core_KE_n2461) );
  XOR2X1 U18689 ( .A(top_core_KE_n2333), .B(top_core_KE_n2501), .Y(
        top_core_KE_n2500) );
  XNOR2X1 U18690 ( .A(top_core_KE_new_sboxw_192_25_), .B(n1738), .Y(
        top_core_KE_n2501) );
  XOR2X1 U18691 ( .A(top_core_KE_n2288), .B(top_core_KE_n2456), .Y(
        top_core_KE_n2455) );
  XNOR2X1 U18692 ( .A(top_core_KE_new_sboxw_192_2_), .B(n1702), .Y(
        top_core_KE_n2456) );
  XOR2X1 U18693 ( .A(top_core_KE_n2328), .B(top_core_KE_n2496), .Y(
        top_core_KE_n2495) );
  XNOR2X1 U18694 ( .A(top_core_KE_new_sboxw_192_26_), .B(n1731), .Y(
        top_core_KE_n2496) );
  XOR2X1 U18695 ( .A(top_core_KE_n2273), .B(top_core_KE_n2441), .Y(
        top_core_KE_n2440) );
  XNOR2X1 U18696 ( .A(top_core_KE_new_sboxw_192_5_), .B(n1695), .Y(
        top_core_KE_n2441) );
  XOR2X1 U18697 ( .A(top_core_KE_n2313), .B(top_core_KE_n2481), .Y(
        top_core_KE_n2480) );
  XNOR2X1 U18698 ( .A(top_core_KE_new_sboxw_192_29_), .B(n1724), .Y(
        top_core_KE_n2481) );
  XOR2X1 U18699 ( .A(top_core_KE_n2258), .B(top_core_KE_n2426), .Y(
        top_core_KE_n2425) );
  XNOR2X1 U18700 ( .A(top_core_KE_new_sboxw_192_8_), .B(n1687), .Y(
        top_core_KE_n2426) );
  XOR2X1 U18701 ( .A(top_core_KE_n2253), .B(top_core_KE_n2421), .Y(
        top_core_KE_n2420) );
  XNOR2X1 U18702 ( .A(top_core_KE_new_sboxw_192_9_), .B(n1680), .Y(
        top_core_KE_n2421) );
  XOR2X1 U18703 ( .A(top_core_KE_n2248), .B(top_core_KE_n2416), .Y(
        top_core_KE_n2415) );
  XNOR2X1 U18704 ( .A(top_core_KE_new_sboxw_192_10_), .B(n1673), .Y(
        top_core_KE_n2416) );
  XOR2X1 U18705 ( .A(top_core_KE_n2233), .B(top_core_KE_n2401), .Y(
        top_core_KE_n2400) );
  XNOR2X1 U18706 ( .A(top_core_KE_new_sboxw_192_13_), .B(n1666), .Y(
        top_core_KE_n2401) );
  AOI222X1 U18707 ( .A0(n6915), .A1(n1810), .B0(n11819), .B1(n665), .C0(n6920), 
        .C1(n1223), .Y(n11931) );
  AOI222X1 U18708 ( .A0(n6869), .A1(n1831), .B0(top_core_KE_sb1_n247), .B1(
        n666), .C0(n6874), .C1(n1217), .Y(top_core_KE_sb1_n360) );
  AOI222X1 U18709 ( .A0(n6622), .A1(n1768), .B0(n12450), .B1(n667), .C0(n6627), 
        .C1(n1182), .Y(n12562) );
  AOI222X1 U18710 ( .A0(n6575), .A1(n1789), .B0(n12135), .B1(n668), .C0(n6580), 
        .C1(n1177), .Y(n12247) );
  AOI222X1 U18711 ( .A0(n6550), .A1(n1688), .B0(n13395), .B1(n670), .C0(n6556), 
        .C1(n610), .Y(n13507) );
  AOI222X1 U18712 ( .A0(n6845), .A1(n1746), .B0(n12765), .B1(n688), .C0(n6851), 
        .C1(n611), .Y(n12877) );
  AOI222X1 U18713 ( .A0(n6598), .A1(n1659), .B0(n13710), .B1(n685), .C0(n6604), 
        .C1(n616), .Y(n13822) );
  AOI222X1 U18714 ( .A0(n6891), .A1(n1717), .B0(n13080), .B1(n687), .C0(n6897), 
        .C1(n612), .Y(n13192) );
  AND2X2 U18715 ( .A(n2866), .B(n1505), .Y(n698) );
  AND2X2 U18716 ( .A(n3467), .B(n1517), .Y(n699) );
  AND2X2 U18717 ( .A(n2624), .B(n1529), .Y(n700) );
  AND2X2 U18718 ( .A(n3226), .B(n1519), .Y(n701) );
  AND2X2 U18719 ( .A(n3165), .B(n1516), .Y(n702) );
  AND2X2 U18720 ( .A(n2927), .B(n1508), .Y(n703) );
  AND2X2 U18721 ( .A(n2563), .B(n1526), .Y(n704) );
  AND2X2 U18722 ( .A(n3287), .B(n1521), .Y(n705) );
  AND2X2 U18723 ( .A(n2988), .B(n1510), .Y(n706) );
  AND2X2 U18724 ( .A(n2685), .B(n1531), .Y(n707) );
  AND2X2 U18725 ( .A(n3348), .B(n1523), .Y(n708) );
  AND2X2 U18726 ( .A(n3046), .B(n1512), .Y(n709) );
  AND2X2 U18727 ( .A(n2745), .B(n1501), .Y(n710) );
  AND2X2 U18728 ( .A(n3406), .B(n1527), .Y(n711) );
  AND2X2 U18729 ( .A(n3107), .B(n1514), .Y(n712) );
  AND2X2 U18730 ( .A(n2806), .B(n1503), .Y(n713) );
  AND2X2 U18731 ( .A(n1505), .B(n2868), .Y(n722) );
  AND2X2 U18732 ( .A(n1517), .B(n3470), .Y(n723) );
  AND2X2 U18733 ( .A(n1529), .B(n2626), .Y(n724) );
  AND2X2 U18734 ( .A(n1519), .B(n3228), .Y(n725) );
  AND2X2 U18735 ( .A(n1516), .B(n3167), .Y(n726) );
  AND2X2 U18736 ( .A(n1508), .B(n2929), .Y(n727) );
  AND2X2 U18737 ( .A(n1526), .B(n2565), .Y(n728) );
  AND2X2 U18738 ( .A(n1521), .B(n3289), .Y(n729) );
  AND2X2 U18739 ( .A(n1510), .B(n2990), .Y(n730) );
  AND2X2 U18740 ( .A(n1531), .B(n2687), .Y(n731) );
  AND2X2 U18741 ( .A(n1523), .B(n3350), .Y(n732) );
  AND2X2 U18742 ( .A(n1512), .B(n3048), .Y(n733) );
  AND2X2 U18743 ( .A(n1501), .B(n2747), .Y(n734) );
  AND2X2 U18744 ( .A(n1527), .B(n3408), .Y(n735) );
  AND2X2 U18745 ( .A(n1514), .B(n3109), .Y(n736) );
  AND2X2 U18746 ( .A(n1503), .B(n2808), .Y(n737) );
  AOI211X1 U18747 ( .A0(n6556), .A1(n1682), .B0(n13441), .C0(n13442), .Y(
        n13436) );
  OAI21XL U18748 ( .A0(n13443), .A1(n13268), .B0(n13444), .Y(n13442) );
  OAI2BB1XL U18749 ( .A0N(n1768), .A1N(n12450), .B0(n184), .Y(n12449) );
  OAI2BB1XL U18750 ( .A0N(n1810), .A1N(n11819), .B0(n77), .Y(n11818) );
  OAI2BB1XL U18751 ( .A0N(n1831), .A1N(top_core_KE_sb1_n247), .B0(n78), .Y(
        top_core_KE_sb1_n246) );
  OAI2BB1XL U18752 ( .A0N(n1789), .A1N(n12135), .B0(n79), .Y(n12134) );
  AOI221X1 U18753 ( .A0(n13272), .A1(n13433), .B0(n6469), .B1(n13434), .C0(
        n13435), .Y(n13432) );
  NAND4BXL U18754 ( .AN(n13280), .B(n13311), .C(n13446), .D(n13447), .Y(n13433) );
  NAND4X1 U18755 ( .A(n13311), .B(n13363), .C(n13234), .D(n13445), .Y(n13434)
         );
  OAI2BB2X1 U18756 ( .B0(n13436), .B1(n13307), .A0N(n13437), .A1N(n6462), .Y(
        n13435) );
  INVX1 U18757 ( .A(n13207), .Y(n6701) );
  INVX1 U18758 ( .A(n12577), .Y(n6988) );
  INVX1 U18759 ( .A(n12892), .Y(n6712) );
  INVX1 U18760 ( .A(n13522), .Y(n6431) );
  INVX1 U18761 ( .A(n12262), .Y(n6372) );
  INVX1 U18762 ( .A(n11630), .Y(n6743) );
  INVX1 U18763 ( .A(top_core_KE_sb1_n55), .Y(n6986) );
  INVX1 U18764 ( .A(n11946), .Y(n6699) );
  AOI222X1 U18765 ( .A0(n6636), .A1(n1674), .B0(n13240), .B1(n686), .C0(n6552), 
        .C1(n1685), .Y(n13474) );
  AOI222X1 U18766 ( .A0(n6928), .A1(n1732), .B0(n12610), .B1(n671), .C0(n6847), 
        .C1(n1743), .Y(n12844) );
  AOI222X1 U18767 ( .A0(n6943), .A1(n1703), .B0(n12925), .B1(n672), .C0(n6893), 
        .C1(n1714), .Y(n13159) );
  AOI222X1 U18768 ( .A0(n6653), .A1(n1647), .B0(n13555), .B1(n669), .C0(n6600), 
        .C1(n1657), .Y(n13789) );
  AOI211X1 U18769 ( .A0(n6920), .A1(n681), .B0(n11900), .C0(n11901), .Y(n11889) );
  OAI21XL U18770 ( .A0(n577), .A1(n11867), .B0(n11902), .Y(n11901) );
  OAI21XL U18771 ( .A0(n6919), .A1(n6914), .B0(n1809), .Y(n11902) );
  AOI211X1 U18772 ( .A0(n6874), .A1(n682), .B0(top_core_KE_sb1_n329), .C0(
        top_core_KE_sb1_n330), .Y(top_core_KE_sb1_n318) );
  OAI21XL U18773 ( .A0(n578), .A1(top_core_KE_sb1_n296), .B0(
        top_core_KE_sb1_n331), .Y(top_core_KE_sb1_n330) );
  OAI21XL U18774 ( .A0(n6873), .A1(n6868), .B0(n1830), .Y(top_core_KE_sb1_n331) );
  AOI211X1 U18775 ( .A0(n6627), .A1(n683), .B0(n12531), .C0(n12532), .Y(n12520) );
  OAI21XL U18776 ( .A0(n579), .A1(n12498), .B0(n12533), .Y(n12532) );
  OAI21XL U18777 ( .A0(n6626), .A1(n6621), .B0(n1768), .Y(n12533) );
  AOI211X1 U18778 ( .A0(n6556), .A1(n686), .B0(n13476), .C0(n13477), .Y(n13465) );
  OAI21XL U18779 ( .A0(n580), .A1(n13443), .B0(n13478), .Y(n13477) );
  OAI21XL U18780 ( .A0(n6554), .A1(n6549), .B0(n1688), .Y(n13478) );
  AOI211X1 U18781 ( .A0(n6580), .A1(n684), .B0(n12216), .C0(n12217), .Y(n12205) );
  OAI21XL U18782 ( .A0(n581), .A1(n12183), .B0(n12218), .Y(n12217) );
  OAI21XL U18783 ( .A0(n6579), .A1(n6574), .B0(n1788), .Y(n12218) );
  AOI211X1 U18784 ( .A0(n6851), .A1(n671), .B0(n12846), .C0(n12847), .Y(n12835) );
  OAI21XL U18785 ( .A0(n584), .A1(n12813), .B0(n12848), .Y(n12847) );
  OAI21XL U18786 ( .A0(n6849), .A1(n6844), .B0(n1746), .Y(n12848) );
  AOI211X1 U18787 ( .A0(n6604), .A1(n669), .B0(n13791), .C0(n13792), .Y(n13780) );
  OAI21XL U18788 ( .A0(n583), .A1(n13758), .B0(n13793), .Y(n13792) );
  OAI21XL U18789 ( .A0(n6602), .A1(n6597), .B0(n1659), .Y(n13793) );
  AOI211X1 U18790 ( .A0(n6897), .A1(n672), .B0(n13161), .C0(n13162), .Y(n13150) );
  OAI21XL U18791 ( .A0(n582), .A1(n13128), .B0(n13163), .Y(n13162) );
  OAI21XL U18792 ( .A0(n6895), .A1(n6890), .B0(n1717), .Y(n13163) );
  AOI211X1 U18793 ( .A0(n1223), .A1(n1204), .B0(n11798), .C0(n1203), .Y(n11793) );
  AOI211X1 U18794 ( .A0(n1217), .A1(n1195), .B0(top_core_KE_sb1_n226), .C0(
        n1194), .Y(top_core_KE_sb1_n221) );
  AOI211X1 U18795 ( .A0(n1182), .A1(n1164), .B0(n12429), .C0(n1163), .Y(n12424) );
  AOI211X1 U18796 ( .A0(n602), .A1(n1150), .B0(n13374), .C0(n1149), .Y(n13369)
         );
  AOI211X1 U18797 ( .A0(n1177), .A1(n1155), .B0(n12114), .C0(n1154), .Y(n12109) );
  AOI211X1 U18798 ( .A0(n603), .A1(n1190), .B0(n12744), .C0(n1189), .Y(n12739)
         );
  AOI211X1 U18799 ( .A0(n609), .A1(n1159), .B0(n13689), .C0(n1158), .Y(n13684)
         );
  AOI211X1 U18800 ( .A0(n604), .A1(n1199), .B0(n13059), .C0(n1198), .Y(n13054)
         );
  AOI211X1 U18801 ( .A0(n6830), .A1(n11894), .B0(n11895), .C0(n11896), .Y(
        n11890) );
  AOI31X1 U18802 ( .A0(n11897), .A1(n11727), .A2(n11898), .B0(n1800), .Y(
        n11895) );
  AOI31X1 U18803 ( .A0(n11757), .A1(n11808), .A2(n11671), .B0(n1796), .Y(
        n11896) );
  AOI211X1 U18804 ( .A0(n6809), .A1(top_core_KE_sb1_n323), .B0(
        top_core_KE_sb1_n324), .C0(top_core_KE_sb1_n325), .Y(
        top_core_KE_sb1_n319) );
  AOI31X1 U18805 ( .A0(top_core_KE_sb1_n326), .A1(top_core_KE_sb1_n154), .A2(
        top_core_KE_sb1_n327), .B0(n1821), .Y(top_core_KE_sb1_n324) );
  AOI31X1 U18806 ( .A0(top_core_KE_sb1_n185), .A1(top_core_KE_sb1_n236), .A2(
        top_core_KE_sb1_n96), .B0(n1817), .Y(top_core_KE_sb1_n325) );
  AOI211X1 U18807 ( .A0(n6534), .A1(n12525), .B0(n12526), .C0(n12527), .Y(
        n12521) );
  AOI31X1 U18808 ( .A0(n12528), .A1(n12358), .A2(n12529), .B0(n1757), .Y(
        n12526) );
  AOI31X1 U18809 ( .A0(n12388), .A1(n12439), .A2(n12302), .B0(n1753), .Y(
        n12527) );
  AOI211X1 U18810 ( .A0(n6477), .A1(n13470), .B0(n13471), .C0(n13472), .Y(
        n13466) );
  AOI31X1 U18811 ( .A0(n13334), .A1(n13384), .A2(n13248), .B0(n1668), .Y(
        n13472) );
  AOI31X1 U18812 ( .A0(n13473), .A1(n13304), .A2(n13474), .B0(n1667), .Y(
        n13471) );
  AOI211X1 U18813 ( .A0(n6512), .A1(n12210), .B0(n12211), .C0(n12212), .Y(
        n12206) );
  AOI31X1 U18814 ( .A0(n12213), .A1(n12043), .A2(n12214), .B0(n1779), .Y(
        n12211) );
  AOI31X1 U18815 ( .A0(n12073), .A1(n12124), .A2(n11987), .B0(n1775), .Y(
        n12212) );
  AOI211X1 U18816 ( .A0(n6780), .A1(n12840), .B0(n12841), .C0(n12842), .Y(
        n12836) );
  AOI31X1 U18817 ( .A0(n12704), .A1(n12754), .A2(n12618), .B0(n1730), .Y(
        n12842) );
  AOI31X1 U18818 ( .A0(n12843), .A1(n12674), .A2(n12844), .B0(n1725), .Y(
        n12841) );
  AOI211X1 U18819 ( .A0(n6523), .A1(n13785), .B0(n13786), .C0(n13787), .Y(
        n13781) );
  AOI31X1 U18820 ( .A0(n13788), .A1(n13619), .A2(n13789), .B0(n1641), .Y(
        n13786) );
  AOI31X1 U18821 ( .A0(n13649), .A1(n13699), .A2(n13563), .B0(n1636), .Y(
        n13787) );
  AOI211X1 U18822 ( .A0(n6819), .A1(n13155), .B0(n13156), .C0(n13157), .Y(
        n13151) );
  AOI31X1 U18823 ( .A0(n13019), .A1(n13069), .A2(n12933), .B0(n1701), .Y(
        n13157) );
  AOI31X1 U18824 ( .A0(n13158), .A1(n12989), .A2(n13159), .B0(n1696), .Y(
        n13156) );
  AOI222X1 U18825 ( .A0(n1801), .A1(n11776), .B0(n11777), .B1(n1796), .C0(
        n1223), .C1(n6824), .Y(n11775) );
  OAI21XL U18826 ( .A0(n11778), .A1(n1258), .B0(n11690), .Y(n11777) );
  OAI211XL U18827 ( .A0(n11779), .A1(n11661), .B0(n11772), .C0(n11780), .Y(
        n11776) );
  AOI222X1 U18828 ( .A0(n1822), .A1(top_core_KE_sb1_n204), .B0(
        top_core_KE_sb1_n205), .B1(n1817), .C0(n1217), .C1(n6802), .Y(
        top_core_KE_sb1_n203) );
  OAI21XL U18829 ( .A0(top_core_KE_sb1_n206), .A1(n1330), .B0(
        top_core_KE_sb1_n115), .Y(top_core_KE_sb1_n205) );
  OAI211XL U18830 ( .A0(top_core_KE_sb1_n207), .A1(top_core_KE_sb1_n86), .B0(
        top_core_KE_sb1_n200), .C0(top_core_KE_sb1_n208), .Y(
        top_core_KE_sb1_n204) );
  AOI222X1 U18831 ( .A0(n1758), .A1(n12407), .B0(n12408), .B1(n1753), .C0(
        n1182), .C1(n6528), .Y(n12406) );
  OAI21XL U18832 ( .A0(n12409), .A1(n1265), .B0(n12321), .Y(n12408) );
  OAI211XL U18833 ( .A0(n12410), .A1(n1264), .B0(n12403), .C0(n12411), .Y(
        n12407) );
  AOI222X1 U18834 ( .A0(n1780), .A1(n12092), .B0(n12093), .B1(n1775), .C0(
        n1177), .C1(n6505), .Y(n12091) );
  OAI21XL U18835 ( .A0(n12094), .A1(n1261), .B0(n12006), .Y(n12093) );
  OAI211XL U18836 ( .A0(n12095), .A1(n11977), .B0(n12088), .C0(n12096), .Y(
        n12092) );
  AOI222X1 U18837 ( .A0(n1641), .A1(n13668), .B0(n13669), .B1(n1636), .C0(n609), .C1(n6517), .Y(n13667) );
  OAI21XL U18838 ( .A0(n13670), .A1(n1277), .B0(n13582), .Y(n13669) );
  AOI222X1 U18839 ( .A0(n1725), .A1(n12723), .B0(n12724), .B1(n1727), .C0(n603), .C1(n6773), .Y(n12722) );
  OAI21XL U18840 ( .A0(n12725), .A1(n1268), .B0(n12637), .Y(n12724) );
  AOI222X1 U18841 ( .A0(n1696), .A1(n13038), .B0(n13039), .B1(n1698), .C0(n604), .C1(n6813), .Y(n13037) );
  OAI21XL U18842 ( .A0(n13040), .A1(n1271), .B0(n12952), .Y(n13039) );
  CLKINVX3 U18843 ( .A(n1648), .Y(n1644) );
  INVX1 U18844 ( .A(top_core_KE_prev_key1_reg_25_), .Y(n1762) );
  INVX1 U18845 ( .A(n13421), .Y(n6468) );
  AOI22X1 U18846 ( .A0(n6475), .A1(n13422), .B0(n6469), .B1(n13423), .Y(n13421) );
  NAND4XL U18847 ( .A(n13383), .B(n13295), .C(n13301), .D(n13424), .Y(n13423)
         );
  NAND4BXL U18848 ( .AN(n13426), .B(n13248), .C(n13363), .D(n13427), .Y(n13422) );
  INVX1 U18849 ( .A(top_core_KE_n1133), .Y(n6339) );
  INVX1 U18850 ( .A(top_core_KE_n1168), .Y(n6370) );
  INVX1 U18851 ( .A(top_core_KE_n1147), .Y(n6362) );
  INVX1 U18852 ( .A(top_core_KE_n1182), .Y(n6356) );
  INVX1 U18853 ( .A(top_core_KE_n1140), .Y(n6348) );
  INVX1 U18854 ( .A(top_core_KE_n1175), .Y(n6312) );
  INVX1 U18855 ( .A(top_core_KE_n1161), .Y(n6366) );
  INVX1 U18856 ( .A(top_core_KE_n1154), .Y(n6352) );
  INVX1 U18857 ( .A(n2335), .Y(n2334) );
  INVX1 U18858 ( .A(n1652), .Y(n1653) );
  INVX1 U18859 ( .A(n1810), .Y(n1811) );
  INVX1 U18860 ( .A(n1831), .Y(n1832) );
  INVX1 U18861 ( .A(n1789), .Y(n1790) );
  INVX1 U18862 ( .A(top_core_KE_prev_key1_reg_88_), .Y(n1660) );
  INVX1 U18863 ( .A(top_core_KE_prev_key1_reg_88_), .Y(n1661) );
  INVX1 U18864 ( .A(top_core_KE_prev_key1_reg_89_), .Y(n1655) );
  INVX1 U18865 ( .A(n1803), .Y(n1804) );
  INVX1 U18866 ( .A(n1824), .Y(n1825) );
  INVX1 U18867 ( .A(n1680), .Y(n1682) );
  INVX1 U18868 ( .A(n1782), .Y(n1783) );
  INVX1 U18869 ( .A(n1738), .Y(n1740) );
  INVX1 U18870 ( .A(n1709), .Y(n1711) );
  INVX1 U18871 ( .A(top_core_KE_prev_key1_reg_9_), .Y(n1805) );
  INVX1 U18872 ( .A(top_core_KE_prev_key1_reg_1_), .Y(n1826) );
  INVX1 U18873 ( .A(top_core_KE_prev_key1_reg_81_), .Y(n1683) );
  INVX1 U18874 ( .A(top_core_KE_prev_key1_reg_17_), .Y(n1784) );
  INVX1 U18875 ( .A(top_core_KE_prev_key1_reg_65_), .Y(n1741) );
  INVX1 U18876 ( .A(top_core_KE_prev_key1_reg_73_), .Y(n1712) );
  INVX1 U18877 ( .A(n1761), .Y(n1763) );
  INVX1 U18878 ( .A(n1810), .Y(n1812) );
  INVX1 U18879 ( .A(n1831), .Y(n1833) );
  INVX1 U18880 ( .A(n1789), .Y(n1791) );
  INVX1 U18881 ( .A(n1666), .Y(n1671) );
  INVX1 U18882 ( .A(n1761), .Y(n1764) );
  INVX1 U18883 ( .A(top_core_KE_prev_key1_reg_24_), .Y(n1769) );
  OR2X2 U18884 ( .A(n7019), .B(n7016), .Y(n738) );
  NOR2BX1 U18885 ( .AN(top_core_EC_n868), .B(n4259), .Y(top_core_EC_n733) );
  NOR2BX1 U18886 ( .AN(top_core_KE_n2693), .B(n2291), .Y(top_core_KE_n2179) );
  OAI22X1 U18887 ( .A0(n1857), .A1(n7021), .B0(n7020), .B1(n1845), .Y(
        top_core_KE_n2693) );
  INVX1 U18888 ( .A(n2365), .Y(n2541) );
  INVX1 U18889 ( .A(n2365), .Y(n2542) );
  INVX1 U18890 ( .A(n2289), .Y(n2284) );
  INVX1 U18891 ( .A(top_core_KE_prev_key1_reg_8_), .Y(n1813) );
  INVX1 U18892 ( .A(top_core_KE_prev_key1_reg_0_), .Y(n1834) );
  INVX1 U18893 ( .A(top_core_KE_prev_key1_reg_80_), .Y(n1689) );
  INVX1 U18894 ( .A(top_core_KE_prev_key1_reg_16_), .Y(n1792) );
  INVX1 U18895 ( .A(top_core_KE_prev_key1_reg_64_), .Y(n1747) );
  INVX1 U18896 ( .A(top_core_KE_prev_key1_reg_72_), .Y(n1718) );
  INVX1 U18897 ( .A(n1724), .Y(n1729) );
  INVX1 U18898 ( .A(n1695), .Y(n1700) );
  INVX1 U18899 ( .A(top_core_KE_prev_key1_reg_89_), .Y(n1656) );
  INVX1 U18900 ( .A(top_core_Addr[2]), .Y(n3985) );
  INVX1 U18901 ( .A(n4088), .Y(n4110) );
  INVX1 U18902 ( .A(top_core_KE_prev_key1_reg_8_), .Y(n1814) );
  INVX1 U18903 ( .A(top_core_KE_prev_key1_reg_0_), .Y(n1835) );
  INVX1 U18904 ( .A(top_core_KE_prev_key1_reg_80_), .Y(n1690) );
  INVX1 U18905 ( .A(top_core_KE_prev_key1_reg_16_), .Y(n1793) );
  INVX1 U18906 ( .A(top_core_KE_prev_key1_reg_72_), .Y(n1719) );
  INVX1 U18907 ( .A(top_core_KE_prev_key1_reg_88_), .Y(n1662) );
  INVX1 U18908 ( .A(top_core_KE_prev_key1_reg_64_), .Y(n1748) );
  INVX1 U18909 ( .A(n1803), .Y(n1806) );
  INVX1 U18910 ( .A(n1824), .Y(n1827) );
  INVX1 U18911 ( .A(n1782), .Y(n1785) );
  INVX1 U18912 ( .A(n1688), .Y(n1691) );
  INVX1 U18913 ( .A(n1746), .Y(n1749) );
  INVX1 U18914 ( .A(top_core_KE_prev_key1_reg_88_), .Y(n1663) );
  INVX1 U18915 ( .A(n1717), .Y(n1720) );
  INVX1 U18916 ( .A(top_core_KE_prev_key1_reg_24_), .Y(n1770) );
  INVX1 U18917 ( .A(top_core_KE_prev_key1_reg_88_), .Y(n1664) );
  INVX1 U18918 ( .A(n1688), .Y(n1692) );
  INVX1 U18919 ( .A(n1717), .Y(n1721) );
  INVX1 U18920 ( .A(n1746), .Y(n1750) );
  INVX1 U18921 ( .A(top_core_KE_prev_key1_reg_8_), .Y(n1815) );
  INVX1 U18922 ( .A(top_core_KE_prev_key1_reg_0_), .Y(n1836) );
  INVX1 U18923 ( .A(top_core_KE_prev_key1_reg_16_), .Y(n1794) );
  INVX1 U18924 ( .A(n1768), .Y(n1771) );
  INVX1 U18925 ( .A(n1674), .Y(n1675) );
  INVX1 U18926 ( .A(n1731), .Y(n1733) );
  INVX1 U18927 ( .A(n1702), .Y(n1704) );
  INVX1 U18928 ( .A(n2540), .Y(n2538) );
  INVX1 U18930 ( .A(n2904), .Y(n2906) );
  INVX1 U18931 ( .A(n3264), .Y(n3266) );
  INVX1 U18932 ( .A(n2722), .Y(n2724) );
  INVX1 U18933 ( .A(n3203), .Y(n3205) );
  INVX1 U18934 ( .A(n2965), .Y(n2967) );
  INVX1 U18935 ( .A(n3444), .Y(n3446) );
  INVX1 U18936 ( .A(top_core_KE_prev_key1_reg_82_), .Y(n1676) );
  INVX1 U18937 ( .A(top_core_KE_prev_key1_reg_66_), .Y(n1734) );
  INVX1 U18938 ( .A(top_core_KE_prev_key1_reg_74_), .Y(n1705) );
  INVX1 U18939 ( .A(top_core_KE_prev_key1_reg_66_), .Y(n1735) );
  INVX1 U18940 ( .A(top_core_KE_prev_key1_reg_74_), .Y(n1706) );
  INVX1 U18941 ( .A(top_core_KE_prev_key1_reg_82_), .Y(n1677) );
  INVX1 U18942 ( .A(top_core_KE_prev_key1_reg_66_), .Y(n1736) );
  INVX1 U18943 ( .A(top_core_KE_prev_key1_reg_74_), .Y(n1707) );
  INVX1 U18944 ( .A(n1768), .Y(n1772) );
  INVX1 U18945 ( .A(top_core_KE_prev_key1_reg_89_), .Y(n1657) );
  INVX1 U18946 ( .A(top_core_KE_n907), .Y(n2169) );
  INVX1 U18947 ( .A(top_core_KE_n910), .Y(n2188) );
  INVX1 U18948 ( .A(top_core_KE_n1877), .Y(n2282) );
  INVX1 U18949 ( .A(top_core_KE_n1875), .Y(n2263) );
  INVX1 U18950 ( .A(top_core_KE_n1875), .Y(n2262) );
  INVX1 U18951 ( .A(top_core_KE_prev_key1_reg_82_), .Y(n1678) );
  INVX1 U18952 ( .A(top_core_KE_prev_key1_reg_66_), .Y(n1737) );
  INVX1 U18953 ( .A(top_core_KE_prev_key1_reg_74_), .Y(n1708) );
  INVX1 U18954 ( .A(top_core_EC_n869), .Y(n3548) );
  INVX1 U18955 ( .A(top_core_KE_n2176), .Y(n2311) );
  INVX1 U18956 ( .A(n1626), .Y(n1634) );
  INVX1 U18957 ( .A(top_core_KE_prev_key1_reg_9_), .Y(n1807) );
  INVX1 U18958 ( .A(top_core_KE_prev_key1_reg_1_), .Y(n1828) );
  INVX1 U18959 ( .A(top_core_KE_prev_key1_reg_81_), .Y(n1684) );
  INVX1 U18960 ( .A(top_core_KE_prev_key1_reg_17_), .Y(n1786) );
  INVX1 U18961 ( .A(top_core_KE_prev_key1_reg_65_), .Y(n1742) );
  INVX1 U18962 ( .A(top_core_KE_prev_key1_reg_73_), .Y(n1713) );
  INVX1 U18963 ( .A(top_core_KE_prev_key1_reg_25_), .Y(n1765) );
  INVX1 U18964 ( .A(top_core_KE_prev_key1_reg_25_), .Y(n1766) );
  INVX1 U18965 ( .A(top_core_KE_prev_key1_reg_81_), .Y(n1685) );
  INVX1 U18966 ( .A(top_core_KE_prev_key1_reg_65_), .Y(n1743) );
  INVX1 U18967 ( .A(top_core_KE_prev_key1_reg_73_), .Y(n1714) );
  INVX1 U18968 ( .A(top_core_KE_prev_key1_reg_24_), .Y(n1773) );
  INVX1 U18969 ( .A(top_core_KE_prev_key1_reg_9_), .Y(n1808) );
  INVX1 U18970 ( .A(top_core_KE_prev_key1_reg_1_), .Y(n1829) );
  INVX1 U18971 ( .A(top_core_KE_prev_key1_reg_81_), .Y(n1686) );
  INVX1 U18972 ( .A(top_core_KE_prev_key1_reg_17_), .Y(n1787) );
  INVX1 U18973 ( .A(top_core_KE_prev_key1_reg_65_), .Y(n1744) );
  INVX1 U18974 ( .A(top_core_KE_prev_key1_reg_73_), .Y(n1715) );
  INVX1 U18975 ( .A(top_core_KE_prev_key1_reg_80_), .Y(n1693) );
  INVX1 U18976 ( .A(top_core_KE_prev_key1_reg_64_), .Y(n1751) );
  INVX1 U18977 ( .A(top_core_KE_prev_key1_reg_72_), .Y(n1722) );
  INVX1 U18978 ( .A(top_core_KE_prev_key1_reg_85_), .Y(n1672) );
  INVX1 U18979 ( .A(top_core_KE_prev_key1_reg_69_), .Y(n1730) );
  INVX1 U18980 ( .A(top_core_KE_prev_key1_reg_77_), .Y(n1701) );
  INVX1 U18981 ( .A(n2366), .Y(n2539) );
  INVX1 U18982 ( .A(n2221), .Y(n2220) );
  INVX1 U18984 ( .A(n4033), .Y(n4115) );
  INVX1 U18985 ( .A(n4032), .Y(n4112) );
  INVX1 U18986 ( .A(n4032), .Y(n4113) );
  INVX1 U18987 ( .A(n4033), .Y(n4111) );
  INVX1 U18988 ( .A(n4033), .Y(n4114) );
  INVX1 U18989 ( .A(top_core_c_ready), .Y(n3686) );
  INVX1 U18990 ( .A(n3948), .Y(n3962) );
  INVX1 U18991 ( .A(n3960), .Y(n3961) );
  INVX1 U18992 ( .A(top_core_k_ready), .Y(n3706) );
  INVX1 U18993 ( .A(top_core_k_ready), .Y(n3705) );
  INVX1 U18994 ( .A(n3704), .Y(n3708) );
  INVX1 U18995 ( .A(n3704), .Y(n3707) );
  INVX1 U18996 ( .A(top_core_KE_prev_key1_reg_82_), .Y(n1679) );
  OR3XL U18997 ( .A(top_core_KE_n2509), .B(top_core_KE_n2510), .C(n2292), .Y(
        n741) );
  INVX1 U18998 ( .A(top_core_EC_ss_in[85]), .Y(n2865) );
  INVX1 U18999 ( .A(top_core_EC_ss_in[5]), .Y(n3466) );
  INVX1 U19000 ( .A(top_core_EC_ss_in[37]), .Y(n3225) );
  INVX1 U19001 ( .A(top_core_EC_ss_in[45]), .Y(n3164) );
  INVX1 U19002 ( .A(top_core_EC_ss_in[77]), .Y(n2926) );
  INVX1 U19003 ( .A(top_core_EC_ss_in[125]), .Y(n2562) );
  INVX1 U19004 ( .A(top_core_EC_ss_in[109]), .Y(n2684) );
  INVX1 U19005 ( .A(top_core_EC_ss_in[29]), .Y(n3286) );
  INVX1 U19006 ( .A(top_core_EC_ss_in[69]), .Y(n2987) );
  INVX1 U19007 ( .A(top_core_EC_ss_in[101]), .Y(n2744) );
  INVX1 U19008 ( .A(top_core_EC_ss_in[53]), .Y(n3106) );
  INVX1 U19009 ( .A(top_core_EC_ss_in[93]), .Y(n2805) );
  NOR4X2 U19010 ( .A(n4192), .B(n_ADDR[6]), .C(n_ADDR[4]), .D(n_ADDR[5]), .Y(
        top_core_io_n621) );
  NOR2BX1 U19011 ( .AN(top_core_io_n189), .B(n_ADDR[4]), .Y(top_core_io_n324)
         );
  NOR3BX1 U19012 ( .AN(n_ADDR[5]), .B(n4192), .C(n_ADDR[6]), .Y(
        top_core_io_n189) );
  AND2X2 U19013 ( .A(top_core_io_n189), .B(n_ADDR[4]), .Y(top_core_io_n154) );
  OAI22X1 U19014 ( .A0(n1557), .A1(n274), .B0(n4176), .B1(n4774), .Y(
        top_core_io_n1178) );
  OAI22X1 U19015 ( .A0(n1560), .A1(n274), .B0(n4176), .B1(n4773), .Y(
        top_core_io_n1177) );
  OAI22X1 U19016 ( .A0(n1563), .A1(n274), .B0(n4176), .B1(n4772), .Y(
        top_core_io_n1176) );
  OAI22X1 U19017 ( .A0(n1566), .A1(n274), .B0(n4176), .B1(n4771), .Y(
        top_core_io_n1175) );
  OAI22X1 U19018 ( .A0(n1569), .A1(n274), .B0(n4176), .B1(n4770), .Y(
        top_core_io_n1174) );
  OAI22X1 U19019 ( .A0(n1572), .A1(n274), .B0(n4176), .B1(n4769), .Y(
        top_core_io_n1173) );
  OAI22X1 U19020 ( .A0(n1575), .A1(n274), .B0(n4176), .B1(n4768), .Y(
        top_core_io_n1172) );
  OAI22X1 U19021 ( .A0(n1580), .A1(n274), .B0(n4176), .B1(n4767), .Y(
        top_core_io_n1171) );
  OAI22X1 U19022 ( .A0(n1557), .A1(n275), .B0(n4180), .B1(n4766), .Y(
        top_core_io_n1170) );
  OAI22X1 U19023 ( .A0(n1560), .A1(n275), .B0(n4180), .B1(n4765), .Y(
        top_core_io_n1169) );
  OAI22X1 U19024 ( .A0(n1563), .A1(n275), .B0(n4180), .B1(n4764), .Y(
        top_core_io_n1168) );
  OAI22X1 U19025 ( .A0(n1566), .A1(n275), .B0(n4180), .B1(n4763), .Y(
        top_core_io_n1167) );
  OAI22X1 U19026 ( .A0(n1569), .A1(n275), .B0(n4180), .B1(n4762), .Y(
        top_core_io_n1166) );
  OAI22X1 U19027 ( .A0(n1572), .A1(n275), .B0(n4180), .B1(n4761), .Y(
        top_core_io_n1165) );
  OAI22X1 U19028 ( .A0(n1575), .A1(n275), .B0(n4180), .B1(n4760), .Y(
        top_core_io_n1164) );
  OAI22X1 U19029 ( .A0(n1580), .A1(n275), .B0(n4180), .B1(n4759), .Y(
        top_core_io_n1163) );
  OAI22X1 U19030 ( .A0(n1557), .A1(n276), .B0(n4184), .B1(n4758), .Y(
        top_core_io_n1162) );
  OAI22X1 U19031 ( .A0(n1560), .A1(n276), .B0(n4184), .B1(n4757), .Y(
        top_core_io_n1161) );
  OAI22X1 U19032 ( .A0(n1563), .A1(n276), .B0(n4184), .B1(n4756), .Y(
        top_core_io_n1160) );
  OAI22X1 U19033 ( .A0(n1566), .A1(n276), .B0(n4184), .B1(n4755), .Y(
        top_core_io_n1159) );
  OAI22X1 U19034 ( .A0(n1569), .A1(n276), .B0(n4184), .B1(n4754), .Y(
        top_core_io_n1158) );
  OAI22X1 U19035 ( .A0(n1572), .A1(n276), .B0(n4184), .B1(n4753), .Y(
        top_core_io_n1157) );
  OAI22X1 U19036 ( .A0(n1575), .A1(n276), .B0(n4184), .B1(n4752), .Y(
        top_core_io_n1156) );
  OAI22X1 U19037 ( .A0(n1580), .A1(n276), .B0(n4184), .B1(n4751), .Y(
        top_core_io_n1155) );
  OAI22X1 U19038 ( .A0(n1557), .A1(n277), .B0(n4188), .B1(n4750), .Y(
        top_core_io_n1154) );
  OAI22X1 U19039 ( .A0(n1560), .A1(n277), .B0(n4188), .B1(n4749), .Y(
        top_core_io_n1153) );
  OAI22X1 U19040 ( .A0(n1563), .A1(n277), .B0(n4188), .B1(n4748), .Y(
        top_core_io_n1152) );
  OAI22X1 U19041 ( .A0(n1566), .A1(n277), .B0(n4188), .B1(n4747), .Y(
        top_core_io_n1151) );
  OAI22X1 U19042 ( .A0(n1569), .A1(n277), .B0(n4188), .B1(n4746), .Y(
        top_core_io_n1150) );
  OAI22X1 U19043 ( .A0(n1572), .A1(n277), .B0(n4188), .B1(n4745), .Y(
        top_core_io_n1149) );
  OAI22X1 U19044 ( .A0(n1575), .A1(n277), .B0(n4188), .B1(n4744), .Y(
        top_core_io_n1148) );
  OAI22X1 U19045 ( .A0(n1580), .A1(n277), .B0(n4188), .B1(n4743), .Y(
        top_core_io_n1147) );
  OAI22X1 U19046 ( .A0(n1557), .A1(n282), .B0(n4177), .B1(n4742), .Y(
        top_core_io_n1146) );
  OAI22X1 U19047 ( .A0(n1560), .A1(n282), .B0(n4177), .B1(n4741), .Y(
        top_core_io_n1145) );
  OAI22X1 U19048 ( .A0(n1563), .A1(n282), .B0(n4177), .B1(n4740), .Y(
        top_core_io_n1144) );
  OAI22X1 U19049 ( .A0(n1566), .A1(n282), .B0(n4177), .B1(n4739), .Y(
        top_core_io_n1143) );
  OAI22X1 U19050 ( .A0(n1569), .A1(n282), .B0(n4177), .B1(n4738), .Y(
        top_core_io_n1142) );
  OAI22X1 U19051 ( .A0(n1572), .A1(n282), .B0(n4177), .B1(n4737), .Y(
        top_core_io_n1141) );
  OAI22X1 U19052 ( .A0(n1575), .A1(n282), .B0(n4177), .B1(n4736), .Y(
        top_core_io_n1140) );
  OAI22X1 U19053 ( .A0(n1580), .A1(n282), .B0(n4177), .B1(n4735), .Y(
        top_core_io_n1139) );
  OAI22X1 U19054 ( .A0(n1557), .A1(n283), .B0(n4181), .B1(n4734), .Y(
        top_core_io_n1138) );
  OAI22X1 U19055 ( .A0(n1560), .A1(n283), .B0(n4181), .B1(n4733), .Y(
        top_core_io_n1137) );
  OAI22X1 U19056 ( .A0(n1563), .A1(n283), .B0(n4181), .B1(n4732), .Y(
        top_core_io_n1136) );
  OAI22X1 U19057 ( .A0(n1566), .A1(n283), .B0(n4181), .B1(n4731), .Y(
        top_core_io_n1135) );
  OAI22X1 U19058 ( .A0(n1569), .A1(n283), .B0(n4181), .B1(n4730), .Y(
        top_core_io_n1134) );
  OAI22X1 U19059 ( .A0(n1572), .A1(n283), .B0(n4181), .B1(n4729), .Y(
        top_core_io_n1133) );
  OAI22X1 U19060 ( .A0(n1575), .A1(n283), .B0(n4181), .B1(n4728), .Y(
        top_core_io_n1132) );
  OAI22X1 U19061 ( .A0(n1580), .A1(n283), .B0(n4181), .B1(n4727), .Y(
        top_core_io_n1131) );
  OAI22X1 U19062 ( .A0(n1557), .A1(n284), .B0(n4185), .B1(n4726), .Y(
        top_core_io_n1130) );
  OAI22X1 U19063 ( .A0(n1560), .A1(n284), .B0(n4185), .B1(n4725), .Y(
        top_core_io_n1129) );
  OAI22X1 U19064 ( .A0(n1563), .A1(n284), .B0(n4185), .B1(n4724), .Y(
        top_core_io_n1128) );
  OAI22X1 U19065 ( .A0(n1566), .A1(n284), .B0(n4185), .B1(n4723), .Y(
        top_core_io_n1127) );
  OAI22X1 U19066 ( .A0(n1569), .A1(n284), .B0(n4185), .B1(n4722), .Y(
        top_core_io_n1126) );
  OAI22X1 U19067 ( .A0(n1572), .A1(n284), .B0(n4185), .B1(n4721), .Y(
        top_core_io_n1125) );
  OAI22X1 U19068 ( .A0(n1575), .A1(n284), .B0(n4185), .B1(n4720), .Y(
        top_core_io_n1124) );
  OAI22X1 U19069 ( .A0(n1580), .A1(n284), .B0(n4185), .B1(n4719), .Y(
        top_core_io_n1123) );
  OAI22X1 U19070 ( .A0(n1557), .A1(n285), .B0(n4189), .B1(n4718), .Y(
        top_core_io_n1122) );
  OAI22X1 U19071 ( .A0(n1560), .A1(n285), .B0(n4189), .B1(n4717), .Y(
        top_core_io_n1121) );
  OAI22X1 U19072 ( .A0(n1563), .A1(n285), .B0(n4189), .B1(n4716), .Y(
        top_core_io_n1120) );
  OAI22X1 U19073 ( .A0(n1566), .A1(n285), .B0(n4189), .B1(n4715), .Y(
        top_core_io_n1119) );
  OAI22X1 U19074 ( .A0(n1569), .A1(n285), .B0(n4189), .B1(n4714), .Y(
        top_core_io_n1118) );
  OAI22X1 U19075 ( .A0(n1572), .A1(n285), .B0(n4189), .B1(n4713), .Y(
        top_core_io_n1117) );
  OAI22X1 U19076 ( .A0(n1575), .A1(n285), .B0(n4189), .B1(n4712), .Y(
        top_core_io_n1116) );
  OAI22X1 U19077 ( .A0(n1580), .A1(n285), .B0(n4189), .B1(n4711), .Y(
        top_core_io_n1115) );
  OAI22X1 U19078 ( .A0(n1557), .A1(n267), .B0(n4178), .B1(n4710), .Y(
        top_core_io_n1114) );
  OAI22X1 U19079 ( .A0(n1560), .A1(n267), .B0(n4178), .B1(n4709), .Y(
        top_core_io_n1113) );
  OAI22X1 U19080 ( .A0(n1563), .A1(n267), .B0(n4178), .B1(n4708), .Y(
        top_core_io_n1112) );
  OAI22X1 U19081 ( .A0(n1566), .A1(n267), .B0(n4178), .B1(n4707), .Y(
        top_core_io_n1111) );
  OAI22X1 U19082 ( .A0(n1569), .A1(n267), .B0(n4178), .B1(n4706), .Y(
        top_core_io_n1110) );
  OAI22X1 U19083 ( .A0(n1572), .A1(n267), .B0(n4178), .B1(n4705), .Y(
        top_core_io_n1109) );
  OAI22X1 U19084 ( .A0(n1575), .A1(n267), .B0(n4178), .B1(n4704), .Y(
        top_core_io_n1108) );
  OAI22X1 U19085 ( .A0(n1580), .A1(n267), .B0(n4178), .B1(n4703), .Y(
        top_core_io_n1107) );
  OAI22X1 U19086 ( .A0(n1557), .A1(n268), .B0(n4182), .B1(n4702), .Y(
        top_core_io_n1106) );
  OAI22X1 U19087 ( .A0(n1560), .A1(n268), .B0(n4182), .B1(n4701), .Y(
        top_core_io_n1105) );
  OAI22X1 U19088 ( .A0(n1563), .A1(n268), .B0(n4182), .B1(n4700), .Y(
        top_core_io_n1104) );
  OAI22X1 U19089 ( .A0(n1566), .A1(n268), .B0(n4182), .B1(n4699), .Y(
        top_core_io_n1103) );
  OAI22X1 U19090 ( .A0(n1569), .A1(n268), .B0(n4182), .B1(n4698), .Y(
        top_core_io_n1102) );
  OAI22X1 U19091 ( .A0(n1572), .A1(n268), .B0(n4182), .B1(n4697), .Y(
        top_core_io_n1101) );
  OAI22X1 U19092 ( .A0(n1575), .A1(n268), .B0(n4182), .B1(n4696), .Y(
        top_core_io_n1100) );
  OAI22X1 U19093 ( .A0(n1580), .A1(n268), .B0(n4182), .B1(n4695), .Y(
        top_core_io_n1099) );
  OAI22X1 U19094 ( .A0(n1557), .A1(n269), .B0(n4186), .B1(n4694), .Y(
        top_core_io_n1098) );
  OAI22X1 U19095 ( .A0(n1560), .A1(n269), .B0(n4186), .B1(n4693), .Y(
        top_core_io_n1097) );
  OAI22X1 U19096 ( .A0(n1563), .A1(n269), .B0(n4186), .B1(n4692), .Y(
        top_core_io_n1096) );
  OAI22X1 U19097 ( .A0(n1566), .A1(n269), .B0(n4186), .B1(n4691), .Y(
        top_core_io_n1095) );
  OAI22X1 U19098 ( .A0(n1569), .A1(n269), .B0(n4186), .B1(n4690), .Y(
        top_core_io_n1094) );
  OAI22X1 U19099 ( .A0(n1572), .A1(n269), .B0(n4186), .B1(n4689), .Y(
        top_core_io_n1093) );
  OAI22X1 U19100 ( .A0(n1575), .A1(n269), .B0(n4186), .B1(n4688), .Y(
        top_core_io_n1092) );
  OAI22X1 U19101 ( .A0(n1579), .A1(n269), .B0(n4186), .B1(n4687), .Y(
        top_core_io_n1091) );
  OAI22X1 U19102 ( .A0(n1557), .A1(n270), .B0(n4190), .B1(n4686), .Y(
        top_core_io_n1090) );
  OAI22X1 U19103 ( .A0(n1560), .A1(n270), .B0(n4190), .B1(n4685), .Y(
        top_core_io_n1089) );
  OAI22X1 U19104 ( .A0(n1563), .A1(n270), .B0(n4190), .B1(n4684), .Y(
        top_core_io_n1088) );
  OAI22X1 U19105 ( .A0(n1566), .A1(n270), .B0(n4190), .B1(n4683), .Y(
        top_core_io_n1087) );
  OAI22X1 U19106 ( .A0(n1569), .A1(n270), .B0(n4190), .B1(n4682), .Y(
        top_core_io_n1086) );
  OAI22X1 U19107 ( .A0(n1572), .A1(n270), .B0(n4190), .B1(n4681), .Y(
        top_core_io_n1085) );
  OAI22X1 U19108 ( .A0(n1575), .A1(n270), .B0(n4190), .B1(n4680), .Y(
        top_core_io_n1084) );
  OAI22X1 U19109 ( .A0(n1579), .A1(n270), .B0(n4190), .B1(n4679), .Y(
        top_core_io_n1083) );
  OAI22X1 U19110 ( .A0(n1558), .A1(n47), .B0(n4179), .B1(n4678), .Y(
        top_core_io_n1082) );
  OAI22X1 U19111 ( .A0(n1561), .A1(n47), .B0(n4179), .B1(n4677), .Y(
        top_core_io_n1081) );
  OAI22X1 U19112 ( .A0(n1564), .A1(n47), .B0(n4179), .B1(n4676), .Y(
        top_core_io_n1080) );
  OAI22X1 U19113 ( .A0(n1567), .A1(n47), .B0(n4179), .B1(n4675), .Y(
        top_core_io_n1079) );
  OAI22X1 U19114 ( .A0(n1570), .A1(n47), .B0(n4179), .B1(n4674), .Y(
        top_core_io_n1078) );
  OAI22X1 U19115 ( .A0(n1573), .A1(n47), .B0(n4179), .B1(n4673), .Y(
        top_core_io_n1077) );
  OAI22X1 U19116 ( .A0(n1576), .A1(n47), .B0(n4179), .B1(n4672), .Y(
        top_core_io_n1076) );
  OAI22X1 U19117 ( .A0(n1579), .A1(n47), .B0(n4179), .B1(n4671), .Y(
        top_core_io_n1075) );
  OAI22X1 U19118 ( .A0(n1558), .A1(n48), .B0(n4183), .B1(n4670), .Y(
        top_core_io_n1074) );
  OAI22X1 U19119 ( .A0(n1561), .A1(n48), .B0(n4183), .B1(n4669), .Y(
        top_core_io_n1073) );
  OAI22X1 U19120 ( .A0(n1564), .A1(n48), .B0(n4183), .B1(n4668), .Y(
        top_core_io_n1072) );
  OAI22X1 U19121 ( .A0(n1567), .A1(n48), .B0(n4183), .B1(n4667), .Y(
        top_core_io_n1071) );
  OAI22X1 U19122 ( .A0(n1570), .A1(n48), .B0(n4183), .B1(n4666), .Y(
        top_core_io_n1070) );
  OAI22X1 U19123 ( .A0(n1573), .A1(n48), .B0(n4183), .B1(n4665), .Y(
        top_core_io_n1069) );
  OAI22X1 U19124 ( .A0(n1576), .A1(n48), .B0(n4183), .B1(n4664), .Y(
        top_core_io_n1068) );
  OAI22X1 U19125 ( .A0(n1579), .A1(n48), .B0(n4183), .B1(n4663), .Y(
        top_core_io_n1067) );
  OAI22X1 U19126 ( .A0(n1558), .A1(n49), .B0(n4187), .B1(n4662), .Y(
        top_core_io_n1066) );
  OAI22X1 U19127 ( .A0(n1561), .A1(n49), .B0(n4187), .B1(n4661), .Y(
        top_core_io_n1065) );
  OAI22X1 U19128 ( .A0(n1564), .A1(n49), .B0(n4187), .B1(n4660), .Y(
        top_core_io_n1064) );
  OAI22X1 U19129 ( .A0(n1567), .A1(n49), .B0(n4187), .B1(n4659), .Y(
        top_core_io_n1063) );
  OAI22X1 U19130 ( .A0(n1570), .A1(n49), .B0(n4187), .B1(n4658), .Y(
        top_core_io_n1062) );
  OAI22X1 U19131 ( .A0(n1573), .A1(n49), .B0(n4187), .B1(n4657), .Y(
        top_core_io_n1061) );
  OAI22X1 U19132 ( .A0(n1576), .A1(n49), .B0(n4187), .B1(n4656), .Y(
        top_core_io_n1060) );
  OAI22X1 U19133 ( .A0(n1579), .A1(n49), .B0(n4187), .B1(n4655), .Y(
        top_core_io_n1059) );
  OAI22X1 U19134 ( .A0(n1558), .A1(n87), .B0(n4191), .B1(n4654), .Y(
        top_core_io_n1058) );
  OAI22X1 U19135 ( .A0(n1561), .A1(n87), .B0(n4191), .B1(n4653), .Y(
        top_core_io_n1057) );
  OAI22X1 U19136 ( .A0(n1564), .A1(n87), .B0(n4191), .B1(n4652), .Y(
        top_core_io_n1056) );
  OAI22X1 U19137 ( .A0(n1567), .A1(n87), .B0(n4191), .B1(n4651), .Y(
        top_core_io_n1055) );
  OAI22X1 U19138 ( .A0(n1570), .A1(n87), .B0(n4191), .B1(n4650), .Y(
        top_core_io_n1054) );
  OAI22X1 U19139 ( .A0(n1573), .A1(n87), .B0(n4191), .B1(n4649), .Y(
        top_core_io_n1053) );
  OAI22X1 U19140 ( .A0(n1576), .A1(n87), .B0(n4191), .B1(n4648), .Y(
        top_core_io_n1052) );
  OAI22X1 U19141 ( .A0(n1579), .A1(n87), .B0(n4191), .B1(n4647), .Y(
        top_core_io_n1051) );
  OAI22X1 U19142 ( .A0(n1558), .A1(n278), .B0(n4145), .B1(n4518), .Y(
        top_core_io_n922) );
  OAI22X1 U19143 ( .A0(n1561), .A1(n278), .B0(n4145), .B1(n4517), .Y(
        top_core_io_n921) );
  OAI22X1 U19144 ( .A0(n1564), .A1(n278), .B0(n4145), .B1(n4516), .Y(
        top_core_io_n920) );
  OAI22X1 U19145 ( .A0(n1567), .A1(n278), .B0(n4145), .B1(n4515), .Y(
        top_core_io_n919) );
  OAI22X1 U19146 ( .A0(n1570), .A1(n278), .B0(n4145), .B1(n4514), .Y(
        top_core_io_n918) );
  OAI22X1 U19147 ( .A0(n1573), .A1(n278), .B0(n4145), .B1(n4513), .Y(
        top_core_io_n917) );
  OAI22X1 U19148 ( .A0(n1576), .A1(n278), .B0(n4145), .B1(n4512), .Y(
        top_core_io_n916) );
  OAI22X1 U19149 ( .A0(n1579), .A1(n278), .B0(n4145), .B1(n4511), .Y(
        top_core_io_n915) );
  OAI22X1 U19150 ( .A0(n1558), .A1(n279), .B0(n4149), .B1(n4510), .Y(
        top_core_io_n914) );
  OAI22X1 U19151 ( .A0(n1561), .A1(n279), .B0(n4149), .B1(n4509), .Y(
        top_core_io_n913) );
  OAI22X1 U19152 ( .A0(n1564), .A1(n279), .B0(n4149), .B1(n4508), .Y(
        top_core_io_n912) );
  OAI22X1 U19153 ( .A0(n1567), .A1(n279), .B0(n4149), .B1(n4507), .Y(
        top_core_io_n911) );
  OAI22X1 U19154 ( .A0(n1570), .A1(n279), .B0(n4149), .B1(n4506), .Y(
        top_core_io_n910) );
  OAI22X1 U19155 ( .A0(n1573), .A1(n279), .B0(n4149), .B1(n4505), .Y(
        top_core_io_n909) );
  OAI22X1 U19156 ( .A0(n1576), .A1(n279), .B0(n4149), .B1(n4504), .Y(
        top_core_io_n908) );
  OAI22X1 U19157 ( .A0(n1579), .A1(n279), .B0(n4149), .B1(n4503), .Y(
        top_core_io_n907) );
  OAI22X1 U19158 ( .A0(n1558), .A1(n280), .B0(n4153), .B1(n4502), .Y(
        top_core_io_n906) );
  OAI22X1 U19159 ( .A0(n1561), .A1(n280), .B0(n4153), .B1(n4501), .Y(
        top_core_io_n905) );
  OAI22X1 U19160 ( .A0(n1564), .A1(n280), .B0(n4153), .B1(n4500), .Y(
        top_core_io_n904) );
  OAI22X1 U19161 ( .A0(n1567), .A1(n280), .B0(n4153), .B1(n4499), .Y(
        top_core_io_n903) );
  OAI22X1 U19162 ( .A0(n1570), .A1(n280), .B0(n4153), .B1(n4498), .Y(
        top_core_io_n902) );
  OAI22X1 U19163 ( .A0(n1573), .A1(n280), .B0(n4153), .B1(n4497), .Y(
        top_core_io_n901) );
  OAI22X1 U19164 ( .A0(n1576), .A1(n280), .B0(n4153), .B1(n4496), .Y(
        top_core_io_n900) );
  OAI22X1 U19165 ( .A0(n1579), .A1(n280), .B0(n4153), .B1(n4495), .Y(
        top_core_io_n899) );
  OAI22X1 U19166 ( .A0(n1558), .A1(n281), .B0(n4157), .B1(n4494), .Y(
        top_core_io_n898) );
  OAI22X1 U19167 ( .A0(n1561), .A1(n281), .B0(n4157), .B1(n4493), .Y(
        top_core_io_n897) );
  OAI22X1 U19168 ( .A0(n1564), .A1(n281), .B0(n4157), .B1(n4492), .Y(
        top_core_io_n896) );
  OAI22X1 U19169 ( .A0(n1567), .A1(n281), .B0(n4157), .B1(n4491), .Y(
        top_core_io_n895) );
  OAI22X1 U19170 ( .A0(n1570), .A1(n281), .B0(n4157), .B1(n4490), .Y(
        top_core_io_n894) );
  OAI22X1 U19171 ( .A0(n1573), .A1(n281), .B0(n4157), .B1(n4489), .Y(
        top_core_io_n893) );
  OAI22X1 U19172 ( .A0(n1576), .A1(n281), .B0(n4157), .B1(n4488), .Y(
        top_core_io_n892) );
  OAI22X1 U19173 ( .A0(n1579), .A1(n281), .B0(n4157), .B1(n4487), .Y(
        top_core_io_n891) );
  OAI22X1 U19174 ( .A0(n1558), .A1(n286), .B0(n4146), .B1(n4486), .Y(
        top_core_io_n890) );
  OAI22X1 U19175 ( .A0(n1561), .A1(n286), .B0(n4146), .B1(n4485), .Y(
        top_core_io_n889) );
  OAI22X1 U19176 ( .A0(n1564), .A1(n286), .B0(n4146), .B1(n4484), .Y(
        top_core_io_n888) );
  OAI22X1 U19177 ( .A0(n1567), .A1(n286), .B0(n4146), .B1(n4483), .Y(
        top_core_io_n887) );
  OAI22X1 U19178 ( .A0(n1570), .A1(n286), .B0(n4146), .B1(n4482), .Y(
        top_core_io_n886) );
  OAI22X1 U19179 ( .A0(n1573), .A1(n286), .B0(n4146), .B1(n4481), .Y(
        top_core_io_n885) );
  OAI22X1 U19180 ( .A0(n1576), .A1(n286), .B0(n4146), .B1(n4480), .Y(
        top_core_io_n884) );
  OAI22X1 U19181 ( .A0(n1579), .A1(n286), .B0(n4146), .B1(n4479), .Y(
        top_core_io_n883) );
  OAI22X1 U19182 ( .A0(n1558), .A1(n287), .B0(n4150), .B1(n4478), .Y(
        top_core_io_n882) );
  OAI22X1 U19183 ( .A0(n1561), .A1(n287), .B0(n4150), .B1(n4477), .Y(
        top_core_io_n881) );
  OAI22X1 U19184 ( .A0(n1564), .A1(n287), .B0(n4150), .B1(n4476), .Y(
        top_core_io_n880) );
  OAI22X1 U19185 ( .A0(n1567), .A1(n287), .B0(n4150), .B1(n4475), .Y(
        top_core_io_n879) );
  OAI22X1 U19186 ( .A0(n1570), .A1(n287), .B0(n4150), .B1(n4474), .Y(
        top_core_io_n878) );
  OAI22X1 U19187 ( .A0(n1573), .A1(n287), .B0(n4150), .B1(n4473), .Y(
        top_core_io_n877) );
  OAI22X1 U19188 ( .A0(n1576), .A1(n287), .B0(n4150), .B1(n4472), .Y(
        top_core_io_n876) );
  OAI22X1 U19189 ( .A0(n1579), .A1(n287), .B0(n4150), .B1(n4471), .Y(
        top_core_io_n875) );
  OAI22X1 U19190 ( .A0(n1558), .A1(n288), .B0(n4154), .B1(n4470), .Y(
        top_core_io_n874) );
  OAI22X1 U19191 ( .A0(n1561), .A1(n288), .B0(n4154), .B1(n4469), .Y(
        top_core_io_n873) );
  OAI22X1 U19192 ( .A0(n1564), .A1(n288), .B0(n4154), .B1(n4468), .Y(
        top_core_io_n872) );
  OAI22X1 U19193 ( .A0(n1567), .A1(n288), .B0(n4154), .B1(n4467), .Y(
        top_core_io_n871) );
  OAI22X1 U19194 ( .A0(n1570), .A1(n288), .B0(n4154), .B1(n4466), .Y(
        top_core_io_n870) );
  OAI22X1 U19195 ( .A0(n1573), .A1(n288), .B0(n4154), .B1(n4465), .Y(
        top_core_io_n869) );
  OAI22X1 U19196 ( .A0(n1576), .A1(n288), .B0(n4154), .B1(n4464), .Y(
        top_core_io_n868) );
  OAI22X1 U19197 ( .A0(n1579), .A1(n288), .B0(n4154), .B1(n4463), .Y(
        top_core_io_n867) );
  OAI22X1 U19198 ( .A0(n1558), .A1(n289), .B0(n4158), .B1(n4462), .Y(
        top_core_io_n866) );
  OAI22X1 U19199 ( .A0(n1561), .A1(n289), .B0(n4158), .B1(n4461), .Y(
        top_core_io_n865) );
  OAI22X1 U19200 ( .A0(n1564), .A1(n289), .B0(n4158), .B1(n4460), .Y(
        top_core_io_n864) );
  OAI22X1 U19201 ( .A0(n1567), .A1(n289), .B0(n4158), .B1(n4459), .Y(
        top_core_io_n863) );
  OAI22X1 U19202 ( .A0(n1570), .A1(n289), .B0(n4158), .B1(n4458), .Y(
        top_core_io_n862) );
  OAI22X1 U19203 ( .A0(n1573), .A1(n289), .B0(n4158), .B1(n4457), .Y(
        top_core_io_n861) );
  OAI22X1 U19204 ( .A0(n1576), .A1(n289), .B0(n4158), .B1(n4456), .Y(
        top_core_io_n860) );
  OAI22X1 U19205 ( .A0(n1580), .A1(n289), .B0(n4158), .B1(n4455), .Y(
        top_core_io_n859) );
  OAI22X1 U19206 ( .A0(n1559), .A1(n271), .B0(n4147), .B1(n4454), .Y(
        top_core_io_n858) );
  OAI22X1 U19207 ( .A0(n1562), .A1(n271), .B0(n4147), .B1(n4453), .Y(
        top_core_io_n857) );
  OAI22X1 U19208 ( .A0(n1565), .A1(n271), .B0(n4147), .B1(n4452), .Y(
        top_core_io_n856) );
  OAI22X1 U19209 ( .A0(n1568), .A1(n271), .B0(n4147), .B1(n4451), .Y(
        top_core_io_n855) );
  OAI22X1 U19210 ( .A0(n1571), .A1(n271), .B0(n4147), .B1(n4450), .Y(
        top_core_io_n854) );
  OAI22X1 U19211 ( .A0(n1572), .A1(n271), .B0(n4147), .B1(n4449), .Y(
        top_core_io_n853) );
  OAI22X1 U19212 ( .A0(n1575), .A1(n271), .B0(n4147), .B1(n4448), .Y(
        top_core_io_n852) );
  OAI22X1 U19213 ( .A0(n1579), .A1(n271), .B0(n4147), .B1(n4447), .Y(
        top_core_io_n851) );
  OAI22X1 U19214 ( .A0(n1559), .A1(n84), .B0(n4151), .B1(n4446), .Y(
        top_core_io_n850) );
  OAI22X1 U19215 ( .A0(n1562), .A1(n84), .B0(n4151), .B1(n4445), .Y(
        top_core_io_n849) );
  OAI22X1 U19216 ( .A0(n1565), .A1(n84), .B0(n4151), .B1(n4444), .Y(
        top_core_io_n848) );
  OAI22X1 U19217 ( .A0(n1568), .A1(n84), .B0(n4151), .B1(n4443), .Y(
        top_core_io_n847) );
  OAI22X1 U19218 ( .A0(n1571), .A1(n84), .B0(n4151), .B1(n4442), .Y(
        top_core_io_n846) );
  OAI22X1 U19219 ( .A0(n1573), .A1(n84), .B0(n4151), .B1(n4441), .Y(
        top_core_io_n845) );
  OAI22X1 U19220 ( .A0(n1576), .A1(n84), .B0(n4151), .B1(n4440), .Y(
        top_core_io_n844) );
  OAI22X1 U19221 ( .A0(n1578), .A1(n84), .B0(n4151), .B1(n4439), .Y(
        top_core_io_n843) );
  OAI22X1 U19222 ( .A0(n1559), .A1(n272), .B0(n4155), .B1(n4438), .Y(
        top_core_io_n842) );
  OAI22X1 U19223 ( .A0(n1562), .A1(n272), .B0(n4155), .B1(n4437), .Y(
        top_core_io_n841) );
  OAI22X1 U19224 ( .A0(n1565), .A1(n272), .B0(n4155), .B1(n4436), .Y(
        top_core_io_n840) );
  OAI22X1 U19225 ( .A0(n1568), .A1(n272), .B0(n4155), .B1(n4435), .Y(
        top_core_io_n839) );
  OAI22X1 U19226 ( .A0(n1571), .A1(n272), .B0(n4155), .B1(n4434), .Y(
        top_core_io_n838) );
  OAI22X1 U19227 ( .A0(n1573), .A1(n272), .B0(n4155), .B1(n4433), .Y(
        top_core_io_n837) );
  OAI22X1 U19228 ( .A0(n1576), .A1(n272), .B0(n4155), .B1(n4432), .Y(
        top_core_io_n836) );
  OAI22X1 U19229 ( .A0(n1578), .A1(n272), .B0(n4155), .B1(n4431), .Y(
        top_core_io_n835) );
  OAI22X1 U19230 ( .A0(n1559), .A1(n273), .B0(n4159), .B1(n4430), .Y(
        top_core_io_n834) );
  OAI22X1 U19231 ( .A0(n1562), .A1(n273), .B0(n4159), .B1(n4429), .Y(
        top_core_io_n833) );
  OAI22X1 U19232 ( .A0(n1565), .A1(n273), .B0(n4159), .B1(n4428), .Y(
        top_core_io_n832) );
  OAI22X1 U19233 ( .A0(n1568), .A1(n273), .B0(n4159), .B1(n4427), .Y(
        top_core_io_n831) );
  OAI22X1 U19234 ( .A0(n1571), .A1(n273), .B0(n4159), .B1(n4426), .Y(
        top_core_io_n830) );
  OAI22X1 U19235 ( .A0(n1573), .A1(n273), .B0(n4159), .B1(n4425), .Y(
        top_core_io_n829) );
  OAI22X1 U19236 ( .A0(n1576), .A1(n273), .B0(n4159), .B1(n4424), .Y(
        top_core_io_n828) );
  OAI22X1 U19237 ( .A0(n1578), .A1(n273), .B0(n4159), .B1(n4423), .Y(
        top_core_io_n827) );
  OAI22X1 U19238 ( .A0(n1559), .A1(n7), .B0(n4148), .B1(n4422), .Y(
        top_core_io_n826) );
  OAI22X1 U19239 ( .A0(n1562), .A1(n7), .B0(n4148), .B1(n4421), .Y(
        top_core_io_n825) );
  OAI22X1 U19240 ( .A0(n1565), .A1(n7), .B0(n4148), .B1(n4420), .Y(
        top_core_io_n824) );
  OAI22X1 U19241 ( .A0(n1568), .A1(n7), .B0(n4148), .B1(n4419), .Y(
        top_core_io_n823) );
  OAI22X1 U19242 ( .A0(n1571), .A1(n7), .B0(n4148), .B1(n4418), .Y(
        top_core_io_n822) );
  OAI22X1 U19243 ( .A0(n1573), .A1(n7), .B0(n4148), .B1(n4417), .Y(
        top_core_io_n821) );
  OAI22X1 U19244 ( .A0(n1576), .A1(n7), .B0(n4148), .B1(n4416), .Y(
        top_core_io_n820) );
  OAI22X1 U19245 ( .A0(n1578), .A1(n7), .B0(n4148), .B1(n4415), .Y(
        top_core_io_n819) );
  OAI22X1 U19246 ( .A0(n1559), .A1(n9), .B0(n4152), .B1(n4414), .Y(
        top_core_io_n818) );
  OAI22X1 U19247 ( .A0(n1562), .A1(n9), .B0(n4152), .B1(n4413), .Y(
        top_core_io_n817) );
  OAI22X1 U19248 ( .A0(n1565), .A1(n9), .B0(n4152), .B1(n4412), .Y(
        top_core_io_n816) );
  OAI22X1 U19249 ( .A0(n1568), .A1(n9), .B0(n4152), .B1(n4411), .Y(
        top_core_io_n815) );
  OAI22X1 U19250 ( .A0(n1571), .A1(n9), .B0(n4152), .B1(n4410), .Y(
        top_core_io_n814) );
  OAI22X1 U19251 ( .A0(n1573), .A1(n9), .B0(n4152), .B1(n4409), .Y(
        top_core_io_n813) );
  OAI22X1 U19252 ( .A0(n1576), .A1(n9), .B0(n4152), .B1(n4408), .Y(
        top_core_io_n812) );
  OAI22X1 U19253 ( .A0(n1580), .A1(n9), .B0(n4152), .B1(n4407), .Y(
        top_core_io_n811) );
  OAI22X1 U19254 ( .A0(n1559), .A1(n10), .B0(n4156), .B1(n4406), .Y(
        top_core_io_n810) );
  OAI22X1 U19255 ( .A0(n1562), .A1(n10), .B0(n4156), .B1(n4405), .Y(
        top_core_io_n809) );
  OAI22X1 U19256 ( .A0(n1565), .A1(n10), .B0(n4156), .B1(n4404), .Y(
        top_core_io_n808) );
  OAI22X1 U19257 ( .A0(n1568), .A1(n10), .B0(n4156), .B1(n4403), .Y(
        top_core_io_n807) );
  OAI22X1 U19258 ( .A0(n1571), .A1(n10), .B0(n4156), .B1(n4402), .Y(
        top_core_io_n806) );
  OAI22X1 U19259 ( .A0(n1574), .A1(n10), .B0(n4156), .B1(n4401), .Y(
        top_core_io_n805) );
  OAI22X1 U19260 ( .A0(n1577), .A1(n10), .B0(n4156), .B1(n4400), .Y(
        top_core_io_n804) );
  OAI22X1 U19261 ( .A0(n1580), .A1(n10), .B0(n4156), .B1(n4399), .Y(
        top_core_io_n803) );
  OAI22X1 U19262 ( .A0(n1559), .A1(n11), .B0(n4160), .B1(n4398), .Y(
        top_core_io_n802) );
  OAI22X1 U19263 ( .A0(n1562), .A1(n11), .B0(n4160), .B1(n4397), .Y(
        top_core_io_n801) );
  OAI22X1 U19264 ( .A0(n1565), .A1(n11), .B0(n4160), .B1(n4396), .Y(
        top_core_io_n800) );
  OAI22X1 U19265 ( .A0(n1568), .A1(n11), .B0(n4160), .B1(n4395), .Y(
        top_core_io_n799) );
  OAI22X1 U19266 ( .A0(n1571), .A1(n11), .B0(n4160), .B1(n4394), .Y(
        top_core_io_n798) );
  OAI22X1 U19267 ( .A0(n1574), .A1(n11), .B0(n4160), .B1(n4393), .Y(
        top_core_io_n797) );
  OAI22X1 U19268 ( .A0(n1577), .A1(n11), .B0(n4160), .B1(n4392), .Y(
        top_core_io_n796) );
  OAI22X1 U19269 ( .A0(n1580), .A1(n11), .B0(n4160), .B1(n4391), .Y(
        top_core_io_n795) );
  OAI22X1 U19270 ( .A0(n1559), .A1(n294), .B0(n4161), .B1(n4390), .Y(
        top_core_io_n794) );
  OAI22X1 U19271 ( .A0(n1562), .A1(n294), .B0(n4161), .B1(n4389), .Y(
        top_core_io_n793) );
  OAI22X1 U19272 ( .A0(n1565), .A1(n294), .B0(n4161), .B1(n4388), .Y(
        top_core_io_n792) );
  OAI22X1 U19273 ( .A0(n1568), .A1(n294), .B0(n4161), .B1(n4387), .Y(
        top_core_io_n791) );
  OAI22X1 U19274 ( .A0(n1571), .A1(n294), .B0(n4161), .B1(n4386), .Y(
        top_core_io_n790) );
  OAI22X1 U19275 ( .A0(n1574), .A1(n294), .B0(n4161), .B1(n4385), .Y(
        top_core_io_n789) );
  OAI22X1 U19276 ( .A0(n1577), .A1(n294), .B0(n4161), .B1(n4384), .Y(
        top_core_io_n788) );
  OAI22X1 U19277 ( .A0(n1579), .A1(n294), .B0(n4161), .B1(n4383), .Y(
        top_core_io_n787) );
  OAI22X1 U19278 ( .A0(n1559), .A1(n295), .B0(n4165), .B1(n4382), .Y(
        top_core_io_n786) );
  OAI22X1 U19279 ( .A0(n1562), .A1(n295), .B0(n4165), .B1(n4381), .Y(
        top_core_io_n785) );
  OAI22X1 U19280 ( .A0(n1565), .A1(n295), .B0(n4165), .B1(n4380), .Y(
        top_core_io_n784) );
  OAI22X1 U19281 ( .A0(n1568), .A1(n295), .B0(n4165), .B1(n4379), .Y(
        top_core_io_n783) );
  OAI22X1 U19282 ( .A0(n1571), .A1(n295), .B0(n4165), .B1(n4378), .Y(
        top_core_io_n782) );
  OAI22X1 U19283 ( .A0(n1572), .A1(n295), .B0(n4165), .B1(n4377), .Y(
        top_core_io_n781) );
  OAI22X1 U19284 ( .A0(n1575), .A1(n295), .B0(n4165), .B1(n4376), .Y(
        top_core_io_n780) );
  OAI22X1 U19285 ( .A0(n1580), .A1(n295), .B0(n4165), .B1(n4375), .Y(
        top_core_io_n779) );
  OAI22X1 U19286 ( .A0(n1559), .A1(n296), .B0(n4168), .B1(n4374), .Y(
        top_core_io_n778) );
  OAI22X1 U19287 ( .A0(n1562), .A1(n296), .B0(n4168), .B1(n4373), .Y(
        top_core_io_n777) );
  OAI22X1 U19288 ( .A0(n1565), .A1(n296), .B0(n4168), .B1(n4372), .Y(
        top_core_io_n776) );
  OAI22X1 U19289 ( .A0(n1568), .A1(n296), .B0(n4168), .B1(n4371), .Y(
        top_core_io_n775) );
  OAI22X1 U19290 ( .A0(n1571), .A1(n296), .B0(n4168), .B1(n4370), .Y(
        top_core_io_n774) );
  OAI22X1 U19291 ( .A0(n1572), .A1(n296), .B0(n4168), .B1(n4369), .Y(
        top_core_io_n773) );
  OAI22X1 U19292 ( .A0(n1575), .A1(n296), .B0(n4168), .B1(n4368), .Y(
        top_core_io_n772) );
  OAI22X1 U19293 ( .A0(n1579), .A1(n296), .B0(n4168), .B1(n4367), .Y(
        top_core_io_n771) );
  OAI22X1 U19294 ( .A0(n1559), .A1(n297), .B0(n4172), .B1(n4366), .Y(
        top_core_io_n770) );
  OAI22X1 U19295 ( .A0(n1562), .A1(n297), .B0(n4172), .B1(n4365), .Y(
        top_core_io_n769) );
  OAI22X1 U19296 ( .A0(n1565), .A1(n297), .B0(n4172), .B1(n4364), .Y(
        top_core_io_n768) );
  OAI22X1 U19297 ( .A0(n1568), .A1(n297), .B0(n4172), .B1(n4363), .Y(
        top_core_io_n767) );
  OAI22X1 U19298 ( .A0(n1571), .A1(n297), .B0(n4172), .B1(n4362), .Y(
        top_core_io_n766) );
  OAI22X1 U19299 ( .A0(n1574), .A1(n297), .B0(n4172), .B1(n4361), .Y(
        top_core_io_n765) );
  OAI22X1 U19300 ( .A0(n1577), .A1(n297), .B0(n4172), .B1(n4360), .Y(
        top_core_io_n764) );
  OAI22X1 U19301 ( .A0(n1580), .A1(n297), .B0(n4172), .B1(n4359), .Y(
        top_core_io_n763) );
  OAI22X1 U19302 ( .A0(n1558), .A1(n298), .B0(n4162), .B1(n4358), .Y(
        top_core_io_n762) );
  OAI22X1 U19303 ( .A0(n1561), .A1(n298), .B0(n4162), .B1(n4357), .Y(
        top_core_io_n761) );
  OAI22X1 U19304 ( .A0(n1564), .A1(n298), .B0(n4162), .B1(n4356), .Y(
        top_core_io_n760) );
  OAI22X1 U19305 ( .A0(n1567), .A1(n298), .B0(n4162), .B1(n4355), .Y(
        top_core_io_n759) );
  OAI22X1 U19306 ( .A0(n1570), .A1(n298), .B0(n4162), .B1(n4354), .Y(
        top_core_io_n758) );
  OAI22X1 U19307 ( .A0(n1574), .A1(n298), .B0(n4162), .B1(n4353), .Y(
        top_core_io_n757) );
  OAI22X1 U19308 ( .A0(n1577), .A1(n298), .B0(n4162), .B1(n4352), .Y(
        top_core_io_n756) );
  OAI22X1 U19309 ( .A0(n1578), .A1(n298), .B0(n4162), .B1(n4351), .Y(
        top_core_io_n755) );
  OAI22X1 U19310 ( .A0(n1558), .A1(n299), .B0(n4166), .B1(n4350), .Y(
        top_core_io_n754) );
  OAI22X1 U19311 ( .A0(n1561), .A1(n299), .B0(n4166), .B1(n4349), .Y(
        top_core_io_n753) );
  OAI22X1 U19312 ( .A0(n1564), .A1(n299), .B0(n4166), .B1(n4348), .Y(
        top_core_io_n752) );
  OAI22X1 U19313 ( .A0(n1567), .A1(n299), .B0(n4166), .B1(n4347), .Y(
        top_core_io_n751) );
  OAI22X1 U19314 ( .A0(n1570), .A1(n299), .B0(n4166), .B1(n4346), .Y(
        top_core_io_n750) );
  OAI22X1 U19315 ( .A0(n1574), .A1(n299), .B0(n4166), .B1(n4345), .Y(
        top_core_io_n749) );
  OAI22X1 U19316 ( .A0(n1577), .A1(n299), .B0(n4166), .B1(n4344), .Y(
        top_core_io_n748) );
  OAI22X1 U19317 ( .A0(n1578), .A1(n299), .B0(n4166), .B1(n4343), .Y(
        top_core_io_n747) );
  OAI22X1 U19318 ( .A0(n1558), .A1(n300), .B0(n4169), .B1(n4342), .Y(
        top_core_io_n746) );
  OAI22X1 U19319 ( .A0(n1561), .A1(n300), .B0(n4169), .B1(n4341), .Y(
        top_core_io_n745) );
  OAI22X1 U19320 ( .A0(n1564), .A1(n300), .B0(n4169), .B1(n4340), .Y(
        top_core_io_n744) );
  OAI22X1 U19321 ( .A0(n1567), .A1(n300), .B0(n4169), .B1(n4339), .Y(
        top_core_io_n743) );
  OAI22X1 U19322 ( .A0(n1570), .A1(n300), .B0(n4169), .B1(n4338), .Y(
        top_core_io_n742) );
  OAI22X1 U19323 ( .A0(n1574), .A1(n300), .B0(n4169), .B1(n4337), .Y(
        top_core_io_n741) );
  OAI22X1 U19324 ( .A0(n1577), .A1(n300), .B0(n4169), .B1(n4336), .Y(
        top_core_io_n740) );
  OAI22X1 U19325 ( .A0(n1578), .A1(n300), .B0(n4169), .B1(n4335), .Y(
        top_core_io_n739) );
  OAI22X1 U19326 ( .A0(n1557), .A1(n301), .B0(n4173), .B1(n4334), .Y(
        top_core_io_n738) );
  OAI22X1 U19327 ( .A0(n1560), .A1(n301), .B0(n4173), .B1(n4333), .Y(
        top_core_io_n737) );
  OAI22X1 U19328 ( .A0(n1563), .A1(n301), .B0(n4173), .B1(n4332), .Y(
        top_core_io_n736) );
  OAI22X1 U19329 ( .A0(n1566), .A1(n301), .B0(n4173), .B1(n4331), .Y(
        top_core_io_n735) );
  OAI22X1 U19330 ( .A0(n1569), .A1(n301), .B0(n4173), .B1(n4330), .Y(
        top_core_io_n734) );
  OAI22X1 U19331 ( .A0(n1574), .A1(n301), .B0(n4173), .B1(n4329), .Y(
        top_core_io_n733) );
  OAI22X1 U19332 ( .A0(n1577), .A1(n301), .B0(n4173), .B1(n4328), .Y(
        top_core_io_n732) );
  OAI22X1 U19333 ( .A0(n1578), .A1(n301), .B0(n4173), .B1(n4327), .Y(
        top_core_io_n731) );
  OAI22X1 U19334 ( .A0(n1558), .A1(n290), .B0(n4163), .B1(n4326), .Y(
        top_core_io_n730) );
  OAI22X1 U19335 ( .A0(n1561), .A1(n290), .B0(n4163), .B1(n4325), .Y(
        top_core_io_n729) );
  OAI22X1 U19336 ( .A0(n1564), .A1(n290), .B0(n4163), .B1(n4324), .Y(
        top_core_io_n728) );
  OAI22X1 U19337 ( .A0(n1567), .A1(n290), .B0(n4163), .B1(n4323), .Y(
        top_core_io_n727) );
  OAI22X1 U19338 ( .A0(n1570), .A1(n290), .B0(n4163), .B1(n4322), .Y(
        top_core_io_n726) );
  OAI22X1 U19339 ( .A0(n1574), .A1(n290), .B0(n4163), .B1(n4321), .Y(
        top_core_io_n725) );
  OAI22X1 U19340 ( .A0(n1577), .A1(n290), .B0(n4163), .B1(n4320), .Y(
        top_core_io_n724) );
  OAI22X1 U19341 ( .A0(n1578), .A1(n290), .B0(n4163), .B1(n4319), .Y(
        top_core_io_n723) );
  OAI22X1 U19342 ( .A0(n1559), .A1(n291), .B0(n4167), .B1(n4318), .Y(
        top_core_io_n722) );
  OAI22X1 U19343 ( .A0(n1562), .A1(n291), .B0(n4167), .B1(n4317), .Y(
        top_core_io_n721) );
  OAI22X1 U19344 ( .A0(n1565), .A1(n291), .B0(n4167), .B1(n4316), .Y(
        top_core_io_n720) );
  OAI22X1 U19345 ( .A0(n1568), .A1(n291), .B0(n4167), .B1(n4315), .Y(
        top_core_io_n719) );
  OAI22X1 U19346 ( .A0(n1571), .A1(n291), .B0(n4167), .B1(n4314), .Y(
        top_core_io_n718) );
  OAI22X1 U19347 ( .A0(n1574), .A1(n291), .B0(n4167), .B1(n4313), .Y(
        top_core_io_n717) );
  OAI22X1 U19348 ( .A0(n1577), .A1(n291), .B0(n4167), .B1(n4312), .Y(
        top_core_io_n716) );
  OAI22X1 U19349 ( .A0(n1578), .A1(n291), .B0(n4167), .B1(n4311), .Y(
        top_core_io_n715) );
  OAI22X1 U19350 ( .A0(n1559), .A1(n292), .B0(n4170), .B1(n4310), .Y(
        top_core_io_n714) );
  OAI22X1 U19351 ( .A0(n1562), .A1(n292), .B0(n4170), .B1(n4309), .Y(
        top_core_io_n713) );
  OAI22X1 U19352 ( .A0(n1565), .A1(n292), .B0(n4170), .B1(n4308), .Y(
        top_core_io_n712) );
  OAI22X1 U19353 ( .A0(n1568), .A1(n292), .B0(n4170), .B1(n4307), .Y(
        top_core_io_n711) );
  OAI22X1 U19354 ( .A0(n1571), .A1(n292), .B0(n4170), .B1(n4306), .Y(
        top_core_io_n710) );
  OAI22X1 U19355 ( .A0(n1574), .A1(n292), .B0(n4170), .B1(n4305), .Y(
        top_core_io_n709) );
  OAI22X1 U19356 ( .A0(n1577), .A1(n292), .B0(n4170), .B1(n4304), .Y(
        top_core_io_n708) );
  OAI22X1 U19357 ( .A0(n1578), .A1(n292), .B0(n4170), .B1(n4303), .Y(
        top_core_io_n707) );
  OAI22X1 U19358 ( .A0(n1559), .A1(n293), .B0(n4174), .B1(n4302), .Y(
        top_core_io_n706) );
  OAI22X1 U19359 ( .A0(n1562), .A1(n293), .B0(n4174), .B1(n4301), .Y(
        top_core_io_n705) );
  OAI22X1 U19360 ( .A0(n1565), .A1(n293), .B0(n4174), .B1(n4300), .Y(
        top_core_io_n704) );
  OAI22X1 U19361 ( .A0(n1568), .A1(n293), .B0(n4174), .B1(n4299), .Y(
        top_core_io_n703) );
  OAI22X1 U19362 ( .A0(n1571), .A1(n293), .B0(n4174), .B1(n4298), .Y(
        top_core_io_n702) );
  OAI22X1 U19363 ( .A0(n1574), .A1(n293), .B0(n4174), .B1(n4297), .Y(
        top_core_io_n701) );
  OAI22X1 U19364 ( .A0(n1577), .A1(n293), .B0(n4174), .B1(n4296), .Y(
        top_core_io_n700) );
  OAI22X1 U19365 ( .A0(n1578), .A1(n293), .B0(n4174), .B1(n4295), .Y(
        top_core_io_n699) );
  OAI22X1 U19366 ( .A0(n1559), .A1(n8), .B0(n4164), .B1(n4294), .Y(
        top_core_io_n698) );
  OAI22X1 U19367 ( .A0(n1562), .A1(n8), .B0(n4164), .B1(n4293), .Y(
        top_core_io_n697) );
  OAI22X1 U19368 ( .A0(n1565), .A1(n8), .B0(n4164), .B1(n4292), .Y(
        top_core_io_n696) );
  OAI22X1 U19369 ( .A0(n1568), .A1(n8), .B0(n4164), .B1(n4291), .Y(
        top_core_io_n695) );
  OAI22X1 U19370 ( .A0(n1571), .A1(n8), .B0(n4164), .B1(n4290), .Y(
        top_core_io_n694) );
  OAI22X1 U19371 ( .A0(n1574), .A1(n8), .B0(n4164), .B1(n4289), .Y(
        top_core_io_n693) );
  OAI22X1 U19372 ( .A0(n1577), .A1(n8), .B0(n4164), .B1(n4288), .Y(
        top_core_io_n692) );
  OAI22X1 U19373 ( .A0(n1578), .A1(n8), .B0(n4164), .B1(n4287), .Y(
        top_core_io_n691) );
  OAI22X1 U19374 ( .A0(n1557), .A1(n266), .B0(n13), .B1(n4286), .Y(
        top_core_io_n690) );
  OAI22X1 U19375 ( .A0(n1560), .A1(n266), .B0(n13), .B1(n4285), .Y(
        top_core_io_n689) );
  OAI22X1 U19376 ( .A0(n1563), .A1(n266), .B0(n13), .B1(n4284), .Y(
        top_core_io_n688) );
  OAI22X1 U19377 ( .A0(n1566), .A1(n266), .B0(n13), .B1(n4283), .Y(
        top_core_io_n687) );
  OAI22X1 U19378 ( .A0(n1569), .A1(n266), .B0(n13), .B1(n4282), .Y(
        top_core_io_n686) );
  OAI22X1 U19379 ( .A0(n1574), .A1(n266), .B0(n13), .B1(n4281), .Y(
        top_core_io_n685) );
  OAI22X1 U19380 ( .A0(n1577), .A1(n266), .B0(n13), .B1(n4280), .Y(
        top_core_io_n684) );
  OAI22X1 U19381 ( .A0(n1578), .A1(n266), .B0(n13), .B1(n4279), .Y(
        top_core_io_n683) );
  OAI22X1 U19382 ( .A0(n1559), .A1(n12), .B0(n4171), .B1(n4278), .Y(
        top_core_io_n682) );
  OAI22X1 U19383 ( .A0(n1562), .A1(n12), .B0(n4171), .B1(n4277), .Y(
        top_core_io_n681) );
  OAI22X1 U19384 ( .A0(n1565), .A1(n12), .B0(n4171), .B1(n4276), .Y(
        top_core_io_n680) );
  OAI22X1 U19385 ( .A0(n1568), .A1(n12), .B0(n4171), .B1(n4275), .Y(
        top_core_io_n679) );
  OAI22X1 U19386 ( .A0(n1571), .A1(n12), .B0(n4171), .B1(n4274), .Y(
        top_core_io_n678) );
  OAI22X1 U19387 ( .A0(n1574), .A1(n12), .B0(n4171), .B1(n4273), .Y(
        top_core_io_n677) );
  OAI22X1 U19388 ( .A0(n1577), .A1(n12), .B0(n4171), .B1(n4272), .Y(
        top_core_io_n676) );
  OAI22X1 U19389 ( .A0(n1578), .A1(n12), .B0(n4171), .B1(n4271), .Y(
        top_core_io_n675) );
  OAI22X1 U19390 ( .A0(n88), .A1(n1557), .B0(n4175), .B1(n4270), .Y(
        top_core_io_n674) );
  OAI22X1 U19391 ( .A0(n88), .A1(n1560), .B0(n4175), .B1(n4269), .Y(
        top_core_io_n673) );
  OAI22X1 U19392 ( .A0(n88), .A1(n1563), .B0(n4175), .B1(n4268), .Y(
        top_core_io_n672) );
  OAI22X1 U19393 ( .A0(n88), .A1(n1566), .B0(n4175), .B1(n4267), .Y(
        top_core_io_n671) );
  OAI22X1 U19394 ( .A0(n88), .A1(n1569), .B0(n4175), .B1(n4266), .Y(
        top_core_io_n670) );
  OAI22X1 U19395 ( .A0(n1574), .A1(n88), .B0(n4175), .B1(n4265), .Y(
        top_core_io_n669) );
  OAI22X1 U19396 ( .A0(n1577), .A1(n88), .B0(n4175), .B1(n4264), .Y(
        top_core_io_n668) );
  OAI22X1 U19397 ( .A0(n1578), .A1(n88), .B0(n4175), .B1(n4263), .Y(
        top_core_io_n667) );
  OAI31X1 U19398 ( .A0(top_core_io_n657), .A1(n4262), .A2(n4194), .B0(
        top_core_io_n659), .Y(top_core_io_N92) );
  NAND2X1 U19399 ( .A(top_core_io_N79), .B(top_core_io_n656), .Y(
        top_core_io_n659) );
  OAI31X1 U19400 ( .A0(top_core_io_n657), .A1(n4261), .A2(n4194), .B0(
        top_core_io_n660), .Y(top_core_io_N91) );
  NAND2X1 U19401 ( .A(top_core_io_N80), .B(top_core_io_n656), .Y(
        top_core_io_n660) );
  INVX1 U19402 ( .A(n_ADDR[0]), .Y(n4125) );
  INVX1 U19403 ( .A(n_ADDR[0]), .Y(n4126) );
  OAI22X1 U19404 ( .A0(n4193), .A1(n4262), .B0(top_core_io_n5), .B1(n1572), 
        .Y(top_core_io_n666) );
  OAI22X1 U19405 ( .A0(n4193), .A1(n4261), .B0(top_core_io_n5), .B1(n1575), 
        .Y(top_core_io_n665) );
  INVX1 U19406 ( .A(top_core_io_n5), .Y(n4193) );
  INVX1 U19407 ( .A(n_ADDR[3]), .Y(n4143) );
  AND2X2 U19408 ( .A(top_core_io_N74), .B(top_core_io_n656), .Y(
        top_core_io_N97) );
  AND2X2 U19409 ( .A(top_core_io_N75), .B(top_core_io_n656), .Y(
        top_core_io_N96) );
  AND2X2 U19410 ( .A(top_core_io_N76), .B(top_core_io_n656), .Y(
        top_core_io_N95) );
  AND2X2 U19411 ( .A(top_core_io_N77), .B(top_core_io_n656), .Y(
        top_core_io_N94) );
  AND2X2 U19412 ( .A(top_core_io_N78), .B(top_core_io_n656), .Y(
        top_core_io_N93) );
  INVX1 U19413 ( .A(n_ADDR[0]), .Y(n4127) );
  NAND2X1 U19414 ( .A(n_ADDR[6]), .B(n4192), .Y(top_core_io_n657) );
  CLKINVX3 U19415 ( .A(n_DIN[2]), .Y(n1572) );
  CLKINVX3 U19416 ( .A(n_DIN[1]), .Y(n1575) );
  OAI222X4 U19417 ( .A0(n11629), .A1(n11630), .B0(n11631), .B1(n11632), .C0(
        n1338), .C1(n11633), .Y(top_core_KE_new_sboxw_15_) );
  AOI211X1 U19418 ( .A0(n11654), .A1(n1205), .B0(n11682), .C0(n11683), .Y(
        n11629) );
  AOI211X1 U19419 ( .A0(n6745), .A1(n11634), .B0(n11635), .C0(n11636), .Y(
        n11633) );
  NOR4X1 U19420 ( .A(n11665), .B(n11666), .C(n11667), .D(n11668), .Y(n11631)
         );
  OAI222X4 U19421 ( .A0(n11745), .A1(n11632), .B0(n1338), .B1(n11746), .C0(
        n11747), .C1(n11630), .Y(top_core_KE_new_sboxw_13_) );
  AOI222X1 U19422 ( .A0(n1797), .A1(n11748), .B0(n11749), .B1(n1796), .C0(
        n6826), .C1(n11750), .Y(n11747) );
  AOI22X1 U19423 ( .A0(n1354), .A1(n11754), .B0(n11755), .B1(n1187), .Y(n11746) );
  NOR4BBX1 U19424 ( .AN(n11774), .BN(n11775), .C(n11653), .D(n11642), .Y(
        n11745) );
  OAI222X4 U19425 ( .A0(n11854), .A1(n11630), .B0(n11855), .B1(n11632), .C0(
        n1338), .C1(n11856), .Y(top_core_KE_new_sboxw_10_) );
  AOI221X1 U19426 ( .A0(n11827), .A1(n1805), .B0(top_core_KE_prev_key1_reg_13_), .B1(n11872), .C0(n11873), .Y(n11855) );
  AOI221X1 U19427 ( .A0(n1801), .A1(n11880), .B0(n11881), .B1(n1796), .C0(
        n11882), .Y(n11854) );
  AOI221X1 U19428 ( .A0(n11695), .A1(n11857), .B0(n6746), .B1(n11858), .C0(
        n11859), .Y(n11856) );
  OAI222X4 U19429 ( .A0(top_core_KE_sb1_n54), .A1(top_core_KE_sb1_n55), .B0(
        top_core_KE_sb1_n56), .B1(top_core_KE_sb1_n57), .C0(n1335), .C1(
        top_core_KE_sb1_n58), .Y(top_core_KE_new_sboxw_7_) );
  AOI211X1 U19430 ( .A0(top_core_KE_sb1_n79), .A1(n1196), .B0(
        top_core_KE_sb1_n107), .C0(top_core_KE_sb1_n108), .Y(
        top_core_KE_sb1_n54) );
  AOI211X1 U19431 ( .A0(n6807), .A1(top_core_KE_sb1_n59), .B0(
        top_core_KE_sb1_n60), .C0(top_core_KE_sb1_n61), .Y(top_core_KE_sb1_n58) );
  NOR4X1 U19432 ( .A(top_core_KE_sb1_n90), .B(top_core_KE_sb1_n91), .C(
        top_core_KE_sb1_n92), .D(top_core_KE_sb1_n93), .Y(top_core_KE_sb1_n56)
         );
  OAI222X4 U19433 ( .A0(top_core_KE_sb1_n173), .A1(top_core_KE_sb1_n57), .B0(
        n1335), .B1(top_core_KE_sb1_n174), .C0(top_core_KE_sb1_n175), .C1(
        top_core_KE_sb1_n55), .Y(top_core_KE_new_sboxw_5_) );
  AOI222X1 U19434 ( .A0(n1818), .A1(top_core_KE_sb1_n176), .B0(
        top_core_KE_sb1_n177), .B1(n1817), .C0(n6804), .C1(
        top_core_KE_sb1_n178), .Y(top_core_KE_sb1_n175) );
  AOI22X1 U19435 ( .A0(n1343), .A1(top_core_KE_sb1_n182), .B0(
        top_core_KE_sb1_n183), .B1(n1224), .Y(top_core_KE_sb1_n174) );
  NOR4BBX1 U19436 ( .AN(top_core_KE_sb1_n202), .BN(top_core_KE_sb1_n203), .C(
        top_core_KE_sb1_n78), .D(top_core_KE_sb1_n67), .Y(top_core_KE_sb1_n173) );
  OAI222X4 U19437 ( .A0(top_core_KE_sb1_n283), .A1(top_core_KE_sb1_n55), .B0(
        top_core_KE_sb1_n284), .B1(top_core_KE_sb1_n57), .C0(n1335), .C1(
        top_core_KE_sb1_n285), .Y(top_core_KE_new_sboxw_2_) );
  AOI221X1 U19438 ( .A0(top_core_KE_sb1_n256), .A1(n1826), .B0(
        top_core_KE_prev_key1_reg_5_), .B1(top_core_KE_sb1_n301), .C0(
        top_core_KE_sb1_n302), .Y(top_core_KE_sb1_n284) );
  AOI221X1 U19439 ( .A0(n1822), .A1(top_core_KE_sb1_n309), .B0(
        top_core_KE_sb1_n310), .B1(n1817), .C0(top_core_KE_sb1_n311), .Y(
        top_core_KE_sb1_n283) );
  AOI221X1 U19440 ( .A0(top_core_KE_sb1_n120), .A1(top_core_KE_sb1_n286), .B0(
        n6801), .B1(top_core_KE_sb1_n287), .C0(top_core_KE_sb1_n288), .Y(
        top_core_KE_sb1_n285) );
  OAI222X4 U19441 ( .A0(n12261), .A1(n12262), .B0(n12263), .B1(n12264), .C0(
        n1370), .C1(n12265), .Y(top_core_KE_new_sboxw_31_) );
  AOI211X1 U19442 ( .A0(n12286), .A1(n1165), .B0(n12313), .C0(n12314), .Y(
        n12261) );
  AOI211X1 U19443 ( .A0(n6442), .A1(n12266), .B0(n12267), .C0(n12268), .Y(
        n12265) );
  NOR4X1 U19444 ( .A(n12296), .B(n12297), .C(n12298), .D(n12299), .Y(n12263)
         );
  OAI222X4 U19445 ( .A0(n12376), .A1(n12264), .B0(n1370), .B1(n12377), .C0(
        n12378), .C1(n12262), .Y(top_core_KE_new_sboxw_29_) );
  AOI222X1 U19446 ( .A0(n1758), .A1(n12379), .B0(n12380), .B1(n1753), .C0(
        n6530), .C1(n12381), .Y(n12378) );
  AOI22X1 U19447 ( .A0(n1368), .A1(n12385), .B0(n12386), .B1(n1147), .Y(n12377) );
  NOR4BBX1 U19448 ( .AN(n12405), .BN(n12406), .C(n12285), .D(n12274), .Y(
        n12376) );
  OAI222X4 U19449 ( .A0(n12485), .A1(n12262), .B0(n12486), .B1(n12264), .C0(
        n1370), .C1(n12487), .Y(top_core_KE_new_sboxw_26_) );
  AOI221X1 U19450 ( .A0(n12458), .A1(n1766), .B0(n1755), .B1(n12503), .C0(
        n12504), .Y(n12486) );
  AOI221X1 U19451 ( .A0(n1756), .A1(n12511), .B0(n12512), .B1(n1753), .C0(
        n12513), .Y(n12485) );
  AOI221X1 U19452 ( .A0(n12326), .A1(n12488), .B0(n6443), .B1(n12489), .C0(
        n12490), .Y(n12487) );
  OAI222X4 U19453 ( .A0(n12800), .A1(n12577), .B0(n12801), .B1(n12579), .C0(
        n1336), .C1(n12802), .Y(top_core_KE_new_sboxw_192_2_) );
  AOI221X1 U19454 ( .A0(n12773), .A1(n1743), .B0(n1725), .B1(n12818), .C0(
        n12819), .Y(n12801) );
  AOI221X1 U19455 ( .A0(n1725), .A1(n12826), .B0(n12827), .B1(n1726), .C0(
        n12828), .Y(n12800) );
  AOI221X1 U19456 ( .A0(n12642), .A1(n12803), .B0(n6772), .B1(n12804), .C0(
        n12805), .Y(n12802) );
  OAI222X4 U19457 ( .A0(n13745), .A1(n13522), .B0(n13746), .B1(n13524), .C0(
        n1341), .C1(n13747), .Y(top_core_KE_new_sboxw_192_26_) );
  AOI221X1 U19458 ( .A0(n13718), .A1(n1657), .B0(n1638), .B1(n13763), .C0(
        n13764), .Y(n13746) );
  AOI221X1 U19459 ( .A0(n1641), .A1(n13771), .B0(n13772), .B1(n1636), .C0(
        n13773), .Y(n13745) );
  AOI221X1 U19460 ( .A0(n13587), .A1(n13748), .B0(n6434), .B1(n13749), .C0(
        n13750), .Y(n13747) );
  OAI222X4 U19461 ( .A0(n12692), .A1(n12579), .B0(n1336), .B1(n12693), .C0(
        n12694), .C1(n12577), .Y(top_core_KE_new_sboxw_192_5_) );
  AOI222X1 U19462 ( .A0(n1725), .A1(n12695), .B0(n12696), .B1(n1729), .C0(
        n6775), .C1(n12697), .Y(n12694) );
  AOI22X1 U19463 ( .A0(n1342), .A1(n12701), .B0(n12702), .B1(n1225), .Y(n12693) );
  NOR4BBX1 U19464 ( .AN(n12721), .BN(n12722), .C(n12600), .D(n12589), .Y(
        n12692) );
  OAI222X4 U19465 ( .A0(n13637), .A1(n13524), .B0(n1341), .B1(n13638), .C0(
        n13639), .C1(n13522), .Y(top_core_KE_new_sboxw_192_29_) );
  AOI222X1 U19466 ( .A0(n1641), .A1(n13640), .B0(n13641), .B1(n1636), .C0(
        n6519), .C1(n13642), .Y(n13639) );
  AOI22X1 U19467 ( .A0(n1369), .A1(n13646), .B0(n13647), .B1(n1146), .Y(n13638) );
  NOR4BBX1 U19468 ( .AN(n13666), .BN(n13667), .C(n13545), .D(n13534), .Y(
        n13637) );
  OAI222X4 U19469 ( .A0(n13115), .A1(n12892), .B0(n13116), .B1(n12894), .C0(
        n1337), .C1(n13117), .Y(top_core_KE_new_sboxw_192_10_) );
  AOI221X1 U19470 ( .A0(n13088), .A1(n1714), .B0(n1696), .B1(n13133), .C0(
        n13134), .Y(n13116) );
  AOI221X1 U19471 ( .A0(n1696), .A1(n13141), .B0(n13142), .B1(n1697), .C0(
        n13143), .Y(n13115) );
  AOI221X1 U19472 ( .A0(n12957), .A1(n13118), .B0(n6715), .B1(n13119), .C0(
        n13120), .Y(n13117) );
  OAI222X4 U19473 ( .A0(n13007), .A1(n12894), .B0(n1337), .B1(n13008), .C0(
        n13009), .C1(n12892), .Y(top_core_KE_new_sboxw_192_13_) );
  AOI222X1 U19474 ( .A0(n1696), .A1(n13010), .B0(n13011), .B1(n1700), .C0(
        n6815), .C1(n13012), .Y(n13009) );
  AOI22X1 U19475 ( .A0(n1355), .A1(n13016), .B0(n13017), .B1(n1186), .Y(n13008) );
  NOR4BBX1 U19476 ( .AN(n13036), .BN(n13037), .C(n12915), .D(n12904), .Y(
        n13007) );
  OAI222X4 U19477 ( .A0(n12891), .A1(n12892), .B0(n12893), .B1(n12894), .C0(
        n1337), .C1(n12895), .Y(top_core_KE_new_sboxw_192_15_) );
  AOI211X1 U19478 ( .A0(n12916), .A1(n1201), .B0(n12944), .C0(n12945), .Y(
        n12891) );
  AOI211X1 U19479 ( .A0(n6714), .A1(n12896), .B0(n12897), .C0(n12898), .Y(
        n12895) );
  NOR4X1 U19480 ( .A(n12927), .B(n12928), .C(n12929), .D(n12930), .Y(n12893)
         );
  OAI222X4 U19481 ( .A0(n13521), .A1(n13522), .B0(n13523), .B1(n13524), .C0(
        n1341), .C1(n13525), .Y(top_core_KE_new_sboxw_192_31_) );
  AOI211X1 U19482 ( .A0(n13546), .A1(n1161), .B0(n13574), .C0(n13575), .Y(
        n13521) );
  AOI211X1 U19483 ( .A0(n6433), .A1(n13526), .B0(n13527), .C0(n13528), .Y(
        n13525) );
  NOR4X1 U19484 ( .A(n13557), .B(n13558), .C(n13559), .D(n13560), .Y(n13523)
         );
  OAI222X4 U19485 ( .A0(n12576), .A1(n12577), .B0(n12578), .B1(n12579), .C0(
        n1336), .C1(n12580), .Y(top_core_KE_new_sboxw_192_7_) );
  AOI211X1 U19486 ( .A0(n12601), .A1(n1192), .B0(n12629), .C0(n12630), .Y(
        n12576) );
  AOI211X1 U19487 ( .A0(n6778), .A1(n12581), .B0(n12582), .C0(n12583), .Y(
        n12580) );
  NOR4X1 U19488 ( .A(n12612), .B(n12613), .C(n12614), .D(n12615), .Y(n12578)
         );
  OAI222X4 U19489 ( .A0(n11945), .A1(n11946), .B0(n11947), .B1(n11948), .C0(
        n1339), .C1(n11949), .Y(top_core_KE_new_sboxw_23_) );
  AOI211X1 U19490 ( .A0(n11970), .A1(n1156), .B0(n11998), .C0(n11999), .Y(
        n11945) );
  AOI211X1 U19491 ( .A0(n6510), .A1(n11950), .B0(n11951), .C0(n11952), .Y(
        n11949) );
  NOR4X1 U19492 ( .A(n11981), .B(n11982), .C(n11983), .D(n11984), .Y(n11947)
         );
  OAI222X4 U19493 ( .A0(n12061), .A1(n11948), .B0(n1339), .B1(n12062), .C0(
        n12063), .C1(n11946), .Y(top_core_KE_new_sboxw_21_) );
  AOI222X1 U19494 ( .A0(n1776), .A1(n12064), .B0(n12065), .B1(n1775), .C0(
        n6507), .C1(n12066), .Y(n12063) );
  AOI22X1 U19495 ( .A0(n1357), .A1(n12070), .B0(n12071), .B1(n1184), .Y(n12062) );
  NOR4BBX1 U19496 ( .AN(n12090), .BN(n12091), .C(n11969), .D(n11958), .Y(
        n12061) );
  OAI222X4 U19497 ( .A0(n12170), .A1(n11946), .B0(n12171), .B1(n11948), .C0(
        n1339), .C1(n12172), .Y(top_core_KE_new_sboxw_18_) );
  AOI221X1 U19498 ( .A0(n12143), .A1(n1784), .B0(top_core_KE_prev_key1_reg_21_), .B1(n12188), .C0(n12189), .Y(n12171) );
  AOI221X1 U19499 ( .A0(n1780), .A1(n12196), .B0(n12197), .B1(n1775), .C0(
        n12198), .Y(n12170) );
  AOI221X1 U19500 ( .A0(n12011), .A1(n12173), .B0(n6504), .B1(n12174), .C0(
        n12175), .Y(n12172) );
  OAI22X2 U19501 ( .A0(n1338), .A1(n11692), .B0(n11693), .B1(n6993), .Y(
        top_core_KE_new_sboxw_14_) );
  AOI211X1 U19502 ( .A0(n11721), .A1(n1187), .B0(n11722), .C0(n11723), .Y(
        n11692) );
  AOI221X1 U19503 ( .A0(n1354), .A1(n11694), .B0(n11695), .B1(n11696), .C0(
        n11697), .Y(n11693) );
  OAI22X1 U19504 ( .A0(n1187), .A1(n11728), .B0(n11729), .B1(n11730), .Y(
        n11722) );
  OAI22X2 U19505 ( .A0(n11915), .A1(n6993), .B0(n1338), .B1(n11916), .Y(
        top_core_KE_new_sboxw_8_) );
  AOI222X1 U19506 ( .A0(n11932), .A1(n1187), .B0(n6746), .B1(n11933), .C0(
        n1354), .C1(n11934), .Y(n11915) );
  AOI22X1 U19507 ( .A0(n1354), .A1(n11917), .B0(n11918), .B1(n1187), .Y(n11916) );
  OAI21XL U19508 ( .A0(n11935), .A1(n1795), .B0(n11936), .Y(n11934) );
  OAI22X2 U19509 ( .A0(n1335), .A1(top_core_KE_sb1_n117), .B0(
        top_core_KE_sb1_n118), .B1(n6997), .Y(top_core_KE_new_sboxw_6_) );
  AOI211X1 U19510 ( .A0(top_core_KE_sb1_n148), .A1(n1224), .B0(
        top_core_KE_sb1_n149), .C0(top_core_KE_sb1_n150), .Y(
        top_core_KE_sb1_n117) );
  AOI221X1 U19511 ( .A0(n1343), .A1(top_core_KE_sb1_n119), .B0(
        top_core_KE_sb1_n120), .B1(top_core_KE_sb1_n121), .C0(
        top_core_KE_sb1_n122), .Y(top_core_KE_sb1_n118) );
  OAI22X1 U19512 ( .A0(n1224), .A1(top_core_KE_sb1_n155), .B0(
        top_core_KE_sb1_n156), .B1(top_core_KE_sb1_n157), .Y(
        top_core_KE_sb1_n149) );
  OAI22X2 U19513 ( .A0(top_core_KE_sb1_n344), .A1(n6997), .B0(n1335), .B1(
        top_core_KE_sb1_n345), .Y(top_core_KE_new_sboxw_0_) );
  AOI222X1 U19514 ( .A0(top_core_KE_sb1_n361), .A1(n1224), .B0(n6801), .B1(
        top_core_KE_sb1_n362), .C0(n1343), .C1(top_core_KE_sb1_n363), .Y(
        top_core_KE_sb1_n344) );
  AOI22X1 U19515 ( .A0(n1343), .A1(top_core_KE_sb1_n346), .B0(
        top_core_KE_sb1_n347), .B1(n1224), .Y(top_core_KE_sb1_n345) );
  OAI21XL U19516 ( .A0(top_core_KE_sb1_n364), .A1(n1816), .B0(
        top_core_KE_sb1_n365), .Y(top_core_KE_sb1_n363) );
  OAI22X2 U19517 ( .A0(n1370), .A1(n12323), .B0(n12324), .B1(n6358), .Y(
        top_core_KE_new_sboxw_30_) );
  AOI211X1 U19518 ( .A0(n12352), .A1(n1147), .B0(n12353), .C0(n12354), .Y(
        n12323) );
  AOI221X1 U19519 ( .A0(n1368), .A1(n12325), .B0(n12326), .B1(n12327), .C0(
        n12328), .Y(n12324) );
  OAI22X1 U19520 ( .A0(n1147), .A1(n12359), .B0(n12360), .B1(n12361), .Y(
        n12353) );
  OAI22X2 U19521 ( .A0(n12546), .A1(n6358), .B0(n1370), .B1(n12547), .Y(
        top_core_KE_new_sboxw_24_) );
  AOI222X1 U19522 ( .A0(n12563), .A1(n1147), .B0(n6443), .B1(n12564), .C0(
        n1368), .C1(n12565), .Y(n12546) );
  AOI22X1 U19523 ( .A0(n1368), .A1(n12548), .B0(n12549), .B1(n1147), .Y(n12547) );
  OAI21XL U19524 ( .A0(n12566), .A1(n1752), .B0(n12567), .Y(n12565) );
  OAI2BB2X2 U19525 ( .B0(n1338), .B1(n11887), .A0N(n1338), .A1N(n11888), .Y(
        top_core_KE_new_sboxw_9_) );
  AOI222X1 U19526 ( .A0(n11903), .A1(n1187), .B0(n6745), .B1(n11904), .C0(
        n6746), .C1(n11905), .Y(n11887) );
  OAI221XL U19527 ( .A0(n11889), .A1(n11640), .B0(n1354), .B1(n11890), .C0(
        n11891), .Y(n11888) );
  NAND4X1 U19528 ( .A(n11910), .B(n11911), .C(n11912), .D(n11913), .Y(n11903)
         );
  OAI2BB2X2 U19529 ( .B0(n1335), .B1(top_core_KE_sb1_n316), .A0N(n1335), .A1N(
        top_core_KE_sb1_n317), .Y(top_core_KE_new_sboxw_1_) );
  AOI222X1 U19530 ( .A0(top_core_KE_sb1_n332), .A1(n1224), .B0(n6807), .B1(
        top_core_KE_sb1_n333), .C0(n6801), .C1(top_core_KE_sb1_n334), .Y(
        top_core_KE_sb1_n316) );
  OAI221XL U19531 ( .A0(top_core_KE_sb1_n318), .A1(top_core_KE_sb1_n65), .B0(
        n1343), .B1(top_core_KE_sb1_n319), .C0(top_core_KE_sb1_n320), .Y(
        top_core_KE_sb1_n317) );
  NAND4X1 U19532 ( .A(top_core_KE_sb1_n339), .B(top_core_KE_sb1_n340), .C(
        top_core_KE_sb1_n341), .D(top_core_KE_sb1_n342), .Y(
        top_core_KE_sb1_n332) );
  OAI2BB2X2 U19533 ( .B0(n1370), .B1(n12518), .A0N(n1370), .A1N(n12519), .Y(
        top_core_KE_new_sboxw_25_) );
  AOI222X1 U19534 ( .A0(n12534), .A1(n1147), .B0(n6442), .B1(n12535), .C0(
        n6443), .C1(n12536), .Y(n12518) );
  OAI221XL U19535 ( .A0(n12520), .A1(n12272), .B0(n1368), .B1(n12521), .C0(
        n12522), .Y(n12519) );
  NAND4X1 U19536 ( .A(n12541), .B(n12542), .C(n12543), .D(n12544), .Y(n12534)
         );
  OAI21X2 U19537 ( .A0(n11782), .A1(n6993), .B0(n11783), .Y(
        top_core_KE_new_sboxw_12_) );
  AOI222X1 U19538 ( .A0(n1354), .A1(n11801), .B0(n6731), .B1(n11802), .C0(
        n11695), .C1(n11803), .Y(n11782) );
  OAI2BB1X1 U19539 ( .A0N(n11784), .A1N(n11785), .B0(n6993), .Y(n11783) );
  NAND4X1 U19540 ( .A(n11807), .B(n11808), .C(n11809), .D(n11810), .Y(n11802)
         );
  OAI21X2 U19541 ( .A0(n1338), .A1(n11820), .B0(n11821), .Y(
        top_core_KE_new_sboxw_11_) );
  AOI211X1 U19542 ( .A0(n11695), .A1(n11840), .B0(n6744), .C0(n11841), .Y(
        n11820) );
  AOI21X1 U19543 ( .A0(n6743), .A1(n11822), .B0(n11823), .Y(n11821) );
  INVX1 U19544 ( .A(n11845), .Y(n6744) );
  OAI21X2 U19545 ( .A0(top_core_KE_sb1_n210), .A1(n6997), .B0(
        top_core_KE_sb1_n211), .Y(top_core_KE_new_sboxw_4_) );
  AOI222X1 U19546 ( .A0(n1343), .A1(top_core_KE_sb1_n229), .B0(n6794), .B1(
        top_core_KE_sb1_n230), .C0(top_core_KE_sb1_n120), .C1(
        top_core_KE_sb1_n231), .Y(top_core_KE_sb1_n210) );
  OAI2BB1X1 U19547 ( .A0N(top_core_KE_sb1_n212), .A1N(top_core_KE_sb1_n213), 
        .B0(n6997), .Y(top_core_KE_sb1_n211) );
  NAND4X1 U19548 ( .A(top_core_KE_sb1_n235), .B(top_core_KE_sb1_n236), .C(
        top_core_KE_sb1_n237), .D(top_core_KE_sb1_n238), .Y(
        top_core_KE_sb1_n230) );
  OAI21X2 U19549 ( .A0(n1335), .A1(top_core_KE_sb1_n249), .B0(
        top_core_KE_sb1_n250), .Y(top_core_KE_new_sboxw_3_) );
  AOI211X1 U19550 ( .A0(top_core_KE_sb1_n120), .A1(top_core_KE_sb1_n269), .B0(
        n6800), .C0(top_core_KE_sb1_n270), .Y(top_core_KE_sb1_n249) );
  AOI21X1 U19551 ( .A0(n6986), .A1(top_core_KE_sb1_n251), .B0(
        top_core_KE_sb1_n252), .Y(top_core_KE_sb1_n250) );
  INVX1 U19552 ( .A(top_core_KE_sb1_n274), .Y(n6800) );
  OAI21X2 U19553 ( .A0(n12413), .A1(n6358), .B0(n12414), .Y(
        top_core_KE_new_sboxw_28_) );
  AOI222X1 U19554 ( .A0(n1368), .A1(n12432), .B0(n6439), .B1(n12433), .C0(
        n12326), .C1(n12434), .Y(n12413) );
  OAI2BB1X1 U19555 ( .A0N(n12415), .A1N(n12416), .B0(n6358), .Y(n12414) );
  NAND4X1 U19556 ( .A(n12438), .B(n12439), .C(n12440), .D(n12441), .Y(n12433)
         );
  OAI21X2 U19557 ( .A0(n1370), .A1(n12451), .B0(n12452), .Y(
        top_core_KE_new_sboxw_27_) );
  AOI211X1 U19558 ( .A0(n12326), .A1(n12471), .B0(n6441), .C0(n12472), .Y(
        n12451) );
  AOI21X1 U19559 ( .A0(n6372), .A1(n12453), .B0(n12454), .Y(n12452) );
  INVX1 U19560 ( .A(n12476), .Y(n6441) );
  NOR2X2 U19561 ( .A(n7023), .B(n7022), .Y(top_core_KE_n896) );
  OAI22X2 U19562 ( .A0(n1341), .A1(n13584), .B0(n13585), .B1(n6989), .Y(
        top_core_KE_new_sboxw_192_30_) );
  AOI211X1 U19563 ( .A0(n13613), .A1(n1146), .B0(n13614), .C0(n13615), .Y(
        n13584) );
  AOI221X1 U19564 ( .A0(n1369), .A1(n13586), .B0(n13587), .B1(n13588), .C0(
        n13589), .Y(n13585) );
  OAI22X1 U19565 ( .A0(n1146), .A1(n13620), .B0(n13621), .B1(n13622), .Y(
        n13614) );
  OAI22X2 U19566 ( .A0(n12861), .A1(n6995), .B0(n1336), .B1(n12862), .Y(
        top_core_KE_new_sboxw_192_0_) );
  AOI222X1 U19567 ( .A0(n12878), .A1(n1225), .B0(n6772), .B1(n12879), .C0(
        n1342), .C1(n12880), .Y(n12861) );
  AOI22X1 U19568 ( .A0(n1342), .A1(n12863), .B0(n12864), .B1(n1225), .Y(n12862) );
  OAI21XL U19569 ( .A0(n12881), .A1(n1727), .B0(n12882), .Y(n12880) );
  OAI22X2 U19570 ( .A0(n13806), .A1(n6989), .B0(n1341), .B1(n13807), .Y(
        top_core_KE_new_sboxw_192_24_) );
  AOI222X1 U19571 ( .A0(n13823), .A1(n1146), .B0(n6434), .B1(n13824), .C0(
        n1369), .C1(n13825), .Y(n13806) );
  AOI22X1 U19572 ( .A0(n1369), .A1(n13808), .B0(n13809), .B1(n1146), .Y(n13807) );
  OAI21XL U19573 ( .A0(n13826), .A1(n1635), .B0(n13827), .Y(n13825) );
  OAI22X2 U19574 ( .A0(n1336), .A1(n12639), .B0(n12640), .B1(n6995), .Y(
        top_core_KE_new_sboxw_192_6_) );
  AOI211X1 U19575 ( .A0(n12668), .A1(n1225), .B0(n12669), .C0(n12670), .Y(
        n12639) );
  AOI221X1 U19576 ( .A0(n1342), .A1(n12641), .B0(n12642), .B1(n12643), .C0(
        n12644), .Y(n12640) );
  OAI22X1 U19577 ( .A0(n1225), .A1(n12675), .B0(n12676), .B1(n12677), .Y(
        n12669) );
  OAI22X2 U19578 ( .A0(n13176), .A1(n6994), .B0(n1337), .B1(n13177), .Y(
        top_core_KE_new_sboxw_192_8_) );
  AOI222X1 U19579 ( .A0(n13193), .A1(n1186), .B0(n6715), .B1(n13194), .C0(
        n1355), .C1(n13195), .Y(n13176) );
  AOI22X1 U19580 ( .A0(n1355), .A1(n13178), .B0(n13179), .B1(n1186), .Y(n13177) );
  OAI21XL U19581 ( .A0(n13196), .A1(n1698), .B0(n13197), .Y(n13195) );
  OAI22X2 U19582 ( .A0(n1337), .A1(n12954), .B0(n12955), .B1(n6994), .Y(
        top_core_KE_new_sboxw_192_14_) );
  AOI211X1 U19583 ( .A0(n12983), .A1(n1186), .B0(n12984), .C0(n12985), .Y(
        n12954) );
  AOI221X1 U19584 ( .A0(n1355), .A1(n12956), .B0(n12957), .B1(n12958), .C0(
        n12959), .Y(n12955) );
  OAI22X1 U19585 ( .A0(n1186), .A1(n12990), .B0(n12991), .B1(n12992), .Y(
        n12984) );
  NOR3X2 U19586 ( .A(n7016), .B(n1334), .C(n7014), .Y(top_core_KE_n875) );
  NOR3X2 U19587 ( .A(n7016), .B(n1332), .C(n1226), .Y(top_core_KE_n878) );
  OAI2BB2X2 U19588 ( .B0(n1336), .B1(n12833), .A0N(n1336), .A1N(n12834), .Y(
        top_core_KE_new_sboxw_192_1_) );
  AOI222X1 U19589 ( .A0(n12849), .A1(n1225), .B0(n6778), .B1(n12850), .C0(
        n6772), .C1(n12851), .Y(n12833) );
  OAI221XL U19590 ( .A0(n12835), .A1(n12587), .B0(n1342), .B1(n12836), .C0(
        n12837), .Y(n12834) );
  NAND4X1 U19591 ( .A(n12856), .B(n12857), .C(n12858), .D(n12859), .Y(n12849)
         );
  OAI2BB2X2 U19592 ( .B0(n1341), .B1(n13778), .A0N(n1341), .A1N(n13779), .Y(
        top_core_KE_new_sboxw_192_25_) );
  AOI222X1 U19593 ( .A0(n13794), .A1(n1146), .B0(n6433), .B1(n13795), .C0(
        n6434), .C1(n13796), .Y(n13778) );
  OAI221XL U19594 ( .A0(n13780), .A1(n13532), .B0(n1369), .B1(n13781), .C0(
        n13782), .Y(n13779) );
  NAND4X1 U19595 ( .A(n13801), .B(n13802), .C(n13803), .D(n13804), .Y(n13794)
         );
  OAI2BB2X2 U19596 ( .B0(n1337), .B1(n13148), .A0N(n1337), .A1N(n13149), .Y(
        top_core_KE_new_sboxw_192_9_) );
  AOI222X1 U19597 ( .A0(n13164), .A1(n1186), .B0(n6714), .B1(n13165), .C0(
        n6715), .C1(n13166), .Y(n13148) );
  OAI221XL U19598 ( .A0(n13150), .A1(n12902), .B0(n1355), .B1(n13151), .C0(
        n13152), .Y(n13149) );
  NAND4X1 U19599 ( .A(n13171), .B(n13172), .C(n13173), .D(n13174), .Y(n13164)
         );
  OAI21X2 U19600 ( .A0(n13673), .A1(n6989), .B0(n13674), .Y(
        top_core_KE_new_sboxw_192_28_) );
  AOI222X1 U19601 ( .A0(n1369), .A1(n13692), .B0(n6419), .B1(n13693), .C0(
        n13587), .C1(n13694), .Y(n13673) );
  OAI2BB1X1 U19602 ( .A0N(n13675), .A1N(n13676), .B0(n6989), .Y(n13674) );
  NAND4X1 U19603 ( .A(n13698), .B(n13699), .C(n13700), .D(n13701), .Y(n13693)
         );
  OAI21X2 U19604 ( .A0(n12728), .A1(n6995), .B0(n12729), .Y(
        top_core_KE_new_sboxw_192_4_) );
  AOI222X1 U19605 ( .A0(n1342), .A1(n12747), .B0(n6763), .B1(n12748), .C0(
        n12642), .C1(n12749), .Y(n12728) );
  OAI2BB1X1 U19606 ( .A0N(n12730), .A1N(n12731), .B0(n6995), .Y(n12729) );
  NAND4X1 U19607 ( .A(n12753), .B(n12754), .C(n12755), .D(n12756), .Y(n12748)
         );
  OAI21X2 U19608 ( .A0(n13043), .A1(n6994), .B0(n13044), .Y(
        top_core_KE_new_sboxw_192_12_) );
  AOI222X1 U19609 ( .A0(n1355), .A1(n13062), .B0(n6706), .B1(n13063), .C0(
        n12957), .C1(n13064), .Y(n13043) );
  OAI2BB1X1 U19610 ( .A0N(n13045), .A1N(n13046), .B0(n6994), .Y(n13044) );
  NAND4X1 U19611 ( .A(n13068), .B(n13069), .C(n13070), .D(n13071), .Y(n13063)
         );
  OAI21X2 U19612 ( .A0(n1336), .A1(n12766), .B0(n12767), .Y(
        top_core_KE_new_sboxw_192_3_) );
  AOI211X1 U19613 ( .A0(n12642), .A1(n12786), .B0(n6771), .C0(n12787), .Y(
        n12766) );
  AOI21X1 U19614 ( .A0(n6988), .A1(n12768), .B0(n12769), .Y(n12767) );
  INVX1 U19615 ( .A(n12791), .Y(n6771) );
  OAI21X2 U19616 ( .A0(n1341), .A1(n13711), .B0(n13712), .Y(
        top_core_KE_new_sboxw_192_27_) );
  AOI211X1 U19617 ( .A0(n13587), .A1(n13731), .B0(n6432), .C0(n13732), .Y(
        n13711) );
  AOI21X1 U19618 ( .A0(n6431), .A1(n13713), .B0(n13714), .Y(n13712) );
  INVX1 U19619 ( .A(n13736), .Y(n6432) );
  OAI21X2 U19620 ( .A0(n1337), .A1(n13081), .B0(n13082), .Y(
        top_core_KE_new_sboxw_192_11_) );
  AOI211X1 U19621 ( .A0(n12957), .A1(n13101), .B0(n6713), .C0(n13102), .Y(
        n13081) );
  AOI21X1 U19622 ( .A0(n6712), .A1(n13083), .B0(n13084), .Y(n13082) );
  INVX1 U19623 ( .A(n13106), .Y(n6713) );
  OAI22X2 U19624 ( .A0(n1339), .A1(n12008), .B0(n12009), .B1(n6992), .Y(
        top_core_KE_new_sboxw_22_) );
  AOI211X1 U19625 ( .A0(n12037), .A1(n1184), .B0(n12038), .C0(n12039), .Y(
        n12008) );
  AOI221X1 U19626 ( .A0(n1357), .A1(n12010), .B0(n12011), .B1(n12012), .C0(
        n12013), .Y(n12009) );
  OAI22X1 U19627 ( .A0(n1184), .A1(n12044), .B0(n12045), .B1(n12046), .Y(
        n12038) );
  OAI22X2 U19628 ( .A0(n12231), .A1(n6992), .B0(n1339), .B1(n12232), .Y(
        top_core_KE_new_sboxw_16_) );
  AOI222X1 U19629 ( .A0(n12248), .A1(n1184), .B0(n6504), .B1(n12249), .C0(
        n1357), .C1(n12250), .Y(n12231) );
  AOI22X1 U19630 ( .A0(n1357), .A1(n12233), .B0(n12234), .B1(n1184), .Y(n12232) );
  OAI21XL U19631 ( .A0(n12251), .A1(n1774), .B0(n12252), .Y(n12250) );
  NAND2X2 U19632 ( .A(n6915), .B(n1344), .Y(n11716) );
  NAND2X2 U19633 ( .A(n6869), .B(n1345), .Y(top_core_KE_sb1_n143) );
  NAND2X2 U19634 ( .A(n6622), .B(n1358), .Y(n12347) );
  NAND2X2 U19635 ( .A(n6575), .B(n1359), .Y(n12032) );
  OAI222XL U19636 ( .A0(top_core_KE_n2703), .A1(top_core_KE_n2509), .B0(n1866), 
        .B1(top_core_KE_n2712), .C0(n738), .C1(n7020), .Y(top_core_KE_n2696)
         );
  NAND2X1 U19637 ( .A(top_core_KE_n896), .B(top_core_KE_Nk0_0_), .Y(
        top_core_KE_n2712) );
  OAI2BB2X2 U19638 ( .B0(n1339), .B1(n12203), .A0N(n1339), .A1N(n12204), .Y(
        top_core_KE_new_sboxw_17_) );
  AOI222X1 U19639 ( .A0(n12219), .A1(n1184), .B0(n6510), .B1(n12220), .C0(
        n6504), .C1(n12221), .Y(n12203) );
  OAI221XL U19640 ( .A0(n12205), .A1(n11956), .B0(n1357), .B1(n12206), .C0(
        n12207), .Y(n12204) );
  NAND4X1 U19641 ( .A(n12226), .B(n12227), .C(n12228), .D(n12229), .Y(n12219)
         );
  OAI21X2 U19642 ( .A0(n12098), .A1(n6992), .B0(n12099), .Y(
        top_core_KE_new_sboxw_20_) );
  AOI222X1 U19643 ( .A0(n1357), .A1(n12117), .B0(n6495), .B1(n12118), .C0(
        n12011), .C1(n12119), .Y(n12098) );
  OAI2BB1X1 U19644 ( .A0N(n12100), .A1N(n12101), .B0(n6992), .Y(n12099) );
  NAND4X1 U19645 ( .A(n12123), .B(n12124), .C(n12125), .D(n12126), .Y(n12118)
         );
  OAI21X2 U19646 ( .A0(n1339), .A1(n12136), .B0(n12137), .Y(
        top_core_KE_new_sboxw_19_) );
  AOI211X1 U19647 ( .A0(n12011), .A1(n12156), .B0(n6503), .C0(n12157), .Y(
        n12136) );
  AOI21X1 U19648 ( .A0(n6699), .A1(n12138), .B0(n12139), .Y(n12137) );
  INVX1 U19649 ( .A(n12161), .Y(n6503) );
  NOR3X1 U19650 ( .A(top_core_KE_n1866), .B(top_core_KE_n1865), .C(n7021), .Y(
        top_core_KE_n1864) );
  NOR2X2 U19651 ( .A(n1678), .B(n1363), .Y(n13373) );
  NOR2X2 U19652 ( .A(n1737), .B(n1349), .Y(n12743) );
  NOR2X2 U19653 ( .A(n1643), .B(n1361), .Y(n13688) );
  NOR2X2 U19654 ( .A(n1708), .B(n1347), .Y(n13058) );
  NOR2X2 U19655 ( .A(n6964), .B(n1346), .Y(n11797) );
  NOR2X2 U19656 ( .A(n6958), .B(n1348), .Y(top_core_KE_sb1_n225) );
  NOR2X2 U19657 ( .A(n6670), .B(n1362), .Y(n12113) );
  NOR2X2 U19658 ( .A(n1171), .B(n1360), .Y(n12428) );
  NOR2X2 U19659 ( .A(n1669), .B(n1356), .Y(n13272) );
  NOR2X2 U19660 ( .A(n1727), .B(n1342), .Y(n12642) );
  NOR2X2 U19661 ( .A(n1698), .B(n1355), .Y(n12957) );
  NOR2X2 U19662 ( .A(n1635), .B(n1369), .Y(n13587) );
  NOR2X2 U19663 ( .A(n1752), .B(n1368), .Y(n12326) );
  NOR2X2 U19664 ( .A(n1795), .B(n1354), .Y(n11695) );
  NOR2X2 U19665 ( .A(n1816), .B(n1343), .Y(top_core_KE_sb1_n120) );
  NOR2X2 U19666 ( .A(n1774), .B(n1357), .Y(n12011) );
  NOR2X1 U19667 ( .A(n1333), .B(n1332), .Y(top_core_KE_n883) );
  AOI22X1 U19668 ( .A0(n1211), .A1(n1811), .B0(n1344), .B1(n625), .Y(n11717)
         );
  AOI22X1 U19669 ( .A0(n1210), .A1(n1832), .B0(n1345), .B1(n626), .Y(
        top_core_KE_sb1_n144) );
  AOI22X1 U19670 ( .A0(n1171), .A1(n1769), .B0(n1358), .B1(n627), .Y(n12348)
         );
  AOI22X1 U19671 ( .A0(n1170), .A1(n1790), .B0(n1359), .B1(n628), .Y(n12033)
         );
  XOR2X1 U19672 ( .A(top_core_KE_new_sboxw_23_), .B(n7006), .Y(
        top_core_KE_n2183) );
  NOR2X1 U19673 ( .A(n1673), .B(n1363), .Y(n13240) );
  NOR2X1 U19674 ( .A(n1702), .B(n1347), .Y(n12925) );
  NOR2X1 U19675 ( .A(n1731), .B(n1349), .Y(n12610) );
  NOR2X1 U19676 ( .A(n1646), .B(n1361), .Y(n13555) );
  NOR2X1 U19677 ( .A(n1358), .B(n1360), .Y(n12294) );
  NOR2X1 U19678 ( .A(n1344), .B(n1346), .Y(n11663) );
  NOR2X1 U19679 ( .A(n1345), .B(n1348), .Y(top_core_KE_sb1_n88) );
  NOR2X1 U19680 ( .A(n1359), .B(n1362), .Y(n11979) );
  NOR2X1 U19681 ( .A(n1169), .B(n1358), .Y(n12442) );
  NOR2X1 U19682 ( .A(n1209), .B(n1344), .Y(n11811) );
  NOR2X1 U19683 ( .A(n1207), .B(n1345), .Y(top_core_KE_sb1_n239) );
  NOR2X1 U19684 ( .A(n1167), .B(n1359), .Y(n12127) );
  AND2X2 U19685 ( .A(top_core_KE_n894), .B(top_core_KE_n1865), .Y(
        top_core_KE_n907) );
  AND2X2 U19686 ( .A(top_core_KE_n1870), .B(top_core_KE_n894), .Y(
        top_core_KE_n910) );
  AND2X2 U19687 ( .A(top_core_KE_n2699), .B(top_core_KE_n894), .Y(
        top_core_KE_n1877) );
  AND2X2 U19688 ( .A(top_core_KE_n2700), .B(n7011), .Y(top_core_KE_n1875) );
  CLKINVX3 U19689 ( .A(top_core_KE_n2705), .Y(n7016) );
  XNOR2X1 U19690 ( .A(n6337), .B(top_core_KE_n1909), .Y(top_core_KE_n1975) );
  XNOR2X1 U19691 ( .A(n6396), .B(top_core_KE_n1927), .Y(top_core_KE_n2009) );
  XNOR2X1 U19692 ( .A(n6535), .B(top_core_KE_n1931), .Y(top_core_KE_n2015) );
  XNOR2X1 U19693 ( .A(n6630), .B(top_core_KE_n1933), .Y(top_core_KE_n2018) );
  XNOR2X1 U19694 ( .A(n6678), .B(top_core_KE_n1937), .Y(top_core_KE_n2024) );
  XNOR2X1 U19695 ( .A(n6685), .B(top_core_KE_n1939), .Y(top_core_KE_n2027) );
  XNOR2X1 U19696 ( .A(n6388), .B(top_core_KE_n1943), .Y(top_core_KE_n2033) );
  XNOR2X1 U19697 ( .A(n6877), .B(top_core_KE_n1947), .Y(top_core_KE_n2039) );
  XNOR2X1 U19698 ( .A(n6938), .B(top_core_KE_n1949), .Y(top_core_KE_n2042) );
  XNOR2X1 U19699 ( .A(n6970), .B(top_core_KE_n1953), .Y(top_core_KE_n2048) );
  XNOR2X1 U19700 ( .A(n6980), .B(top_core_KE_n1955), .Y(top_core_KE_n2051) );
  XNOR2X1 U19701 ( .A(n6380), .B(top_core_KE_n1959), .Y(top_core_KE_n2057) );
  XNOR2X1 U19702 ( .A(n6831), .B(top_core_KE_n1963), .Y(top_core_KE_n2063) );
  XNOR2X1 U19703 ( .A(n6923), .B(top_core_KE_n1965), .Y(top_core_KE_n2066) );
  XNOR2X1 U19704 ( .A(n6965), .B(top_core_KE_n1969), .Y(top_core_KE_n2072) );
  XNOR2X1 U19705 ( .A(n6975), .B(top_core_KE_n1971), .Y(top_core_KE_n2075) );
  XNOR2X1 U19706 ( .A(n6959), .B(top_core_KE_n1951), .Y(top_core_KE_n2045) );
  XNOR2X1 U19707 ( .A(n6953), .B(top_core_KE_n1967), .Y(top_core_KE_n2069) );
  XNOR2X1 U19708 ( .A(n6810), .B(top_core_KE_n1945), .Y(top_core_KE_n2036) );
  XNOR2X1 U19709 ( .A(n6747), .B(top_core_KE_n1961), .Y(top_core_KE_n2060) );
  XNOR2X1 U19710 ( .A(n6663), .B(top_core_KE_n1935), .Y(top_core_KE_n2021) );
  XNOR2X1 U19711 ( .A(n6444), .B(top_core_KE_n1929), .Y(top_core_KE_n2012) );
  XNOR2X1 U19712 ( .A(n6332), .B(top_core_KE_n1925), .Y(top_core_KE_n2006) );
  XNOR2X1 U19713 ( .A(n6319), .B(top_core_KE_n1957), .Y(top_core_KE_n2054) );
  XNOR2X1 U19714 ( .A(n6323), .B(top_core_KE_n1941), .Y(top_core_KE_n2030) );
  XNOR2X1 U19715 ( .A(n6692), .B(top_core_KE_n1923), .Y(top_core_KE_n2003) );
  XNOR2X1 U19716 ( .A(n6671), .B(top_core_KE_n1919), .Y(top_core_KE_n1995) );
  XNOR2X1 U19717 ( .A(n6647), .B(top_core_KE_n1917), .Y(top_core_KE_n1991) );
  XNOR2X1 U19718 ( .A(n6583), .B(top_core_KE_n1915), .Y(top_core_KE_n1987) );
  XNOR2X1 U19719 ( .A(n6513), .B(top_core_KE_n1913), .Y(top_core_KE_n1983) );
  XNOR2X1 U19720 ( .A(n6405), .B(top_core_KE_n1911), .Y(top_core_KE_n1979) );
  XNOR2X1 U19721 ( .A(n6310), .B(top_core_KE_n1921), .Y(top_core_KE_n1999) );
  NOR2X1 U19722 ( .A(n1679), .B(n1367), .Y(n13395) );
  NOR2X1 U19723 ( .A(n1734), .B(n1353), .Y(n12765) );
  NOR2X1 U19724 ( .A(n1705), .B(n1351), .Y(n13080) );
  NOR2X1 U19725 ( .A(n1643), .B(n1365), .Y(n13710) );
  NOR2X1 U19726 ( .A(n1171), .B(n1364), .Y(n12450) );
  NOR2X1 U19727 ( .A(n1211), .B(n1350), .Y(n11819) );
  NOR2X1 U19728 ( .A(n1210), .B(n1352), .Y(top_core_KE_sb1_n247) );
  NOR2X1 U19729 ( .A(n1170), .B(n1366), .Y(n12135) );
  AOI22X1 U19730 ( .A0(top_core_KE_n1865), .A1(top_core_KE_n897), .B0(
        top_core_KE_n896), .B1(top_core_KE_n1866), .Y(top_core_KE_n915) );
  NOR2X1 U19731 ( .A(n667), .B(n1358), .Y(n12340) );
  NOR2X1 U19732 ( .A(n665), .B(n1344), .Y(n11709) );
  NOR2X1 U19733 ( .A(n666), .B(n1345), .Y(top_core_KE_sb1_n134) );
  NOR2X1 U19734 ( .A(n668), .B(n1359), .Y(n12025) );
  AOI22X1 U19735 ( .A0(n1802), .A1(n1344), .B0(n1211), .B1(n625), .Y(n11736)
         );
  AOI22X1 U19736 ( .A0(n1823), .A1(n1345), .B0(n1210), .B1(n626), .Y(
        top_core_KE_sb1_n163) );
  AOI22X1 U19737 ( .A0(n1760), .A1(n1358), .B0(n1171), .B1(n627), .Y(n12367)
         );
  AOI22X1 U19738 ( .A0(n1781), .A1(n1359), .B0(n1170), .B1(n628), .Y(n12052)
         );
  AOI22X1 U19739 ( .A0(n1651), .A1(top_core_KE_prev_key1_reg_90_), .B0(n1643), 
        .B1(n631), .Y(n13628) );
  XNOR2X1 U19740 ( .A(n6962), .B(top_core_KE_new_sboxw_2_), .Y(
        top_core_KE_n1060) );
  XNOR2X1 U19741 ( .A(n6821), .B(top_core_KE_new_sboxw_5_), .Y(
        top_core_KE_n1039) );
  XNOR2X1 U19742 ( .A(n6668), .B(top_core_KE_new_sboxw_10_), .Y(
        top_core_KE_n1004) );
  XNOR2X1 U19743 ( .A(n6481), .B(top_core_KE_new_sboxw_13_), .Y(
        top_core_KE_n983) );
  XNOR2X1 U19744 ( .A(n6395), .B(top_core_KE_new_sboxw_15_), .Y(
        top_core_KE_n969) );
  XNOR2X1 U19745 ( .A(n6330), .B(top_core_KE_new_sboxw_7_), .Y(
        top_core_KE_n1025) );
  XNOR2X1 U19746 ( .A(n6956), .B(top_core_KE_new_sboxw_26_), .Y(
        top_core_KE_n1116) );
  XNOR2X1 U19747 ( .A(n6783), .B(top_core_KE_new_sboxw_29_), .Y(
        top_core_KE_n1095) );
  XNOR2X1 U19748 ( .A(n6379), .B(top_core_KE_new_sboxw_31_), .Y(
        top_core_KE_n1081) );
  XNOR2X1 U19749 ( .A(n6983), .B(top_core_KE_new_sboxw_0_), .Y(
        top_core_KE_n1074) );
  XNOR2X1 U19750 ( .A(n6978), .B(top_core_KE_new_sboxw_24_), .Y(
        top_core_KE_n1130) );
  XNOR2X1 U19751 ( .A(n6719), .B(top_core_KE_new_sboxw_6_), .Y(
        top_core_KE_n1032) );
  XNOR2X1 U19752 ( .A(n6690), .B(top_core_KE_new_sboxw_8_), .Y(
        top_core_KE_n1018) );
  XNOR2X1 U19753 ( .A(n6403), .B(top_core_KE_new_sboxw_14_), .Y(
        top_core_KE_n976) );
  XNOR2X1 U19754 ( .A(n6386), .B(top_core_KE_new_sboxw_30_), .Y(
        top_core_KE_n1088) );
  XNOR2X1 U19755 ( .A(n6973), .B(top_core_KE_new_sboxw_1_), .Y(
        top_core_KE_n1067) );
  XNOR2X1 U19756 ( .A(n6968), .B(top_core_KE_new_sboxw_25_), .Y(
        top_core_KE_n1123) );
  XNOR2X1 U19757 ( .A(n6946), .B(top_core_KE_new_sboxw_3_), .Y(
        top_core_KE_n1053) );
  XNOR2X1 U19758 ( .A(n6683), .B(top_core_KE_new_sboxw_9_), .Y(
        top_core_KE_n1011) );
  XNOR2X1 U19759 ( .A(n6931), .B(top_core_KE_new_sboxw_27_), .Y(
        top_core_KE_n1109) );
  XNOR2X1 U19760 ( .A(n6901), .B(top_core_KE_new_sboxw_4_), .Y(
        top_core_KE_n1046) );
  XNOR2X1 U19761 ( .A(n6855), .B(top_core_KE_new_sboxw_28_), .Y(
        top_core_KE_n1102) );
  XNOR2X1 U19762 ( .A(n6640), .B(top_core_KE_new_sboxw_11_), .Y(
        top_core_KE_n997) );
  XNOR2X1 U19763 ( .A(n6561), .B(top_core_KE_new_sboxw_12_), .Y(
        top_core_KE_n990) );
  XOR2X1 U19764 ( .A(top_core_KE_new_sboxw_21_), .B(n7000), .Y(
        top_core_KE_n2517) );
  XOR2X1 U19765 ( .A(top_core_KE_new_sboxw_18_), .B(n7003), .Y(
        top_core_KE_n2526) );
  OAI222XL U19766 ( .A0(top_core_EC_n1011), .A1(n4196), .B0(top_core_EC_n1017), 
        .B1(top_core_EC_n1013), .C0(n3986), .C1(n1), .Y(top_core_EC_n1292) );
  NOR2X1 U19767 ( .A(top_core_EC_n1018), .B(top_core_EC_n1019), .Y(
        top_core_EC_n1017) );
  AOI2BB1X1 U19768 ( .A0N(top_core_EC_n1022), .A1N(top_core_EC_n1014), .B0(
        n3976), .Y(top_core_EC_n1018) );
  AOI21X1 U19769 ( .A0(top_core_EC_n1020), .A1(n6307), .B0(n3985), .Y(
        top_core_EC_n1019) );
  OAI222XL U19770 ( .A0(top_core_EC_n1011), .A1(n4197), .B0(top_core_EC_n1012), 
        .B1(top_core_EC_n1013), .C0(n3975), .C1(n1), .Y(top_core_EC_n1291) );
  AOI32X1 U19771 ( .A0(n3984), .A1(n3975), .A2(top_core_EC_n1014), .B0(
        top_core_Addr[3]), .B1(top_core_EC_n1015), .Y(top_core_EC_n1012) );
  XOR2X1 U19772 ( .A(top_core_KE_new_sboxw_22_), .B(n6999), .Y(
        top_core_KE_n2514) );
  XOR2X1 U19773 ( .A(top_core_KE_new_sboxw_16_), .B(n7005), .Y(
        top_core_KE_n2532) );
  XOR2X1 U19774 ( .A(top_core_KE_new_sboxw_17_), .B(n7004), .Y(
        top_core_KE_n2529) );
  XOR2X1 U19775 ( .A(top_core_KE_new_sboxw_20_), .B(n7001), .Y(
        top_core_KE_n2520) );
  XOR2X1 U19776 ( .A(top_core_KE_new_sboxw_19_), .B(n7002), .Y(
        top_core_KE_n2523) );
  NOR2X1 U19777 ( .A(n11849), .B(n1350), .Y(n11701) );
  NOR2X1 U19778 ( .A(top_core_KE_sb1_n278), .B(n1352), .Y(top_core_KE_sb1_n126) );
  NOR2X1 U19779 ( .A(n12480), .B(n1364), .Y(n12332) );
  NOR2X1 U19780 ( .A(n13425), .B(n1367), .Y(n13278) );
  NOR2X1 U19781 ( .A(n12165), .B(n1366), .Y(n12017) );
  NOR2X1 U19782 ( .A(n12795), .B(n1353), .Y(n12648) );
  NOR2X1 U19783 ( .A(n13740), .B(n1365), .Y(n13593) );
  NOR2X1 U19784 ( .A(n13110), .B(n1351), .Y(n12963) );
  NAND2X1 U19785 ( .A(n1356), .B(n1340), .Y(n13207) );
  NAND2X1 U19786 ( .A(n1355), .B(n1337), .Y(n12892) );
  NAND2X1 U19787 ( .A(n1342), .B(n1336), .Y(n12577) );
  NAND2X1 U19788 ( .A(n1369), .B(n1341), .Y(n13522) );
  NAND2X1 U19789 ( .A(n1368), .B(n1370), .Y(n12262) );
  NAND2X1 U19790 ( .A(n1354), .B(n1338), .Y(n11630) );
  NAND2X1 U19791 ( .A(n1343), .B(n1335), .Y(top_core_KE_sb1_n55) );
  NAND2X1 U19792 ( .A(n1357), .B(n1339), .Y(n11946) );
  NAND2X1 U19793 ( .A(n1369), .B(n1635), .Y(n13532) );
  NAND2X1 U19794 ( .A(n1354), .B(n1795), .Y(n11640) );
  NAND2X1 U19795 ( .A(n1343), .B(n1816), .Y(top_core_KE_sb1_n65) );
  NAND2X1 U19796 ( .A(n1368), .B(n1752), .Y(n12272) );
  NAND2X1 U19797 ( .A(n1357), .B(n1774), .Y(n11956) );
  NAND2X1 U19798 ( .A(n1356), .B(n1668), .Y(n13217) );
  NAND2X1 U19799 ( .A(n1342), .B(n1726), .Y(n12587) );
  NAND2X1 U19800 ( .A(n1355), .B(n1697), .Y(n12902) );
  OAI211X1 U19801 ( .A0(n1813), .A1(n11919), .B0(n11925), .C0(n11926), .Y(
        n11917) );
  AOI222X1 U19802 ( .A0(n1800), .A1(n11927), .B0(n11928), .B1(n1796), .C0(
        n6824), .C1(n1808), .Y(n11926) );
  AOI31X1 U19803 ( .A0(n1223), .A1(n1350), .A2(n11652), .B0(n6827), .Y(n11925)
         );
  NAND4X1 U19804 ( .A(n11757), .B(n11716), .C(n11930), .D(n11931), .Y(n11927)
         );
  OAI211X1 U19805 ( .A0(n1834), .A1(top_core_KE_sb1_n348), .B0(
        top_core_KE_sb1_n354), .C0(top_core_KE_sb1_n355), .Y(
        top_core_KE_sb1_n346) );
  AOI222X1 U19806 ( .A0(n1821), .A1(top_core_KE_sb1_n356), .B0(
        top_core_KE_sb1_n357), .B1(n1817), .C0(n6802), .C1(n1829), .Y(
        top_core_KE_sb1_n355) );
  AOI31X1 U19807 ( .A0(n1217), .A1(n1352), .A2(top_core_KE_sb1_n77), .B0(n6805), .Y(top_core_KE_sb1_n354) );
  NAND4X1 U19808 ( .A(top_core_KE_sb1_n185), .B(top_core_KE_sb1_n143), .C(
        top_core_KE_sb1_n359), .D(top_core_KE_sb1_n360), .Y(
        top_core_KE_sb1_n356) );
  OAI211X1 U19809 ( .A0(n1773), .A1(n12550), .B0(n12556), .C0(n12557), .Y(
        n12548) );
  AOI222X1 U19810 ( .A0(n1758), .A1(n12558), .B0(n12559), .B1(n1753), .C0(
        n6528), .C1(n1763), .Y(n12557) );
  AOI31X1 U19811 ( .A0(n1182), .A1(n1364), .A2(n12284), .B0(n6531), .Y(n12556)
         );
  NAND4X1 U19812 ( .A(n12388), .B(n12347), .C(n12561), .D(n12562), .Y(n12558)
         );
  OAI211X1 U19813 ( .A0(n1691), .A1(n13495), .B0(n13501), .C0(n13502), .Y(
        n13493) );
  AOI222X1 U19814 ( .A0(n1667), .A1(n13503), .B0(n13504), .B1(n1672), .C0(
        n6470), .C1(n1686), .Y(n13502) );
  AOI31X1 U19815 ( .A0(n602), .A1(n1367), .A2(n13229), .B0(n6473), .Y(n13501)
         );
  NAND4X1 U19816 ( .A(n13334), .B(n13293), .C(n13506), .D(n13507), .Y(n13503)
         );
  OAI211X1 U19817 ( .A0(n1792), .A1(n12235), .B0(n12241), .C0(n12242), .Y(
        n12233) );
  AOI222X1 U19818 ( .A0(n1779), .A1(n12243), .B0(n12244), .B1(n1775), .C0(
        n6505), .C1(n1787), .Y(n12242) );
  AOI31X1 U19819 ( .A0(n1177), .A1(n1366), .A2(n11968), .B0(n6508), .Y(n12241)
         );
  NAND4X1 U19820 ( .A(n12073), .B(n12032), .C(n12246), .D(n12247), .Y(n12243)
         );
  OAI211X1 U19821 ( .A0(n1749), .A1(n12865), .B0(n12871), .C0(n12872), .Y(
        n12863) );
  AOI222X1 U19822 ( .A0(n1725), .A1(n12873), .B0(n12874), .B1(n1730), .C0(
        n6773), .C1(n1744), .Y(n12872) );
  AOI31X1 U19823 ( .A0(n603), .A1(n1353), .A2(n12599), .B0(n6776), .Y(n12871)
         );
  NAND4X1 U19824 ( .A(n12704), .B(n12663), .C(n12876), .D(n12877), .Y(n12873)
         );
  OAI211X1 U19825 ( .A0(n1663), .A1(n13810), .B0(n13816), .C0(n13817), .Y(
        n13808) );
  AOI222X1 U19826 ( .A0(n1641), .A1(n13818), .B0(n13819), .B1(n1636), .C0(
        n6517), .C1(n1653), .Y(n13817) );
  AOI31X1 U19827 ( .A0(n609), .A1(n1365), .A2(n13544), .B0(n6520), .Y(n13816)
         );
  NAND4X1 U19828 ( .A(n13649), .B(n13608), .C(n13821), .D(n13822), .Y(n13818)
         );
  OAI211X1 U19829 ( .A0(n1720), .A1(n13180), .B0(n13186), .C0(n13187), .Y(
        n13178) );
  AOI222X1 U19830 ( .A0(n1696), .A1(n13188), .B0(n13189), .B1(n1701), .C0(
        n6813), .C1(n1715), .Y(n13187) );
  AOI31X1 U19831 ( .A0(n604), .A1(n1351), .A2(n12914), .B0(n6816), .Y(n13186)
         );
  NAND4X1 U19832 ( .A(n13019), .B(n12978), .C(n13191), .D(n13192), .Y(n13188)
         );
  NAND2X1 U19833 ( .A(n1341), .B(n1146), .Y(n13524) );
  NAND2X1 U19834 ( .A(n1338), .B(n1187), .Y(n11632) );
  NAND2X1 U19835 ( .A(n1335), .B(n1224), .Y(top_core_KE_sb1_n57) );
  NAND2X1 U19836 ( .A(n1340), .B(n1185), .Y(n13209) );
  NAND2X1 U19837 ( .A(n1339), .B(n1184), .Y(n11948) );
  NAND2X1 U19838 ( .A(n1337), .B(n1186), .Y(n12894) );
  NAND2X1 U19839 ( .A(n1336), .B(n1225), .Y(n12579) );
  NAND2X1 U19840 ( .A(n1370), .B(n1147), .Y(n12264) );
  OAI221XL U19841 ( .A0(n1500), .A1(n6999), .B0(n7006), .B1(n151), .C0(
        top_core_KE_n2710), .Y(top_core_KE_n4928) );
  OAI221XL U19842 ( .A0(n1500), .A1(n7006), .B0(n7005), .B1(n151), .C0(
        top_core_KE_n2710), .Y(top_core_KE_n4927) );
  OAI221XL U19843 ( .A0(n1500), .A1(n7004), .B0(n7003), .B1(n151), .C0(
        top_core_KE_n2710), .Y(top_core_KE_n4925) );
  OAI221XL U19844 ( .A0(n686), .A1(n1150), .B0(n1367), .B1(n1688), .C0(n1363), 
        .Y(n13327) );
  OAI221XL U19845 ( .A0(n671), .A1(n1190), .B0(n1353), .B1(n1746), .C0(n1349), 
        .Y(n12697) );
  OAI221XL U19846 ( .A0(n672), .A1(n1199), .B0(n1351), .B1(n1717), .C0(n1347), 
        .Y(n13012) );
  OAI221XL U19847 ( .A0(n669), .A1(n1159), .B0(n1365), .B1(n1659), .C0(n1361), 
        .Y(n13642) );
  OAI221XL U19848 ( .A0(n683), .A1(n1164), .B0(n1364), .B1(n1768), .C0(n1360), 
        .Y(n12381) );
  OAI221XL U19849 ( .A0(n681), .A1(n1204), .B0(n1350), .B1(n1810), .C0(n1346), 
        .Y(n11750) );
  OAI221XL U19850 ( .A0(n682), .A1(n1195), .B0(n1352), .B1(n1831), .C0(n1348), 
        .Y(top_core_KE_sb1_n178) );
  OAI221XL U19851 ( .A0(n684), .A1(n1155), .B0(n1366), .B1(n1789), .C0(n1362), 
        .Y(n12066) );
  AOI21X1 U19852 ( .A0(n6904), .A1(n625), .B0(n11805), .Y(n11804) );
  AOI21X1 U19853 ( .A0(n6858), .A1(n626), .B0(top_core_KE_sb1_n233), .Y(
        top_core_KE_sb1_n232) );
  AOI21X1 U19854 ( .A0(n6611), .A1(n627), .B0(n12436), .Y(n12435) );
  AOI21X1 U19855 ( .A0(n6564), .A1(n628), .B0(n12121), .Y(n12120) );
  NAND3X1 U19856 ( .A(top_core_KE_n2723), .B(top_core_KE_n2705), .C(
        top_core_KE_n2724), .Y(top_core_KE_n2721) );
  NAND3X1 U19857 ( .A(top_core_KE_n875), .B(top_core_KE_round_ctr_reg_0_), .C(
        n1333), .Y(top_core_KE_n881) );
  NAND3X1 U19858 ( .A(top_core_KE_n878), .B(top_core_KE_round_ctr_reg_0_), .C(
        n1334), .Y(top_core_KE_n890) );
  AOI31X1 U19859 ( .A0(n11824), .A1(n11825), .A2(n11826), .B0(n11632), .Y(
        n11823) );
  AOI211X1 U19860 ( .A0(n11827), .A1(n1222), .B0(n11828), .C0(n11829), .Y(
        n11826) );
  AOI31X1 U19861 ( .A0(n1810), .A1(n1350), .A2(n11652), .B0(n11833), .Y(n11824) );
  AOI31X1 U19862 ( .A0(top_core_KE_sb1_n253), .A1(top_core_KE_sb1_n254), .A2(
        top_core_KE_sb1_n255), .B0(top_core_KE_sb1_n57), .Y(
        top_core_KE_sb1_n252) );
  AOI211X1 U19863 ( .A0(top_core_KE_sb1_n256), .A1(n1216), .B0(
        top_core_KE_sb1_n257), .C0(top_core_KE_sb1_n258), .Y(
        top_core_KE_sb1_n255) );
  AOI31X1 U19864 ( .A0(n1831), .A1(n1352), .A2(top_core_KE_sb1_n77), .B0(
        top_core_KE_sb1_n262), .Y(top_core_KE_sb1_n253) );
  AOI31X1 U19865 ( .A0(n12455), .A1(n12456), .A2(n12457), .B0(n12264), .Y(
        n12454) );
  AOI211X1 U19866 ( .A0(n12458), .A1(n1181), .B0(n12459), .C0(n12460), .Y(
        n12457) );
  AOI31X1 U19867 ( .A0(n1768), .A1(n1364), .A2(n12284), .B0(n12464), .Y(n12455) );
  AOI31X1 U19868 ( .A0(n13400), .A1(n13401), .A2(n13402), .B0(n13209), .Y(
        n13399) );
  AOI211X1 U19869 ( .A0(n13403), .A1(n1173), .B0(n13404), .C0(n13405), .Y(
        n13402) );
  AOI31X1 U19870 ( .A0(n1688), .A1(n1367), .A2(n13229), .B0(n13409), .Y(n13400) );
  AOI31X1 U19871 ( .A0(n12140), .A1(n12141), .A2(n12142), .B0(n11948), .Y(
        n12139) );
  AOI211X1 U19872 ( .A0(n12143), .A1(n1176), .B0(n12144), .C0(n12145), .Y(
        n12142) );
  AOI31X1 U19873 ( .A0(n1789), .A1(n1366), .A2(n11968), .B0(n12149), .Y(n12140) );
  AOI31X1 U19874 ( .A0(n12770), .A1(n12771), .A2(n12772), .B0(n12579), .Y(
        n12769) );
  AOI211X1 U19875 ( .A0(n12773), .A1(n1213), .B0(n12774), .C0(n12775), .Y(
        n12772) );
  AOI31X1 U19876 ( .A0(n1746), .A1(n1353), .A2(n12599), .B0(n12779), .Y(n12770) );
  AOI31X1 U19877 ( .A0(n13715), .A1(n13716), .A2(n13717), .B0(n13524), .Y(
        n13714) );
  AOI211X1 U19878 ( .A0(n13718), .A1(n1178), .B0(n13719), .C0(n13720), .Y(
        n13717) );
  AOI31X1 U19879 ( .A0(n1659), .A1(n1365), .A2(n13544), .B0(n13724), .Y(n13715) );
  AOI31X1 U19880 ( .A0(n13085), .A1(n13086), .A2(n13087), .B0(n12894), .Y(
        n13084) );
  AOI211X1 U19881 ( .A0(n13088), .A1(n1219), .B0(n13089), .C0(n13090), .Y(
        n13087) );
  AOI31X1 U19882 ( .A0(n1717), .A1(n1351), .A2(n12914), .B0(n13094), .Y(n13085) );
  INVX1 U19883 ( .A(n11772), .Y(n6910) );
  INVX1 U19884 ( .A(top_core_KE_sb1_n200), .Y(n6864) );
  INVX1 U19885 ( .A(n12403), .Y(n6617) );
  INVX1 U19886 ( .A(n13349), .Y(n6545) );
  INVX1 U19887 ( .A(n12088), .Y(n6570) );
  INVX1 U19888 ( .A(n12719), .Y(n6840) );
  INVX1 U19889 ( .A(n13664), .Y(n6593) );
  INVX1 U19890 ( .A(n13034), .Y(n6886) );
  NAND2X1 U19891 ( .A(n2141), .B(top_core_KE_n894), .Y(top_core_KE_n2509) );
  NAND2X1 U19892 ( .A(top_core_KE_round_ctr_reg_0_), .B(top_core_KE_n2705), 
        .Y(top_core_KE_n2716) );
  NOR2X1 U19893 ( .A(n6308), .B(n3541), .Y(top_core_EC_n862) );
  NOR2X1 U19894 ( .A(n3561), .B(n6308), .Y(top_core_EC_n943) );
  OAI21XL U19895 ( .A0(top_core_KE_round_ctr_reg_0_), .A1(n7016), .B0(
        top_core_KE_n2719), .Y(top_core_KE_n2718) );
  NAND2X1 U19896 ( .A(n1356), .B(n1666), .Y(n13307) );
  NAND2X1 U19897 ( .A(n1355), .B(n1695), .Y(n12992) );
  NAND2X1 U19898 ( .A(n1342), .B(n1724), .Y(n12677) );
  NAND2X1 U19899 ( .A(n1673), .B(n1367), .Y(n13310) );
  NAND2X1 U19900 ( .A(n1731), .B(n1353), .Y(n12680) );
  NAND2X1 U19901 ( .A(n1702), .B(n1351), .Y(n12995) );
  NAND2X1 U19902 ( .A(n1646), .B(n1365), .Y(n13625) );
  NAND2X1 U19903 ( .A(n1358), .B(n1364), .Y(n12364) );
  NAND2X1 U19904 ( .A(n1344), .B(n1350), .Y(n11733) );
  NAND2X1 U19905 ( .A(n1345), .B(n1352), .Y(top_core_KE_sb1_n160) );
  NAND2X1 U19906 ( .A(n1359), .B(n1366), .Y(n12049) );
  NAND2X1 U19907 ( .A(n1354), .B(n1798), .Y(n11730) );
  NAND2X1 U19908 ( .A(n1343), .B(n1819), .Y(top_core_KE_sb1_n157) );
  NAND2X1 U19909 ( .A(n1368), .B(n1755), .Y(n12361) );
  NAND2X1 U19910 ( .A(n1357), .B(n1777), .Y(n12046) );
  NAND2X1 U19911 ( .A(n1369), .B(n1637), .Y(n13622) );
  AOI21X1 U19912 ( .A0(n7014), .A1(top_core_KE_n2705), .B0(top_core_KE_n2718), 
        .Y(top_core_KE_n2717) );
  OAI211X1 U19913 ( .A0(top_core_KE_n2725), .A1(n7017), .B0(top_core_KE_n2720), 
        .C0(top_core_KE_n2721), .Y(top_core_KE_n4932) );
  NAND2X1 U19914 ( .A(n3569), .B(n6308), .Y(top_core_EC_n947) );
  NAND2X1 U19915 ( .A(n1174), .B(n1363), .Y(n13319) );
  NAND2X1 U19916 ( .A(n1214), .B(n1349), .Y(n12689) );
  NAND2X1 U19917 ( .A(n1220), .B(n1347), .Y(n13004) );
  NAND2X1 U19918 ( .A(n1179), .B(n1361), .Y(n13634) );
  NAND2X1 U19919 ( .A(n607), .B(n1360), .Y(n12373) );
  NAND2X1 U19920 ( .A(n605), .B(n1346), .Y(n11742) );
  NAND2X1 U19921 ( .A(n606), .B(n1348), .Y(top_core_KE_sb1_n169) );
  NAND2X1 U19922 ( .A(n608), .B(n1362), .Y(n12058) );
  NAND2XL U19923 ( .A(top_core_KE_n2705), .B(top_core_KE_n1865), .Y(
        top_core_KE_n743) );
  AOI211X1 U19924 ( .A0(n11652), .A1(n11739), .B0(n11740), .C0(n11741), .Y(
        n11738) );
  AOI22X1 U19925 ( .A0(n1798), .A1(n11743), .B0(n11744), .B1(n1795), .Y(n11737) );
  OAI21XL U19926 ( .A0(n1350), .A1(n665), .B0(n1346), .Y(n11739) );
  AOI211X1 U19927 ( .A0(top_core_KE_sb1_n77), .A1(top_core_KE_sb1_n166), .B0(
        top_core_KE_sb1_n167), .C0(top_core_KE_sb1_n168), .Y(
        top_core_KE_sb1_n165) );
  AOI22X1 U19928 ( .A0(n1819), .A1(top_core_KE_sb1_n170), .B0(
        top_core_KE_sb1_n171), .B1(n1816), .Y(top_core_KE_sb1_n164) );
  OAI21XL U19929 ( .A0(n1352), .A1(n666), .B0(n1348), .Y(top_core_KE_sb1_n166)
         );
  AOI211X1 U19930 ( .A0(n12284), .A1(n12370), .B0(n12371), .C0(n12372), .Y(
        n12369) );
  AOI22X1 U19931 ( .A0(top_core_KE_prev_key1_reg_29_), .A1(n12374), .B0(n12375), .B1(n1752), .Y(n12368) );
  OAI21XL U19932 ( .A0(n1364), .A1(n667), .B0(n1360), .Y(n12370) );
  AOI211X1 U19933 ( .A0(n13229), .A1(n13316), .B0(n13317), .C0(n13318), .Y(
        n13315) );
  AOI22X1 U19934 ( .A0(n1666), .A1(n13320), .B0(n13321), .B1(n1668), .Y(n13314) );
  OAI21XL U19935 ( .A0(n1367), .A1(n670), .B0(n1363), .Y(n13316) );
  AOI211X1 U19936 ( .A0(n11968), .A1(n12055), .B0(n12056), .C0(n12057), .Y(
        n12054) );
  AOI22X1 U19937 ( .A0(n1777), .A1(n12059), .B0(n12060), .B1(n1774), .Y(n12053) );
  OAI21XL U19938 ( .A0(n1366), .A1(n668), .B0(n1362), .Y(n12055) );
  AOI211X1 U19939 ( .A0(n12599), .A1(n12686), .B0(n12687), .C0(n12688), .Y(
        n12685) );
  AOI22X1 U19940 ( .A0(n1724), .A1(n12690), .B0(n12691), .B1(n1726), .Y(n12684) );
  OAI21XL U19941 ( .A0(n1353), .A1(n671), .B0(n1349), .Y(n12686) );
  AOI211X1 U19942 ( .A0(n12914), .A1(n13001), .B0(n13002), .C0(n13003), .Y(
        n13000) );
  AOI22X1 U19943 ( .A0(n1695), .A1(n13005), .B0(n13006), .B1(n1697), .Y(n12999) );
  OAI21XL U19944 ( .A0(n1351), .A1(n672), .B0(n1347), .Y(n13001) );
  AOI211X1 U19945 ( .A0(n13544), .A1(n13631), .B0(n13632), .C0(n13633), .Y(
        n13630) );
  AOI22X1 U19946 ( .A0(top_core_KE_prev_key1_reg_93_), .A1(n13635), .B0(n13636), .B1(n1635), .Y(n13629) );
  OAI21XL U19947 ( .A0(n1365), .A1(n669), .B0(n1361), .Y(n13631) );
  CLKINVX3 U19948 ( .A(n1341), .Y(n6989) );
  AOI21X1 U19949 ( .A0(n11673), .A1(n11773), .B0(n11674), .Y(n11781) );
  AOI21X1 U19950 ( .A0(top_core_KE_sb1_n98), .A1(top_core_KE_sb1_n201), .B0(
        top_core_KE_sb1_n99), .Y(top_core_KE_sb1_n209) );
  AOI21X1 U19951 ( .A0(n12304), .A1(n12404), .B0(n12305), .Y(n12412) );
  AOI21X1 U19952 ( .A0(n11989), .A1(n12089), .B0(n11990), .Y(n12097) );
  AOI21X1 U19953 ( .A0(n12620), .A1(n12720), .B0(n12621), .Y(n12727) );
  AOI21X1 U19954 ( .A0(n13565), .A1(n13665), .B0(n13566), .Y(n13672) );
  AOI21X1 U19955 ( .A0(n12935), .A1(n13035), .B0(n12936), .Y(n13042) );
  NAND2X1 U19956 ( .A(top_core_KE_n1864), .B(top_core_KE_round_ctr_reg_0_), 
        .Y(top_core_KE_n914) );
  NAND3X1 U19957 ( .A(top_core_KE_round_ctr_reg_0_), .B(n1226), .C(
        top_core_KE_n875), .Y(top_core_KE_n876) );
  NAND3X1 U19958 ( .A(top_core_KE_round_ctr_reg_0_), .B(n7007), .C(
        top_core_KE_n878), .Y(top_core_KE_n879) );
  NOR4BBX1 U19959 ( .AN(n13351), .BN(n13352), .C(n13230), .D(n13219), .Y(
        n13322) );
  AOI222X1 U19960 ( .A0(n1667), .A1(n13353), .B0(n13354), .B1(n1669), .C0(n602), .C1(n6470), .Y(n13352) );
  OAI21XL U19961 ( .A0(n13355), .A1(n1274), .B0(n13267), .Y(n13354) );
  CLKINVX3 U19962 ( .A(n1336), .Y(n6995) );
  CLKINVX3 U19963 ( .A(n1337), .Y(n6994) );
  CLKINVX3 U19964 ( .A(n1340), .Y(n6990) );
  CLKINVX3 U19965 ( .A(n1339), .Y(n6992) );
  CLKINVX3 U19966 ( .A(n1338), .Y(n6993) );
  CLKINVX3 U19967 ( .A(n1335), .Y(n6997) );
  MX2X1 U19968 ( .A(n1333), .B(n1226), .S0(top_core_KE_r343_quotient_2_), .Y(
        top_core_KE_r343_u_div_PartRem_2__1_) );
  MX2X1 U19969 ( .A(n1332), .B(n7014), .S0(n7010), .Y(
        top_core_KE_r343_u_div_PartRem_1__1_) );
  AOI31X1 U19970 ( .A0(n13220), .A1(n13221), .A2(n13222), .B0(n1356), .Y(
        n13212) );
  AOI2BB2X1 U19971 ( .B0(n13231), .B1(n756), .A0N(n13232), .A1N(n610), .Y(
        n13220) );
  AOI31X1 U19972 ( .A0(n12905), .A1(n12906), .A2(n12907), .B0(n1355), .Y(
        n12897) );
  AOI2BB2X1 U19973 ( .B0(n12916), .B1(n758), .A0N(n12917), .A1N(n612), .Y(
        n12905) );
  AOI31X1 U19974 ( .A0(n12590), .A1(n12591), .A2(n12592), .B0(n1342), .Y(
        n12582) );
  AOI2BB2X1 U19975 ( .B0(n12601), .B1(n757), .A0N(n12602), .A1N(n611), .Y(
        n12590) );
  AOI31X1 U19976 ( .A0(n13535), .A1(n13536), .A2(n13537), .B0(n1369), .Y(
        n13527) );
  AOI2BB2X1 U19977 ( .B0(n13546), .B1(n759), .A0N(n13547), .A1N(n616), .Y(
        n13535) );
  AOI31X1 U19978 ( .A0(n12275), .A1(n12276), .A2(n12277), .B0(n1368), .Y(
        n12267) );
  AOI2BB2X1 U19979 ( .B0(n12286), .B1(n760), .A0N(n12287), .A1N(n1182), .Y(
        n12275) );
  AOI31X1 U19980 ( .A0(n11643), .A1(n11644), .A2(n11645), .B0(n1354), .Y(
        n11635) );
  AOI2BB2X1 U19981 ( .B0(n11654), .B1(n761), .A0N(n11655), .A1N(n1223), .Y(
        n11643) );
  AOI31X1 U19982 ( .A0(top_core_KE_sb1_n68), .A1(top_core_KE_sb1_n69), .A2(
        top_core_KE_sb1_n70), .B0(n1343), .Y(top_core_KE_sb1_n60) );
  AOI2BB2X1 U19983 ( .B0(top_core_KE_sb1_n79), .B1(n762), .A0N(
        top_core_KE_sb1_n80), .A1N(n1217), .Y(top_core_KE_sb1_n68) );
  AOI31X1 U19984 ( .A0(n11959), .A1(n11960), .A2(n11961), .B0(n1357), .Y(
        n11951) );
  AOI2BB2X1 U19985 ( .B0(n11970), .B1(n763), .A0N(n11971), .A1N(n1177), .Y(
        n11959) );
  AOI31X1 U19986 ( .A0(n13214), .A1(n13215), .A2(n13216), .B0(n13217), .Y(
        n13213) );
  NAND3X1 U19987 ( .A(n1174), .B(n1674), .C(n717), .Y(n13215) );
  AOI22X1 U19988 ( .A0(n1687), .A1(n13218), .B0(n6544), .B1(n629), .Y(n13216)
         );
  AOI31X1 U19989 ( .A0(n1367), .A1(n6633), .A2(n1173), .B0(n13219), .Y(n13214)
         );
  AOI31X1 U19990 ( .A0(n12899), .A1(n12900), .A2(n12901), .B0(n12902), .Y(
        n12898) );
  NAND3X1 U19991 ( .A(n1220), .B(n1703), .C(n721), .Y(n12900) );
  AOI22X1 U19992 ( .A0(n1716), .A1(n12903), .B0(n6885), .B1(n632), .Y(n12901)
         );
  AOI31X1 U19993 ( .A0(n1351), .A1(n6940), .A2(n1219), .B0(n12904), .Y(n12899)
         );
  AOI31X1 U19994 ( .A0(n12269), .A1(n12270), .A2(n12271), .B0(n12272), .Y(
        n12268) );
  NAND3X1 U19995 ( .A(n607), .B(n1358), .C(n716), .Y(n12270) );
  AOI22X1 U19996 ( .A0(n1767), .A1(n12273), .B0(n6616), .B1(n627), .Y(n12271)
         );
  AOI31X1 U19997 ( .A0(n1364), .A1(n6658), .A2(n1181), .B0(n12274), .Y(n12269)
         );
  AOI31X1 U19998 ( .A0(n13529), .A1(n13530), .A2(n13531), .B0(n13532), .Y(
        n13528) );
  NAND3X1 U19999 ( .A(n1179), .B(n1649), .C(n720), .Y(n13530) );
  AOI22X1 U20000 ( .A0(n1658), .A1(n13533), .B0(n6592), .B1(n631), .Y(n13531)
         );
  AOI31X1 U20001 ( .A0(n1365), .A1(n6650), .A2(n1178), .B0(n13534), .Y(n13529)
         );
  AOI31X1 U20002 ( .A0(n12584), .A1(n12585), .A2(n12586), .B0(n12587), .Y(
        n12583) );
  NAND3X1 U20003 ( .A(n1214), .B(n1732), .C(n719), .Y(n12585) );
  AOI22X1 U20004 ( .A0(n1745), .A1(n12588), .B0(n6839), .B1(n630), .Y(n12586)
         );
  AOI31X1 U20005 ( .A0(n1353), .A1(n6925), .A2(n1213), .B0(n12589), .Y(n12584)
         );
  AOI31X1 U20006 ( .A0(n11637), .A1(n11638), .A2(n11639), .B0(n11640), .Y(
        n11636) );
  NAND3X1 U20007 ( .A(n605), .B(n1344), .C(n714), .Y(n11638) );
  AOI22X1 U20008 ( .A0(n1809), .A1(n11641), .B0(n6909), .B1(n625), .Y(n11639)
         );
  AOI31X1 U20009 ( .A0(n1350), .A1(n6948), .A2(n1222), .B0(n11642), .Y(n11637)
         );
  AOI31X1 U20010 ( .A0(top_core_KE_sb1_n62), .A1(top_core_KE_sb1_n63), .A2(
        top_core_KE_sb1_n64), .B0(top_core_KE_sb1_n65), .Y(top_core_KE_sb1_n61) );
  NAND3X1 U20011 ( .A(n606), .B(n1345), .C(n715), .Y(top_core_KE_sb1_n63) );
  AOI22X1 U20012 ( .A0(n1830), .A1(top_core_KE_sb1_n66), .B0(n6863), .B1(n626), 
        .Y(top_core_KE_sb1_n64) );
  AOI31X1 U20013 ( .A0(n1352), .A1(n6933), .A2(n1216), .B0(top_core_KE_sb1_n67), .Y(top_core_KE_sb1_n62) );
  AOI31X1 U20014 ( .A0(n11953), .A1(n11954), .A2(n11955), .B0(n11956), .Y(
        n11952) );
  NAND3X1 U20015 ( .A(n608), .B(n1359), .C(n718), .Y(n11954) );
  AOI22X1 U20016 ( .A0(n1788), .A1(n11957), .B0(n6569), .B1(n628), .Y(n11955)
         );
  AOI31X1 U20017 ( .A0(n1366), .A1(n6642), .A2(n1176), .B0(n11958), .Y(n11953)
         );
  NAND3X1 U20018 ( .A(n1367), .B(n1678), .C(n610), .Y(n13383) );
  NAND3X1 U20019 ( .A(n1350), .B(n1211), .C(n1223), .Y(n11807) );
  NAND3X1 U20020 ( .A(n1352), .B(n1210), .C(n1217), .Y(top_core_KE_sb1_n235)
         );
  NAND3X1 U20021 ( .A(n1364), .B(n1171), .C(n1182), .Y(n12438) );
  NAND3X1 U20022 ( .A(n1366), .B(n1170), .C(n1177), .Y(n12123) );
  NAND3X1 U20023 ( .A(n1353), .B(n1737), .C(n611), .Y(n12753) );
  NAND3X1 U20024 ( .A(n1365), .B(n1644), .C(n616), .Y(n13698) );
  NAND3X1 U20025 ( .A(n1351), .B(n1708), .C(n612), .Y(n13068) );
  NAND2X1 U20026 ( .A(top_core_EC_n943), .B(top_core_EC_n944), .Y(
        top_core_EC_n869) );
  CLKINVX3 U20027 ( .A(n1332), .Y(n7014) );
  NAND2X1 U20028 ( .A(top_core_KE_n1866), .B(top_core_KE_n2705), .Y(
        top_core_KE_n873) );
  AND2X2 U20029 ( .A(top_core_KE_n884), .B(n1332), .Y(top_core_KE_n887) );
  NAND3X1 U20030 ( .A(top_core_KE_round_ctr_reg_0_), .B(top_core_KE_n883), .C(
        top_core_KE_n884), .Y(top_core_KE_n885) );
  AND3X2 U20031 ( .A(top_core_KE_n2506), .B(top_core_KE_n894), .C(n2286), .Y(
        top_core_KE_n2176) );
  NAND3X1 U20032 ( .A(top_core_KE_round_ctr_reg_0_), .B(n1226), .C(
        top_core_KE_n887), .Y(top_core_KE_n888) );
  NOR2X1 U20033 ( .A(n1582), .B(n4262), .Y(top_core_io_n1179) );
  NOR2X1 U20034 ( .A(n1582), .B(n4261), .Y(top_core_io_n1180) );
  AND2X2 U20035 ( .A(top_core_EC_n1009), .B(top_core_EC_n944), .Y(
        top_core_EC_n950) );
  AND2X2 U20036 ( .A(top_core_EC_n1009), .B(n6306), .Y(top_core_EC_n951) );
  OAI22XL U20037 ( .A0(n1360), .A1(n627), .B0(n12367), .B1(n12349), .Y(n12375)
         );
  OAI22XL U20038 ( .A0(n1361), .A1(n631), .B0(n13628), .B1(n13610), .Y(n13636)
         );
  OAI22XL U20039 ( .A0(n1346), .A1(n625), .B0(n11736), .B1(n11718), .Y(n11744)
         );
  OAI22XL U20040 ( .A0(n1348), .A1(n626), .B0(top_core_KE_sb1_n163), .B1(
        top_core_KE_sb1_n145), .Y(top_core_KE_sb1_n171) );
  OAI22XL U20041 ( .A0(n1363), .A1(n629), .B0(n13313), .B1(n13295), .Y(n13321)
         );
  OAI22XL U20042 ( .A0(n1362), .A1(n628), .B0(n12052), .B1(n12034), .Y(n12060)
         );
  OAI22XL U20043 ( .A0(n1349), .A1(n630), .B0(n12683), .B1(n12665), .Y(n12691)
         );
  OAI22XL U20044 ( .A0(n1347), .A1(n632), .B0(n12998), .B1(n12980), .Y(n13006)
         );
  INVX1 U20045 ( .A(top_core_KE_Nk0_0_), .Y(n7019) );
  NAND2X1 U20046 ( .A(n7016), .B(top_core_KE_n2720), .Y(top_core_KE_n2719) );
  INVX1 U20047 ( .A(n1358), .Y(n6677) );
  XNOR2X1 U20048 ( .A(n6961), .B(top_core_KE_new_sboxw_2_), .Y(
        top_core_KE_n1058) );
  XNOR2X1 U20049 ( .A(n6820), .B(top_core_KE_new_sboxw_5_), .Y(
        top_core_KE_n1037) );
  XNOR2X1 U20050 ( .A(n6328), .B(top_core_KE_new_sboxw_7_), .Y(
        top_core_KE_n1023) );
  XNOR2X1 U20051 ( .A(n6955), .B(top_core_KE_new_sboxw_26_), .Y(
        top_core_KE_n1114) );
  XNOR2X1 U20052 ( .A(n6781), .B(top_core_KE_new_sboxw_29_), .Y(
        top_core_KE_n1093) );
  XNOR2X1 U20053 ( .A(n6377), .B(top_core_KE_new_sboxw_31_), .Y(
        top_core_KE_n1079) );
  XNOR2X1 U20054 ( .A(top_core_KE_n2147), .B(n6983), .Y(top_core_KE_n2298) );
  XNOR2X1 U20055 ( .A(top_core_KE_n2171), .B(n6978), .Y(top_core_KE_n2338) );
  XNOR2X1 U20056 ( .A(top_core_KE_n2144), .B(n6973), .Y(top_core_KE_n2293) );
  XNOR2X1 U20057 ( .A(top_core_KE_n2168), .B(n6968), .Y(top_core_KE_n2333) );
  XNOR2X1 U20058 ( .A(top_core_KE_n2141), .B(n6962), .Y(top_core_KE_n2288) );
  XNOR2X1 U20059 ( .A(top_core_KE_n2165), .B(n6956), .Y(top_core_KE_n2328) );
  XNOR2X1 U20060 ( .A(top_core_KE_n2138), .B(n6946), .Y(top_core_KE_n2283) );
  XNOR2X1 U20061 ( .A(top_core_KE_n2162), .B(n6931), .Y(top_core_KE_n2323) );
  XNOR2X1 U20062 ( .A(top_core_KE_n2135), .B(n6901), .Y(top_core_KE_n2278) );
  XNOR2X1 U20063 ( .A(top_core_KE_n2159), .B(n6855), .Y(top_core_KE_n2318) );
  XNOR2X1 U20064 ( .A(top_core_KE_n2132), .B(n6821), .Y(top_core_KE_n2273) );
  XNOR2X1 U20065 ( .A(top_core_KE_n2156), .B(n6783), .Y(top_core_KE_n2313) );
  XNOR2X1 U20066 ( .A(top_core_KE_n2129), .B(n6719), .Y(top_core_KE_n2268) );
  XNOR2X1 U20067 ( .A(top_core_KE_n2099), .B(n6696), .Y(top_core_KE_n2218) );
  XNOR2X1 U20068 ( .A(top_core_KE_n2123), .B(n6690), .Y(top_core_KE_n2258) );
  XNOR2X1 U20069 ( .A(top_core_KE_n2120), .B(n6683), .Y(top_core_KE_n2253) );
  XNOR2X1 U20070 ( .A(top_core_KE_n2093), .B(n6675), .Y(top_core_KE_n2208) );
  XNOR2X1 U20071 ( .A(top_core_KE_n2117), .B(n6668), .Y(top_core_KE_n2248) );
  XNOR2X1 U20072 ( .A(top_core_KE_n2090), .B(n6656), .Y(top_core_KE_n2203) );
  XNOR2X1 U20073 ( .A(top_core_KE_n2114), .B(n6640), .Y(top_core_KE_n2243) );
  XNOR2X1 U20074 ( .A(top_core_KE_n2087), .B(n6608), .Y(top_core_KE_n2198) );
  XNOR2X1 U20075 ( .A(top_core_KE_n2111), .B(n6561), .Y(top_core_KE_n2238) );
  XNOR2X1 U20076 ( .A(top_core_KE_n2084), .B(n6525), .Y(top_core_KE_n2193) );
  XNOR2X1 U20077 ( .A(top_core_KE_n2108), .B(n6481), .Y(top_core_KE_n2233) );
  XNOR2X1 U20078 ( .A(top_core_KE_n2081), .B(n6437), .Y(top_core_KE_n2188) );
  XNOR2X1 U20079 ( .A(top_core_KE_n2105), .B(n6403), .Y(top_core_KE_n2228) );
  XNOR2X1 U20080 ( .A(top_core_KE_n2102), .B(n6395), .Y(top_core_KE_n2223) );
  XNOR2X1 U20081 ( .A(top_core_KE_n2153), .B(n6386), .Y(top_core_KE_n2308) );
  XNOR2X1 U20082 ( .A(top_core_KE_n2150), .B(n6379), .Y(top_core_KE_n2303) );
  XNOR2X1 U20083 ( .A(top_core_KE_n2078), .B(n6344), .Y(top_core_KE_n2180) );
  XNOR2X1 U20084 ( .A(top_core_KE_n2126), .B(n6330), .Y(top_core_KE_n2263) );
  XNOR2X1 U20085 ( .A(top_core_KE_n2096), .B(n6317), .Y(top_core_KE_n2213) );
  XNOR2X1 U20086 ( .A(top_core_KE_new_sboxw_31_), .B(top_core_KE_n1909), .Y(
        top_core_KE_n1133) );
  XNOR2X1 U20087 ( .A(top_core_KE_new_sboxw_26_), .B(top_core_KE_n1919), .Y(
        top_core_KE_n1168) );
  XNOR2X1 U20088 ( .A(top_core_KE_new_sboxw_29_), .B(top_core_KE_n1913), .Y(
        top_core_KE_n1147) );
  INVX1 U20089 ( .A(top_core_KE_n1974), .Y(n6448) );
  INVX1 U20090 ( .A(top_core_KE_n2002), .Y(n6466) );
  INVX1 U20091 ( .A(top_core_KE_n1994), .Y(n6461) );
  INVX1 U20092 ( .A(top_core_KE_n1990), .Y(n6458) );
  INVX1 U20093 ( .A(top_core_KE_n1998), .Y(n6463) );
  INVX1 U20094 ( .A(top_core_KE_n1986), .Y(n6455) );
  INVX1 U20095 ( .A(top_core_KE_n1982), .Y(n6452) );
  INVX1 U20096 ( .A(top_core_KE_n1978), .Y(n6449) );
  XOR2X1 U20097 ( .A(top_core_Key[121]), .B(top_core_EC_add_in_r[1]), .Y(
        top_core_EC_add_out_r_1_) );
  OAI22X1 U20098 ( .A0(n3619), .A1(n6303), .B0(top_core_EC_ss_n218), .B1(n3606), .Y(top_core_EC_add_in_r[1]) );
  XOR2X1 U20099 ( .A(top_core_Key[106]), .B(top_core_EC_add_in_r[18]), .Y(
        top_core_EC_add_out_r_18_) );
  OAI22X1 U20100 ( .A0(n3618), .A1(n6286), .B0(top_core_EC_ss_n220), .B1(n3607), .Y(top_core_EC_add_in_r[18]) );
  XOR2X1 U20101 ( .A(top_core_Key[122]), .B(top_core_EC_add_in_r[2]), .Y(
        top_core_EC_add_out_r_2_) );
  OAI22X1 U20102 ( .A0(n3582), .A1(n6302), .B0(top_core_EC_ss_n207), .B1(n3598), .Y(top_core_EC_add_in_r[2]) );
  XOR2X1 U20103 ( .A(top_core_Key[90]), .B(top_core_EC_add_in_r[34]), .Y(
        top_core_EC_add_out_r_34_) );
  OAI22X1 U20104 ( .A0(n3582), .A1(n6270), .B0(top_core_EC_ss_n202), .B1(n3596), .Y(top_core_EC_add_in_r[34]) );
  XOR2X1 U20105 ( .A(top_core_Key[74]), .B(top_core_EC_add_in_r[50]), .Y(
        top_core_EC_add_out_r_50_) );
  OAI22X1 U20106 ( .A0(n3584), .A1(n6254), .B0(top_core_EC_ss_n184), .B1(n3596), .Y(top_core_EC_add_in_r[50]) );
  XOR2X1 U20107 ( .A(top_core_Key[104]), .B(top_core_EC_add_in_r[16]), .Y(
        top_core_EC_add_out_r_16_) );
  OAI22X1 U20108 ( .A0(n3582), .A1(n6288), .B0(top_core_EC_ss_n222), .B1(n3624), .Y(top_core_EC_add_in_r[16]) );
  XOR2X1 U20109 ( .A(top_core_Key[120]), .B(top_core_EC_add_in_r[0]), .Y(
        top_core_EC_add_out_r_0_) );
  OAI22X1 U20110 ( .A0(n3622), .A1(n6304), .B0(top_core_EC_ss_n257), .B1(n3608), .Y(top_core_EC_add_in_r[0]) );
  XOR2X1 U20111 ( .A(top_core_Key[107]), .B(top_core_EC_add_in_r[19]), .Y(
        top_core_EC_add_out_r_19_) );
  OAI22X1 U20112 ( .A0(n3614), .A1(n6285), .B0(top_core_EC_ss_n219), .B1(n3606), .Y(top_core_EC_add_in_r[19]) );
  XOR2X1 U20113 ( .A(top_core_Key[127]), .B(top_core_EC_add_in_r[7]), .Y(
        top_core_EC_add_out_r_7_) );
  OAI22X1 U20114 ( .A0(n3585), .A1(n6297), .B0(top_core_EC_ss_n152), .B1(n3589), .Y(top_core_EC_add_in_r[7]) );
  XOR2X1 U20115 ( .A(top_core_Key[123]), .B(top_core_EC_add_in_r[3]), .Y(
        top_core_EC_add_out_r_3_) );
  OAI22X1 U20116 ( .A0(n3583), .A1(n6301), .B0(top_core_EC_ss_n196), .B1(n3602), .Y(top_core_EC_add_in_r[3]) );
  XOR2X1 U20117 ( .A(top_core_Key[88]), .B(top_core_EC_add_in_r[32]), .Y(
        top_core_EC_add_out_r_32_) );
  OAI22X1 U20118 ( .A0(n3582), .A1(n6272), .B0(top_core_EC_ss_n204), .B1(n3610), .Y(top_core_EC_add_in_r[32]) );
  XOR2X1 U20119 ( .A(top_core_Key[72]), .B(top_core_EC_add_in_r[48]), .Y(
        top_core_EC_add_out_r_48_) );
  OAI22X1 U20120 ( .A0(n3583), .A1(n6256), .B0(top_core_EC_ss_n187), .B1(n3597), .Y(top_core_EC_add_in_r[48]) );
  XOR2X1 U20121 ( .A(top_core_Key[75]), .B(top_core_EC_add_in_r[51]), .Y(
        top_core_EC_add_out_r_51_) );
  OAI22X1 U20122 ( .A0(n3584), .A1(n6253), .B0(top_core_EC_ss_n183), .B1(n3595), .Y(top_core_EC_add_in_r[51]) );
  XOR2X1 U20123 ( .A(top_core_Key[91]), .B(top_core_EC_add_in_r[35]), .Y(
        top_core_EC_add_out_r_35_) );
  OAI22X1 U20124 ( .A0(n3582), .A1(n6269), .B0(top_core_EC_ss_n201), .B1(n3627), .Y(top_core_EC_add_in_r[35]) );
  XOR2X1 U20125 ( .A(top_core_Key[105]), .B(top_core_EC_add_in_r[17]), .Y(
        top_core_EC_add_out_r_17_) );
  OAI22X1 U20126 ( .A0(n3620), .A1(n6287), .B0(top_core_EC_ss_n221), .B1(n3607), .Y(top_core_EC_add_in_r[17]) );
  XOR2X1 U20127 ( .A(top_core_Key[114]), .B(top_core_EC_add_in_r[10]), .Y(
        top_core_EC_add_out_r_10_) );
  OAI22X1 U20128 ( .A0(n237), .A1(n6294), .B0(top_core_EC_ss_n246), .B1(n3611), 
        .Y(top_core_EC_add_in_r[10]) );
  XOR2X1 U20129 ( .A(top_core_Key[115]), .B(top_core_EC_add_in_r[11]), .Y(
        top_core_EC_add_out_r_11_) );
  OAI22X1 U20130 ( .A0(n237), .A1(n6293), .B0(top_core_EC_ss_n235), .B1(n3612), 
        .Y(top_core_EC_add_in_r[11]) );
  XOR2X1 U20131 ( .A(top_core_Key[108]), .B(top_core_EC_add_in_r[20]), .Y(
        top_core_EC_add_out_r_20_) );
  OAI22X1 U20132 ( .A0(n3621), .A1(n6284), .B0(top_core_EC_ss_n217), .B1(n3599), .Y(top_core_EC_add_in_r[20]) );
  XOR2X1 U20133 ( .A(top_core_Key[124]), .B(top_core_EC_add_in_r[4]), .Y(
        top_core_EC_add_out_r_4_) );
  OAI22X1 U20134 ( .A0(n3584), .A1(n6300), .B0(top_core_EC_ss_n185), .B1(n3596), .Y(top_core_EC_add_in_r[4]) );
  XOR2X1 U20135 ( .A(top_core_Key[109]), .B(top_core_EC_add_in_r[21]), .Y(
        top_core_EC_add_out_r_21_) );
  OAI22X1 U20136 ( .A0(n3622), .A1(n6283), .B0(top_core_EC_ss_n216), .B1(n3602), .Y(top_core_EC_add_in_r[21]) );
  XOR2X1 U20137 ( .A(top_core_Key[125]), .B(top_core_EC_add_in_r[5]), .Y(
        top_core_EC_add_out_r_5_) );
  OAI22X1 U20138 ( .A0(n3584), .A1(n6299), .B0(top_core_EC_ss_n174), .B1(n3591), .Y(top_core_EC_add_in_r[5]) );
  XOR2X1 U20139 ( .A(top_core_Key[110]), .B(top_core_EC_add_in_r[22]), .Y(
        top_core_EC_add_out_r_22_) );
  OAI22X1 U20140 ( .A0(n3622), .A1(n6282), .B0(top_core_EC_ss_n215), .B1(n3605), .Y(top_core_EC_add_in_r[22]) );
  XOR2X1 U20141 ( .A(top_core_Key[126]), .B(top_core_EC_add_in_r[6]), .Y(
        top_core_EC_add_out_r_6_) );
  OAI22X1 U20142 ( .A0(n3623), .A1(n6298), .B0(top_core_EC_ss_n163), .B1(n3592), .Y(top_core_EC_add_in_r[6]) );
  XOR2X1 U20143 ( .A(top_core_Key[111]), .B(top_core_EC_add_in_r[23]), .Y(
        top_core_EC_add_out_r_23_) );
  OAI22X1 U20144 ( .A0(n3585), .A1(n6281), .B0(top_core_EC_ss_n214), .B1(n3605), .Y(top_core_EC_add_in_r[23]) );
  XOR2X1 U20145 ( .A(top_core_Key[73]), .B(top_core_EC_add_in_r[49]), .Y(
        top_core_EC_add_out_r_49_) );
  OAI22X1 U20146 ( .A0(n3583), .A1(n6255), .B0(top_core_EC_ss_n186), .B1(n3597), .Y(top_core_EC_add_in_r[49]) );
  XOR2X1 U20147 ( .A(top_core_Key[89]), .B(top_core_EC_add_in_r[33]), .Y(
        top_core_EC_add_out_r_33_) );
  OAI22X1 U20148 ( .A0(n3582), .A1(n6271), .B0(top_core_EC_ss_n203), .B1(n3595), .Y(top_core_EC_add_in_r[33]) );
  XOR2X1 U20149 ( .A(top_core_Key[76]), .B(top_core_EC_add_in_r[52]), .Y(
        top_core_EC_add_out_r_52_) );
  OAI22X1 U20150 ( .A0(n3584), .A1(n6252), .B0(top_core_EC_ss_n182), .B1(n3595), .Y(top_core_EC_add_in_r[52]) );
  XOR2X1 U20151 ( .A(top_core_Key[77]), .B(top_core_EC_add_in_r[53]), .Y(
        top_core_EC_add_out_r_53_) );
  OAI22X1 U20152 ( .A0(n3584), .A1(n6251), .B0(top_core_EC_ss_n181), .B1(n3594), .Y(top_core_EC_add_in_r[53]) );
  XOR2X1 U20153 ( .A(top_core_Key[92]), .B(top_core_EC_add_in_r[36]), .Y(
        top_core_EC_add_out_r_36_) );
  OAI22X1 U20154 ( .A0(n3582), .A1(n6268), .B0(top_core_EC_ss_n200), .B1(n3593), .Y(top_core_EC_add_in_r[36]) );
  XOR2X1 U20155 ( .A(top_core_Key[78]), .B(top_core_EC_add_in_r[54]), .Y(
        top_core_EC_add_out_r_54_) );
  OAI22X1 U20156 ( .A0(n3584), .A1(n6250), .B0(top_core_EC_ss_n180), .B1(n3594), .Y(top_core_EC_add_in_r[54]) );
  XOR2X1 U20157 ( .A(top_core_Key[93]), .B(top_core_EC_add_in_r[37]), .Y(
        top_core_EC_add_out_r_37_) );
  OAI22X1 U20158 ( .A0(n3582), .A1(n6267), .B0(top_core_EC_ss_n199), .B1(n3608), .Y(top_core_EC_add_in_r[37]) );
  XOR2X1 U20159 ( .A(top_core_Key[79]), .B(top_core_EC_add_in_r[55]), .Y(
        top_core_EC_add_out_r_55_) );
  OAI22X1 U20160 ( .A0(n3584), .A1(n6249), .B0(top_core_EC_ss_n179), .B1(n3593), .Y(top_core_EC_add_in_r[55]) );
  XOR2X1 U20161 ( .A(top_core_Key[95]), .B(top_core_EC_add_in_r[39]), .Y(
        top_core_EC_add_out_r_39_) );
  OAI22X1 U20162 ( .A0(n3583), .A1(n6265), .B0(top_core_EC_ss_n197), .B1(n3602), .Y(top_core_EC_add_in_r[39]) );
  XOR2X1 U20163 ( .A(top_core_Key[94]), .B(top_core_EC_add_in_r[38]), .Y(
        top_core_EC_add_out_r_38_) );
  OAI22X1 U20164 ( .A0(n3582), .A1(n6266), .B0(top_core_EC_ss_n198), .B1(n3625), .Y(top_core_EC_add_in_r[38]) );
  XOR2X1 U20165 ( .A(top_core_Key[119]), .B(top_core_EC_add_in_r[15]), .Y(
        top_core_EC_add_out_r_15_) );
  OAI22X1 U20166 ( .A0(n3583), .A1(n6289), .B0(top_core_EC_ss_n223), .B1(n3592), .Y(top_core_EC_add_in_r[15]) );
  XOR2X1 U20167 ( .A(top_core_Key[112]), .B(top_core_EC_add_in_r[8]), .Y(
        top_core_EC_add_out_r_8_) );
  OAI22X1 U20168 ( .A0(n3586), .A1(n6296), .B0(top_core_EC_ss_n141), .B1(n3588), .Y(top_core_EC_add_in_r[8]) );
  XOR2X1 U20169 ( .A(top_core_Key[117]), .B(top_core_EC_add_in_r[13]), .Y(
        top_core_EC_add_out_r_13_) );
  OAI22X1 U20170 ( .A0(n3587), .A1(n6291), .B0(top_core_EC_ss_n225), .B1(n3588), .Y(top_core_EC_add_in_r[13]) );
  XOR2X1 U20171 ( .A(top_core_Key[118]), .B(top_core_EC_add_in_r[14]), .Y(
        top_core_EC_add_out_r_14_) );
  OAI22X1 U20172 ( .A0(n3584), .A1(n6290), .B0(top_core_EC_ss_n224), .B1(n3597), .Y(top_core_EC_add_in_r[14]) );
  XOR2X1 U20173 ( .A(top_core_Key[103]), .B(top_core_EC_add_in_r[31]), .Y(
        top_core_EC_add_out_r_31_) );
  OAI22X1 U20174 ( .A0(n3582), .A1(n6273), .B0(top_core_EC_ss_n205), .B1(n3609), .Y(top_core_EC_add_in_r[31]) );
  XOR2X1 U20175 ( .A(top_core_Key[101]), .B(top_core_EC_add_in_r[29]), .Y(
        top_core_EC_add_out_r_29_) );
  OAI22X1 U20176 ( .A0(n3582), .A1(n6275), .B0(top_core_EC_ss_n208), .B1(n3593), .Y(top_core_EC_add_in_r[29]) );
  XOR2X1 U20177 ( .A(top_core_Key[102]), .B(top_core_EC_add_in_r[30]), .Y(
        top_core_EC_add_out_r_30_) );
  OAI22X1 U20178 ( .A0(n3582), .A1(n6274), .B0(top_core_EC_ss_n206), .B1(n3599), .Y(top_core_EC_add_in_r[30]) );
  XOR2X1 U20179 ( .A(top_core_Key[87]), .B(top_core_EC_add_in_r[47]), .Y(
        top_core_EC_add_out_r_47_) );
  OAI22X1 U20180 ( .A0(n3583), .A1(n6257), .B0(top_core_EC_ss_n188), .B1(n3598), .Y(top_core_EC_add_in_r[47]) );
  XOR2X1 U20181 ( .A(top_core_Key[80]), .B(top_core_EC_add_in_r[40]), .Y(
        top_core_EC_add_out_r_40_) );
  OAI22X1 U20182 ( .A0(n3583), .A1(n6264), .B0(top_core_EC_ss_n195), .B1(n3601), .Y(top_core_EC_add_in_r[40]) );
  XOR2X1 U20183 ( .A(top_core_Key[82]), .B(top_core_EC_add_in_r[42]), .Y(
        top_core_EC_add_out_r_42_) );
  OAI22X1 U20184 ( .A0(n3583), .A1(n6262), .B0(top_core_EC_ss_n193), .B1(n3600), .Y(top_core_EC_add_in_r[42]) );
  XOR2X1 U20185 ( .A(top_core_Key[83]), .B(top_core_EC_add_in_r[43]), .Y(
        top_core_EC_add_out_r_43_) );
  OAI22X1 U20186 ( .A0(n3583), .A1(n6261), .B0(top_core_EC_ss_n192), .B1(n3600), .Y(top_core_EC_add_in_r[43]) );
  XOR2X1 U20187 ( .A(top_core_Key[85]), .B(top_core_EC_add_in_r[45]), .Y(
        top_core_EC_add_out_r_45_) );
  OAI22X1 U20188 ( .A0(n3583), .A1(n6259), .B0(top_core_EC_ss_n190), .B1(n3599), .Y(top_core_EC_add_in_r[45]) );
  XOR2X1 U20189 ( .A(top_core_Key[86]), .B(top_core_EC_add_in_r[46]), .Y(
        top_core_EC_add_out_r_46_) );
  OAI22X1 U20190 ( .A0(n3583), .A1(n6258), .B0(top_core_EC_ss_n189), .B1(n3598), .Y(top_core_EC_add_in_r[46]) );
  XOR2X1 U20191 ( .A(top_core_Key[96]), .B(top_core_EC_add_in_r[24]), .Y(
        top_core_EC_add_out_r_24_) );
  OAI22X1 U20192 ( .A0(n3587), .A1(n6280), .B0(top_core_EC_ss_n213), .B1(n3604), .Y(top_core_EC_add_in_r[24]) );
  XOR2X1 U20193 ( .A(top_core_Key[98]), .B(top_core_EC_add_in_r[26]), .Y(
        top_core_EC_add_out_r_26_) );
  OAI22X1 U20194 ( .A0(n3587), .A1(n6278), .B0(top_core_EC_ss_n211), .B1(n3603), .Y(top_core_EC_add_in_r[26]) );
  XOR2X1 U20195 ( .A(top_core_Key[99]), .B(top_core_EC_add_in_r[27]), .Y(
        top_core_EC_add_out_r_27_) );
  OAI22X1 U20196 ( .A0(n3587), .A1(n6277), .B0(top_core_EC_ss_n210), .B1(n3603), .Y(top_core_EC_add_in_r[27]) );
  XOR2X1 U20197 ( .A(top_core_Key[113]), .B(top_core_EC_add_in_r[9]), .Y(
        top_core_EC_add_out_r_9_) );
  OAI22X1 U20198 ( .A0(n3587), .A1(n6295), .B0(top_core_EC_ss_n130), .B1(n3599), .Y(top_core_EC_add_in_r[9]) );
  XOR2X1 U20199 ( .A(top_core_Key[116]), .B(top_core_EC_add_in_r[12]), .Y(
        top_core_EC_add_out_r_12_) );
  OAI22X1 U20200 ( .A0(n3622), .A1(n6292), .B0(top_core_EC_ss_n226), .B1(n3627), .Y(top_core_EC_add_in_r[12]) );
  XOR2X1 U20201 ( .A(top_core_Key[97]), .B(top_core_EC_add_in_r[25]), .Y(
        top_core_EC_add_out_r_25_) );
  OAI22X1 U20202 ( .A0(n3587), .A1(n6279), .B0(top_core_EC_ss_n212), .B1(n3604), .Y(top_core_EC_add_in_r[25]) );
  XOR2X1 U20203 ( .A(top_core_Key[100]), .B(top_core_EC_add_in_r[28]), .Y(
        top_core_EC_add_out_r_28_) );
  OAI22X1 U20204 ( .A0(n3582), .A1(n6276), .B0(top_core_EC_ss_n209), .B1(n3592), .Y(top_core_EC_add_in_r[28]) );
  XOR2X1 U20205 ( .A(top_core_Key[64]), .B(top_core_EC_add_in_r[56]), .Y(
        top_core_EC_add_out_r_56_) );
  OAI22X1 U20206 ( .A0(n3584), .A1(n6248), .B0(top_core_EC_ss_n178), .B1(n3593), .Y(top_core_EC_add_in_r[56]) );
  XOR2X1 U20207 ( .A(top_core_Key[81]), .B(top_core_EC_add_in_r[41]), .Y(
        top_core_EC_add_out_r_41_) );
  OAI22X1 U20208 ( .A0(n3583), .A1(n6263), .B0(top_core_EC_ss_n194), .B1(n3601), .Y(top_core_EC_add_in_r[41]) );
  XOR2X1 U20209 ( .A(top_core_Key[84]), .B(top_core_EC_add_in_r[44]), .Y(
        top_core_EC_add_out_r_44_) );
  OAI22X1 U20210 ( .A0(n3583), .A1(n6260), .B0(top_core_EC_ss_n191), .B1(n3599), .Y(top_core_EC_add_in_r[44]) );
  XOR2X1 U20211 ( .A(top_core_Key[65]), .B(top_core_EC_add_in_r[57]), .Y(
        top_core_EC_add_out_r_57_) );
  OAI22X1 U20212 ( .A0(n3584), .A1(n6247), .B0(top_core_EC_ss_n177), .B1(n3592), .Y(top_core_EC_add_in_r[57]) );
  XNOR2X1 U20213 ( .A(n6982), .B(top_core_KE_new_sboxw_0_), .Y(
        top_core_KE_n1072) );
  XNOR2X1 U20214 ( .A(n6717), .B(top_core_KE_new_sboxw_6_), .Y(
        top_core_KE_n1030) );
  XNOR2X1 U20215 ( .A(n6977), .B(top_core_KE_new_sboxw_24_), .Y(
        top_core_KE_n1128) );
  XNOR2X1 U20216 ( .A(n6384), .B(top_core_KE_new_sboxw_30_), .Y(
        top_core_KE_n1086) );
  XNOR2X1 U20217 ( .A(n6972), .B(top_core_KE_new_sboxw_1_), .Y(
        top_core_KE_n1065) );
  XNOR2X1 U20218 ( .A(n6967), .B(top_core_KE_new_sboxw_25_), .Y(
        top_core_KE_n1121) );
  XNOR2X1 U20219 ( .A(n6945), .B(top_core_KE_new_sboxw_3_), .Y(
        top_core_KE_n1051) );
  XNOR2X1 U20220 ( .A(n6900), .B(top_core_KE_new_sboxw_4_), .Y(
        top_core_KE_n1044) );
  XNOR2X1 U20221 ( .A(n6930), .B(top_core_KE_new_sboxw_27_), .Y(
        top_core_KE_n1107) );
  XNOR2X1 U20222 ( .A(n6854), .B(top_core_KE_new_sboxw_28_), .Y(
        top_core_KE_n1100) );
  OAI22X1 U20223 ( .A0(n1185), .A1(n13305), .B0(n13306), .B1(n13307), .Y(
        n13299) );
  AOI211X1 U20224 ( .A0(n6554), .A1(n1690), .B0(n13308), .C0(n13309), .Y(
        n13306) );
  OAI21XL U20225 ( .A0(n13238), .A1(n13310), .B0(n13311), .Y(n13309) );
  OAI22XL U20226 ( .A0(n7000), .A1(n151), .B0(n1500), .B1(n7001), .Y(
        top_core_KE_n4922) );
  OAI22XL U20227 ( .A0(n6999), .A1(n151), .B0(n1500), .B1(n7000), .Y(
        top_core_KE_n4921) );
  XNOR2X1 U20228 ( .A(n6695), .B(n6499), .Y(top_core_KE_n960) );
  XNOR2X1 U20229 ( .A(n6674), .B(n6492), .Y(top_core_KE_n946) );
  XNOR2X1 U20230 ( .A(n6655), .B(n6489), .Y(top_core_KE_n939) );
  XNOR2X1 U20231 ( .A(n6607), .B(n6486), .Y(top_core_KE_n932) );
  XNOR2X1 U20232 ( .A(n6524), .B(n6485), .Y(top_core_KE_n925) );
  XNOR2X1 U20233 ( .A(n6435), .B(n6484), .Y(top_core_KE_n917) );
  XNOR2X1 U20234 ( .A(n6314), .B(n6496), .Y(top_core_KE_n953) );
  XOR2X1 U20235 ( .A(top_core_KE_n1921), .B(n6496), .Y(top_core_KE_n1177) );
  XOR2X1 U20236 ( .A(top_core_KE_n1909), .B(n6483), .Y(top_core_KE_n1135) );
  XOR2X1 U20237 ( .A(top_core_KE_n1923), .B(n6499), .Y(top_core_KE_n1184) );
  XOR2X1 U20238 ( .A(top_core_KE_n1919), .B(n6492), .Y(top_core_KE_n1170) );
  XOR2X1 U20239 ( .A(top_core_KE_n1917), .B(n6489), .Y(top_core_KE_n1163) );
  XOR2X1 U20240 ( .A(top_core_KE_n1915), .B(n6486), .Y(top_core_KE_n1156) );
  XOR2X1 U20241 ( .A(top_core_KE_n1913), .B(n6485), .Y(top_core_KE_n1149) );
  XOR2X1 U20242 ( .A(top_core_KE_n1911), .B(n6484), .Y(top_core_KE_n1142) );
  XNOR2X1 U20243 ( .A(top_core_KE_new_sboxw_24_), .B(top_core_KE_n1923), .Y(
        top_core_KE_n1182) );
  XNOR2X1 U20244 ( .A(top_core_KE_new_sboxw_30_), .B(top_core_KE_n1911), .Y(
        top_core_KE_n1140) );
  BUFX4 U20245 ( .A(top_core_EC_ss_in[7]), .Y(n1506) );
  OAI22X1 U20246 ( .A0(n2385), .A1(n6297), .B0(n2421), .B1(n880), .Y(
        top_core_EC_ss_in[7]) );
  BUFX4 U20247 ( .A(top_core_EC_ss_in[87]), .Y(n1504) );
  OAI22X1 U20248 ( .A0(n2385), .A1(n6217), .B0(n2423), .B1(n881), .Y(
        top_core_EC_ss_in[87]) );
  BUFX4 U20249 ( .A(top_core_EC_ss_in[119]), .Y(n1528) );
  OAI22X1 U20250 ( .A0(n2391), .A1(n6185), .B0(n2455), .B1(n882), .Y(
        top_core_EC_ss_in[119]) );
  BUFX4 U20251 ( .A(top_core_EC_ss_in[39]), .Y(n1518) );
  OAI22X1 U20252 ( .A0(n2389), .A1(n6265), .B0(n2405), .B1(n883), .Y(
        top_core_EC_ss_in[39]) );
  BUFX4 U20253 ( .A(top_core_EC_ss_in[71]), .Y(n1509) );
  OAI22X1 U20254 ( .A0(n2386), .A1(n6233), .B0(n2418), .B1(n884), .Y(
        top_core_EC_ss_in[71]) );
  BUFX4 U20255 ( .A(top_core_EC_ss_in[111]), .Y(n1530) );
  OAI22X1 U20256 ( .A0(n2392), .A1(n6193), .B0(n2526), .B1(n885), .Y(
        top_core_EC_ss_in[111]) );
  BUFX4 U20257 ( .A(top_core_EC_ss_in[47]), .Y(n1515) );
  OAI22X1 U20258 ( .A0(n2388), .A1(n6257), .B0(n2409), .B1(n886), .Y(
        top_core_EC_ss_in[47]) );
  BUFX4 U20259 ( .A(top_core_EC_ss_in[23]), .Y(n1522) );
  OAI22X1 U20260 ( .A0(n2390), .A1(n6281), .B0(n2400), .B1(n887), .Y(
        top_core_EC_ss_in[23]) );
  BUFX4 U20261 ( .A(top_core_EC_ss_in[63]), .Y(n1511) );
  OAI22X1 U20262 ( .A0(n2387), .A1(n6241), .B0(n2415), .B1(n888), .Y(
        top_core_EC_ss_in[63]) );
  BUFX4 U20263 ( .A(top_core_EC_ss_in[127]), .Y(n1525) );
  OAI22X1 U20264 ( .A0(n2391), .A1(n6177), .B0(n2424), .B1(n889), .Y(
        top_core_EC_ss_in[127]) );
  BUFX4 U20265 ( .A(top_core_EC_ss_in[103]), .Y(n1532) );
  OAI22X1 U20266 ( .A0(n2393), .A1(n6201), .B0(n2397), .B1(n890), .Y(
        top_core_EC_ss_in[103]) );
  BUFX4 U20267 ( .A(top_core_EC_ss_in[15]), .Y(n1524) );
  OAI22X1 U20268 ( .A0(n2390), .A1(n6289), .B0(n2522), .B1(n891), .Y(
        top_core_EC_ss_in[15]) );
  BUFX4 U20269 ( .A(top_core_EC_ss_in[79]), .Y(n1507) );
  OAI22X1 U20270 ( .A0(n2385), .A1(n6225), .B0(n2420), .B1(n892), .Y(
        top_core_EC_ss_in[79]) );
  BUFX4 U20271 ( .A(top_core_EC_ss_in[55]), .Y(n1513) );
  OAI22X1 U20272 ( .A0(n2387), .A1(n6249), .B0(n2412), .B1(n893), .Y(
        top_core_EC_ss_in[55]) );
  BUFX4 U20273 ( .A(top_core_EC_ss_in[95]), .Y(n1502) );
  OAI22X1 U20274 ( .A0(n2384), .A1(n6209), .B0(n2411), .B1(n894), .Y(
        top_core_EC_ss_in[95]) );
  BUFX4 U20275 ( .A(top_core_EC_ss_in[31]), .Y(n1520) );
  OAI22X1 U20276 ( .A0(n2389), .A1(n6273), .B0(n2403), .B1(n895), .Y(
        top_core_EC_ss_in[31]) );
  OAI22X1 U20277 ( .A0(n824), .A1(n3631), .B0(n192), .B1(n3639), .Y(
        top_core_EC_N207) );
  OAI22X1 U20278 ( .A0(n875), .A1(n3628), .B0(n193), .B1(n3636), .Y(
        top_core_EC_N208) );
  OAI22X1 U20279 ( .A0(n848), .A1(n3632), .B0(n128), .B1(n3640), .Y(
        top_core_EC_N209) );
  OAI22X1 U20280 ( .A0(n834), .A1(n3632), .B0(n194), .B1(n3640), .Y(
        top_core_EC_N210) );
  OAI22X1 U20281 ( .A0(n857), .A1(n3632), .B0(n195), .B1(n3640), .Y(
        top_core_EC_N211) );
  OAI22X1 U20282 ( .A0(n888), .A1(n3632), .B0(n196), .B1(n3640), .Y(
        top_core_EC_N212) );
  OAI22X1 U20283 ( .A0(n816), .A1(n3632), .B0(n197), .B1(n3640), .Y(
        top_core_EC_N213) );
  OAI22X1 U20284 ( .A0(n788), .A1(n3632), .B0(n198), .B1(n3640), .Y(
        top_core_EC_N214) );
  OAI22X1 U20285 ( .A0(n787), .A1(n3632), .B0(n199), .B1(n3640), .Y(
        top_core_EC_N215) );
  OAI22X1 U20286 ( .A0(n872), .A1(n3632), .B0(n200), .B1(n3640), .Y(
        top_core_EC_N216) );
  OAI22X1 U20287 ( .A0(n838), .A1(n3632), .B0(n152), .B1(n3640), .Y(
        top_core_EC_N217) );
  OAI22X1 U20288 ( .A0(n839), .A1(n3632), .B0(n127), .B1(n3640), .Y(
        top_core_EC_N218) );
  OAI22X1 U20289 ( .A0(n862), .A1(n3632), .B0(n126), .B1(n3640), .Y(
        top_core_EC_N219) );
  OAI22X1 U20290 ( .A0(n884), .A1(n3632), .B0(n153), .B1(n3640), .Y(
        top_core_EC_N220) );
  OAI22X1 U20291 ( .A0(n809), .A1(n3633), .B0(n201), .B1(n3641), .Y(
        top_core_EC_N221) );
  OAI22X1 U20292 ( .A0(n810), .A1(n3633), .B0(n154), .B1(n3641), .Y(
        top_core_EC_N222) );
  OAI22X1 U20293 ( .A0(n776), .A1(n3633), .B0(n202), .B1(n3641), .Y(
        top_core_EC_N223) );
  OAI22X1 U20294 ( .A0(n869), .A1(n3633), .B0(n203), .B1(n3641), .Y(
        top_core_EC_N224) );
  OAI22X1 U20295 ( .A0(n829), .A1(n3633), .B0(n155), .B1(n3641), .Y(
        top_core_EC_N225) );
  OAI22X1 U20296 ( .A0(n828), .A1(n3633), .B0(n204), .B1(n3641), .Y(
        top_core_EC_N226) );
  OAI22X1 U20297 ( .A0(n853), .A1(n3633), .B0(n205), .B1(n3641), .Y(
        top_core_EC_N227) );
  OAI22X1 U20298 ( .A0(n892), .A1(n3633), .B0(n206), .B1(n3641), .Y(
        top_core_EC_N228) );
  OAI22X1 U20299 ( .A0(n775), .A1(n3633), .B0(n207), .B1(n3641), .Y(
        top_core_EC_N229) );
  OAI22X1 U20300 ( .A0(n772), .A1(n3633), .B0(n208), .B1(n3641), .Y(
        top_core_EC_N230) );
  OAI22X1 U20301 ( .A0(n782), .A1(n3633), .B0(n209), .B1(n3641), .Y(
        top_core_EC_N231) );
  OAI22X1 U20302 ( .A0(n855), .A1(n3633), .B0(n210), .B1(n3641), .Y(
        top_core_EC_N232) );
  OAI22X1 U20303 ( .A0(n802), .A1(n3634), .B0(n156), .B1(n3642), .Y(
        top_core_EC_N233) );
  OAI22X1 U20304 ( .A0(n801), .A1(n3634), .B0(n125), .B1(n3642), .Y(
        top_core_EC_N234) );
  OAI22X1 U20305 ( .A0(n833), .A1(n3634), .B0(n124), .B1(n3642), .Y(
        top_core_EC_N235) );
  OAI22X1 U20306 ( .A0(n881), .A1(n3634), .B0(n123), .B1(n3642), .Y(
        top_core_EC_N236) );
  OAI22X1 U20307 ( .A0(n820), .A1(n3634), .B0(n211), .B1(n3642), .Y(
        top_core_EC_N237) );
  OAI22X1 U20308 ( .A0(n786), .A1(n3634), .B0(n157), .B1(n3642), .Y(
        top_core_EC_N238) );
  OAI22X1 U20309 ( .A0(n796), .A1(n3634), .B0(n212), .B1(n3642), .Y(
        top_core_EC_N239) );
  OAI22X1 U20310 ( .A0(n879), .A1(n3634), .B0(n213), .B1(n3642), .Y(
        top_core_EC_N240) );
  OAI22X1 U20311 ( .A0(n846), .A1(n3634), .B0(n122), .B1(n3642), .Y(
        top_core_EC_N241) );
  OAI22X1 U20312 ( .A0(n851), .A1(n3634), .B0(n214), .B1(n3642), .Y(
        top_core_EC_N242) );
  OAI22X1 U20313 ( .A0(n866), .A1(n3634), .B0(n215), .B1(n3642), .Y(
        top_core_EC_N243) );
  OAI22X1 U20314 ( .A0(n894), .A1(n3634), .B0(n216), .B1(n3642), .Y(
        top_core_EC_N244) );
  OAI22X1 U20315 ( .A0(n818), .A1(n3632), .B0(n217), .B1(n3640), .Y(
        top_core_EC_N245) );
  OAI22X1 U20316 ( .A0(n793), .A1(n3633), .B0(n218), .B1(n3641), .Y(
        top_core_EC_N246) );
  OAI22X1 U20317 ( .A0(n792), .A1(n3634), .B0(n219), .B1(n3642), .Y(
        top_core_EC_N247) );
  OAI22X1 U20318 ( .A0(n876), .A1(n3629), .B0(n220), .B1(n3637), .Y(
        top_core_EC_N248) );
  OAI22X1 U20319 ( .A0(n842), .A1(n3632), .B0(n158), .B1(n3640), .Y(
        top_core_EC_N249) );
  OAI22X1 U20320 ( .A0(n843), .A1(n3632), .B0(n134), .B1(n3640), .Y(
        top_core_EC_N250) );
  OAI22X1 U20321 ( .A0(n864), .A1(n3630), .B0(n133), .B1(n3638), .Y(
        top_core_EC_N251) );
  OAI22X1 U20322 ( .A0(n890), .A1(n3631), .B0(n159), .B1(n3639), .Y(
        top_core_EC_N252) );
  OAI22X1 U20323 ( .A0(n798), .A1(n3628), .B0(n221), .B1(n3636), .Y(
        top_core_EC_N253) );
  OAI22X1 U20324 ( .A0(n800), .A1(n3635), .B0(n160), .B1(n3643), .Y(
        top_core_EC_N254) );
  OAI22X1 U20325 ( .A0(n821), .A1(n3633), .B0(n222), .B1(n3641), .Y(
        top_core_EC_N255) );
  OAI22X1 U20326 ( .A0(n873), .A1(n3634), .B0(n223), .B1(n3642), .Y(
        top_core_EC_N256) );
  OAI22X1 U20327 ( .A0(n832), .A1(n3635), .B0(n161), .B1(n3643), .Y(
        top_core_EC_N257) );
  OAI22X1 U20328 ( .A0(n831), .A1(n3635), .B0(n224), .B1(n3643), .Y(
        top_core_EC_N258) );
  OAI22X1 U20329 ( .A0(n854), .A1(n3635), .B0(n225), .B1(n3643), .Y(
        top_core_EC_N259) );
  OAI22X1 U20330 ( .A0(n885), .A1(n3635), .B0(n226), .B1(n3643), .Y(
        top_core_EC_N260) );
  OAI22X1 U20331 ( .A0(n777), .A1(n3635), .B0(n227), .B1(n3643), .Y(
        top_core_EC_N261) );
  OAI22X1 U20332 ( .A0(n773), .A1(n3635), .B0(n228), .B1(n3643), .Y(
        top_core_EC_N262) );
  OAI22X1 U20333 ( .A0(n783), .A1(n3635), .B0(n229), .B1(n3643), .Y(
        top_core_EC_N263) );
  OAI22X1 U20334 ( .A0(n860), .A1(n3635), .B0(n230), .B1(n3643), .Y(
        top_core_EC_N264) );
  OAI22X1 U20335 ( .A0(n812), .A1(n3635), .B0(n162), .B1(n3643), .Y(
        top_core_EC_N265) );
  OAI22X1 U20336 ( .A0(n811), .A1(n3635), .B0(n132), .B1(n3643), .Y(
        top_core_EC_N266) );
  OAI22X1 U20337 ( .A0(n836), .A1(n3635), .B0(n131), .B1(n3643), .Y(
        top_core_EC_N267) );
  OAI22X1 U20338 ( .A0(n882), .A1(n3635), .B0(n130), .B1(n3643), .Y(
        top_core_EC_N268) );
  OAI22X1 U20339 ( .A0(n807), .A1(n3633), .B0(n231), .B1(n3641), .Y(
        top_core_EC_N269) );
  OAI22X1 U20340 ( .A0(n791), .A1(n3634), .B0(n163), .B1(n3642), .Y(
        top_core_EC_N270) );
  OAI22X1 U20341 ( .A0(n779), .A1(n3629), .B0(n232), .B1(n3637), .Y(
        top_core_EC_N271) );
  OAI22X1 U20342 ( .A0(n870), .A1(n3630), .B0(n233), .B1(n3638), .Y(
        top_core_EC_N272) );
  OAI22X1 U20343 ( .A0(n827), .A1(n3630), .B0(n129), .B1(n3638), .Y(
        top_core_EC_N273) );
  OAI22X1 U20344 ( .A0(n830), .A1(n3631), .B0(n234), .B1(n3639), .Y(
        top_core_EC_N274) );
  OAI22X1 U20345 ( .A0(n858), .A1(n3628), .B0(n235), .B1(n3636), .Y(
        top_core_EC_N275) );
  OAI22X1 U20346 ( .A0(n889), .A1(n3635), .B0(n236), .B1(n3643), .Y(
        top_core_EC_N276) );
  XNOR2X1 U20347 ( .A(top_core_KE_new_sboxw_25_), .B(top_core_KE_n1921), .Y(
        top_core_KE_n1175) );
  XNOR2X1 U20348 ( .A(top_core_KE_new_sboxw_27_), .B(top_core_KE_n1917), .Y(
        top_core_KE_n1161) );
  XNOR2X1 U20349 ( .A(top_core_KE_new_sboxw_28_), .B(top_core_KE_n1915), .Y(
        top_core_KE_n1154) );
  XOR2X1 U20350 ( .A(top_core_KE_new_sboxw_192_15_), .B(top_core_KE_n1925), 
        .Y(top_core_KE_n1682) );
  XOR2X1 U20351 ( .A(top_core_KE_new_sboxw_192_13_), .B(top_core_KE_n1929), 
        .Y(top_core_KE_n1698) );
  XOR2X1 U20352 ( .A(top_core_KE_new_sboxw_192_10_), .B(top_core_KE_n1935), 
        .Y(top_core_KE_n1722) );
  XOR2X1 U20353 ( .A(top_core_KE_new_sboxw_192_7_), .B(top_core_KE_n1941), .Y(
        top_core_KE_n1746) );
  XOR2X1 U20354 ( .A(top_core_KE_new_sboxw_192_5_), .B(top_core_KE_n1945), .Y(
        top_core_KE_n1762) );
  XOR2X1 U20355 ( .A(top_core_KE_new_sboxw_192_2_), .B(top_core_KE_n1951), .Y(
        top_core_KE_n1786) );
  XOR2X1 U20356 ( .A(top_core_KE_new_sboxw_192_31_), .B(top_core_KE_n1957), 
        .Y(top_core_KE_n1810) );
  XOR2X1 U20357 ( .A(top_core_KE_new_sboxw_192_29_), .B(top_core_KE_n1961), 
        .Y(top_core_KE_n1826) );
  XOR2X1 U20358 ( .A(top_core_KE_new_sboxw_192_26_), .B(top_core_KE_n1967), 
        .Y(top_core_KE_n1850) );
  OAI22X1 U20359 ( .A0(n769), .A1(n3628), .B0(n6095), .B1(n3636), .Y(
        top_core_EC_N149) );
  OAI22X1 U20360 ( .A0(n771), .A1(n3628), .B0(n6102), .B1(n3636), .Y(
        top_core_EC_N150) );
  OAI22X1 U20361 ( .A0(n780), .A1(n3628), .B0(n6100), .B1(n3636), .Y(
        top_core_EC_N151) );
  OAI22X1 U20362 ( .A0(n856), .A1(n3628), .B0(n6098), .B1(n3636), .Y(
        top_core_EC_N152) );
  OAI22X1 U20363 ( .A0(n806), .A1(n3628), .B0(n6094), .B1(n3636), .Y(
        top_core_EC_N153) );
  OAI22X1 U20364 ( .A0(n805), .A1(n3628), .B0(n6097), .B1(n3636), .Y(
        top_core_EC_N154) );
  OAI22X1 U20365 ( .A0(n826), .A1(n3628), .B0(n6093), .B1(n3636), .Y(
        top_core_EC_N155) );
  OAI22X1 U20366 ( .A0(n880), .A1(n3628), .B0(n6096), .B1(n3636), .Y(
        top_core_EC_N156) );
  OAI22X1 U20367 ( .A0(n808), .A1(n3628), .B0(n5047), .B1(n3636), .Y(
        top_core_EC_N157) );
  OAI22X1 U20368 ( .A0(n768), .A1(n3628), .B0(n5046), .B1(n3636), .Y(
        top_core_EC_N158) );
  OAI22X1 U20369 ( .A0(n825), .A1(n3628), .B0(n5045), .B1(n3636), .Y(
        top_core_EC_N159) );
  OAI22X1 U20370 ( .A0(n877), .A1(n3628), .B0(n5043), .B1(n3636), .Y(
        top_core_EC_N160) );
  OAI22X1 U20371 ( .A0(n852), .A1(n3629), .B0(n5042), .B1(n3637), .Y(
        top_core_EC_N161) );
  OAI22X1 U20372 ( .A0(n835), .A1(n3629), .B0(n5041), .B1(n3637), .Y(
        top_core_EC_N162) );
  OAI22X1 U20373 ( .A0(n859), .A1(n3629), .B0(n5040), .B1(n3637), .Y(
        top_core_EC_N163) );
  OAI22X1 U20374 ( .A0(n891), .A1(n3629), .B0(n5039), .B1(n3637), .Y(
        top_core_EC_N164) );
  OAI22X1 U20375 ( .A0(n817), .A1(n3629), .B0(n5314), .B1(n3637), .Y(
        top_core_EC_N165) );
  OAI22X1 U20376 ( .A0(n790), .A1(n3629), .B0(n5317), .B1(n3637), .Y(
        top_core_EC_N166) );
  OAI22X1 U20377 ( .A0(n789), .A1(n3629), .B0(n5316), .B1(n3637), .Y(
        top_core_EC_N167) );
  OAI22X1 U20378 ( .A0(n874), .A1(n3629), .B0(n5313), .B1(n3637), .Y(
        top_core_EC_N168) );
  OAI22X1 U20379 ( .A0(n840), .A1(n3629), .B0(n5312), .B1(n3637), .Y(
        top_core_EC_N169) );
  OAI22X1 U20380 ( .A0(n841), .A1(n3629), .B0(n5311), .B1(n3637), .Y(
        top_core_EC_N170) );
  OAI22X1 U20381 ( .A0(n863), .A1(n3629), .B0(n5310), .B1(n3637), .Y(
        top_core_EC_N171) );
  OAI22X1 U20382 ( .A0(n887), .A1(n3629), .B0(n5309), .B1(n3637), .Y(
        top_core_EC_N172) );
  OAI22X1 U20383 ( .A0(n815), .A1(n3630), .B0(n4841), .B1(n3638), .Y(
        top_core_EC_N173) );
  OAI22X1 U20384 ( .A0(n797), .A1(n3630), .B0(n4850), .B1(n3638), .Y(
        top_core_EC_N174) );
  OAI22X1 U20385 ( .A0(n785), .A1(n3630), .B0(n4848), .B1(n3638), .Y(
        top_core_EC_N175) );
  OAI22X1 U20386 ( .A0(n871), .A1(n3630), .B0(n4847), .B1(n3638), .Y(
        top_core_EC_N176) );
  OAI22X1 U20387 ( .A0(n850), .A1(n3630), .B0(n4836), .B1(n3638), .Y(
        top_core_EC_N177) );
  OAI22X1 U20388 ( .A0(n849), .A1(n3630), .B0(n4846), .B1(n3638), .Y(
        top_core_EC_N178) );
  OAI22X1 U20389 ( .A0(n867), .A1(n3630), .B0(n4832), .B1(n3638), .Y(
        top_core_EC_N179) );
  OAI22X1 U20390 ( .A0(n895), .A1(n3630), .B0(n4845), .B1(n3638), .Y(
        top_core_EC_N180) );
  OAI22X1 U20391 ( .A0(n778), .A1(n3630), .B0(n5786), .B1(n3638), .Y(
        top_core_EC_N181) );
  OAI22X1 U20392 ( .A0(n774), .A1(n3630), .B0(n5789), .B1(n3638), .Y(
        top_core_EC_N182) );
  OAI22X1 U20393 ( .A0(n784), .A1(n3630), .B0(n5788), .B1(n3638), .Y(
        top_core_EC_N183) );
  OAI22X1 U20394 ( .A0(n861), .A1(n3630), .B0(n5785), .B1(n3638), .Y(
        top_core_EC_N184) );
  OAI22X1 U20395 ( .A0(n814), .A1(n3631), .B0(n5784), .B1(n3639), .Y(
        top_core_EC_N185) );
  OAI22X1 U20396 ( .A0(n813), .A1(n3631), .B0(n5783), .B1(n3639), .Y(
        top_core_EC_N186) );
  OAI22X1 U20397 ( .A0(n837), .A1(n3631), .B0(n5782), .B1(n3639), .Y(
        top_core_EC_N187) );
  OAI22X1 U20398 ( .A0(n883), .A1(n3631), .B0(n5781), .B1(n3639), .Y(
        top_core_EC_N188) );
  OAI22X1 U20399 ( .A0(n799), .A1(n3631), .B0(n5395), .B1(n3639), .Y(
        top_core_EC_N189) );
  OAI22X1 U20400 ( .A0(n804), .A1(n3631), .B0(n5404), .B1(n3639), .Y(
        top_core_EC_N190) );
  OAI22X1 U20401 ( .A0(n770), .A1(n3631), .B0(n5402), .B1(n3639), .Y(
        top_core_EC_N191) );
  OAI22X1 U20402 ( .A0(n868), .A1(n3631), .B0(n5401), .B1(n3639), .Y(
        top_core_EC_N192) );
  OAI22X1 U20403 ( .A0(n823), .A1(n3631), .B0(n5394), .B1(n3639), .Y(
        top_core_EC_N193) );
  OAI22X1 U20404 ( .A0(n822), .A1(n3631), .B0(n5400), .B1(n3639), .Y(
        top_core_EC_N194) );
  OAI22X1 U20405 ( .A0(n847), .A1(n3631), .B0(n5393), .B1(n3639), .Y(
        top_core_EC_N195) );
  OAI22X1 U20406 ( .A0(n886), .A1(n3631), .B0(n5399), .B1(n3639), .Y(
        top_core_EC_N196) );
  OAI22X1 U20407 ( .A0(n819), .A1(n3635), .B0(n4960), .B1(n3643), .Y(
        top_core_EC_N197) );
  OAI22X1 U20408 ( .A0(n795), .A1(n3629), .B0(n4963), .B1(n3637), .Y(
        top_core_EC_N198) );
  OAI22X1 U20409 ( .A0(n794), .A1(n3632), .B0(n4962), .B1(n3640), .Y(
        top_core_EC_N199) );
  OAI22X1 U20410 ( .A0(n878), .A1(n3630), .B0(n4959), .B1(n3638), .Y(
        top_core_EC_N200) );
  OAI22X1 U20411 ( .A0(n844), .A1(n3631), .B0(n4958), .B1(n3639), .Y(
        top_core_EC_N201) );
  OAI22X1 U20412 ( .A0(n845), .A1(n3628), .B0(n4957), .B1(n3636), .Y(
        top_core_EC_N202) );
  OAI22X1 U20413 ( .A0(n865), .A1(n3635), .B0(n4955), .B1(n3643), .Y(
        top_core_EC_N203) );
  OAI22X1 U20414 ( .A0(n893), .A1(n3633), .B0(n4950), .B1(n3641), .Y(
        top_core_EC_N204) );
  OAI22X1 U20415 ( .A0(n803), .A1(n3634), .B0(n5233), .B1(n3642), .Y(
        top_core_EC_N205) );
  OAI22X1 U20416 ( .A0(n781), .A1(n3629), .B0(n5232), .B1(n3637), .Y(
        top_core_EC_N206) );
  XNOR2X1 U20417 ( .A(n6667), .B(top_core_KE_new_sboxw_10_), .Y(
        top_core_KE_n1002) );
  XNOR2X1 U20418 ( .A(n6480), .B(top_core_KE_new_sboxw_13_), .Y(
        top_core_KE_n981) );
  XNOR2X1 U20419 ( .A(n6394), .B(top_core_KE_new_sboxw_15_), .Y(
        top_core_KE_n967) );
  INVX1 U20420 ( .A(top_core_EC_n944), .Y(n6306) );
  OAI22XL U20421 ( .A0(n2), .A1(n4256), .B0(n4259), .B1(n2451), .Y(
        top_core_EC_n1295) );
  XNOR2X1 U20422 ( .A(top_core_KE_new_sboxw_192_15_), .B(n6394), .Y(
        top_core_KE_n1426) );
  XNOR2X1 U20423 ( .A(top_core_KE_new_sboxw_192_13_), .B(n6480), .Y(
        top_core_KE_n1442) );
  XNOR2X1 U20424 ( .A(top_core_KE_new_sboxw_192_10_), .B(n6667), .Y(
        top_core_KE_n1466) );
  XNOR2X1 U20425 ( .A(top_core_KE_new_sboxw_192_7_), .B(n6328), .Y(
        top_core_KE_n1490) );
  XNOR2X1 U20426 ( .A(top_core_KE_new_sboxw_192_5_), .B(n6820), .Y(
        top_core_KE_n1506) );
  XNOR2X1 U20427 ( .A(top_core_KE_new_sboxw_192_2_), .B(n6961), .Y(
        top_core_KE_n1530) );
  XNOR2X1 U20428 ( .A(top_core_KE_new_sboxw_192_31_), .B(n6377), .Y(
        top_core_KE_n1554) );
  XNOR2X1 U20429 ( .A(top_core_KE_new_sboxw_192_29_), .B(n6781), .Y(
        top_core_KE_n1570) );
  XNOR2X1 U20430 ( .A(top_core_KE_new_sboxw_192_26_), .B(n6955), .Y(
        top_core_KE_n1594) );
  XNOR2X1 U20431 ( .A(n6341), .B(top_core_KE_new_sboxw_31_), .Y(
        top_core_KE_n902) );
  NAND2BX1 U20432 ( .AN(top_core_EC_n946), .B(n2391), .Y(top_core_EC_n868) );
  XNOR2X1 U20433 ( .A(top_core_KE_new_sboxw_15_), .B(top_core_KE_n2631), .Y(
        top_core_KE_n1741) );
  XNOR2X1 U20434 ( .A(top_core_KE_new_sboxw_13_), .B(top_core_KE_n2639), .Y(
        top_core_KE_n1757) );
  XNOR2X1 U20435 ( .A(top_core_KE_new_sboxw_10_), .B(top_core_KE_n2651), .Y(
        top_core_KE_n1781) );
  XNOR2X1 U20436 ( .A(top_core_KE_new_sboxw_7_), .B(top_core_KE_n2663), .Y(
        top_core_KE_n1805) );
  XNOR2X1 U20437 ( .A(top_core_KE_new_sboxw_5_), .B(top_core_KE_n2671), .Y(
        top_core_KE_n1821) );
  XNOR2X1 U20438 ( .A(top_core_KE_new_sboxw_2_), .B(top_core_KE_n2683), .Y(
        top_core_KE_n1845) );
  OAI21XL U20439 ( .A0(n6308), .A1(n1), .B0(top_core_EC_n1027), .Y(
        top_core_EC_n1299) );
  OAI21XL U20440 ( .A0(top_core_EC_n1024), .A1(n6308), .B0(n1), .Y(
        top_core_EC_n1027) );
  XNOR2X1 U20441 ( .A(top_core_KE_new_sboxw_31_), .B(top_core_KE_n2559), .Y(
        top_core_KE_n1613) );
  XNOR2X1 U20442 ( .A(top_core_KE_new_sboxw_29_), .B(top_core_KE_n2569), .Y(
        top_core_KE_n1629) );
  XNOR2X1 U20443 ( .A(top_core_KE_new_sboxw_26_), .B(top_core_KE_n2584), .Y(
        top_core_KE_n1653) );
  XOR2X1 U20444 ( .A(top_core_KE_new_sboxw_192_14_), .B(top_core_KE_n1927), 
        .Y(top_core_KE_n1690) );
  XOR2X1 U20445 ( .A(top_core_KE_new_sboxw_192_8_), .B(top_core_KE_n1939), .Y(
        top_core_KE_n1738) );
  XOR2X1 U20446 ( .A(top_core_KE_new_sboxw_192_6_), .B(top_core_KE_n1943), .Y(
        top_core_KE_n1754) );
  XOR2X1 U20447 ( .A(top_core_KE_new_sboxw_192_0_), .B(top_core_KE_n1955), .Y(
        top_core_KE_n1802) );
  XOR2X1 U20448 ( .A(top_core_KE_new_sboxw_192_30_), .B(top_core_KE_n1959), 
        .Y(top_core_KE_n1818) );
  XOR2X1 U20449 ( .A(top_core_KE_new_sboxw_192_24_), .B(top_core_KE_n1971), 
        .Y(top_core_KE_n1869) );
  XOR2X1 U20450 ( .A(top_core_KE_new_sboxw_192_9_), .B(top_core_KE_n1937), .Y(
        top_core_KE_n1730) );
  XOR2X1 U20451 ( .A(top_core_KE_new_sboxw_192_1_), .B(top_core_KE_n1953), .Y(
        top_core_KE_n1794) );
  XOR2X1 U20452 ( .A(top_core_KE_new_sboxw_192_25_), .B(top_core_KE_n1969), 
        .Y(top_core_KE_n1858) );
  XOR2X1 U20453 ( .A(top_core_KE_new_sboxw_192_12_), .B(top_core_KE_n1931), 
        .Y(top_core_KE_n1706) );
  XOR2X1 U20454 ( .A(top_core_KE_new_sboxw_192_11_), .B(top_core_KE_n1933), 
        .Y(top_core_KE_n1714) );
  XOR2X1 U20455 ( .A(top_core_KE_new_sboxw_192_4_), .B(top_core_KE_n1947), .Y(
        top_core_KE_n1770) );
  XOR2X1 U20456 ( .A(top_core_KE_new_sboxw_192_3_), .B(top_core_KE_n1949), .Y(
        top_core_KE_n1778) );
  XOR2X1 U20457 ( .A(top_core_KE_new_sboxw_192_28_), .B(top_core_KE_n1963), 
        .Y(top_core_KE_n1834) );
  XOR2X1 U20458 ( .A(top_core_KE_new_sboxw_192_27_), .B(top_core_KE_n1965), 
        .Y(top_core_KE_n1842) );
  XNOR2X1 U20459 ( .A(top_core_KE_new_sboxw_192_14_), .B(n6402), .Y(
        top_core_KE_n1434) );
  XNOR2X1 U20460 ( .A(top_core_KE_new_sboxw_192_8_), .B(n6689), .Y(
        top_core_KE_n1482) );
  XNOR2X1 U20461 ( .A(top_core_KE_new_sboxw_192_6_), .B(n6717), .Y(
        top_core_KE_n1498) );
  XNOR2X1 U20462 ( .A(top_core_KE_new_sboxw_192_0_), .B(n6982), .Y(
        top_core_KE_n1546) );
  XNOR2X1 U20463 ( .A(top_core_KE_new_sboxw_192_30_), .B(n6384), .Y(
        top_core_KE_n1562) );
  XNOR2X1 U20464 ( .A(top_core_KE_new_sboxw_192_24_), .B(n6977), .Y(
        top_core_KE_n1610) );
  XNOR2X1 U20465 ( .A(n6689), .B(top_core_KE_new_sboxw_8_), .Y(
        top_core_KE_n1016) );
  XNOR2X1 U20466 ( .A(n6402), .B(top_core_KE_new_sboxw_14_), .Y(
        top_core_KE_n974) );
  XNOR2X1 U20467 ( .A(top_core_KE_new_sboxw_192_9_), .B(n6682), .Y(
        top_core_KE_n1474) );
  XNOR2X1 U20468 ( .A(top_core_KE_new_sboxw_192_1_), .B(n6972), .Y(
        top_core_KE_n1538) );
  XNOR2X1 U20469 ( .A(top_core_KE_new_sboxw_192_25_), .B(n6967), .Y(
        top_core_KE_n1602) );
  XNOR2X1 U20470 ( .A(top_core_KE_new_sboxw_192_12_), .B(n6560), .Y(
        top_core_KE_n1450) );
  XNOR2X1 U20471 ( .A(top_core_KE_new_sboxw_192_11_), .B(n6639), .Y(
        top_core_KE_n1458) );
  XNOR2X1 U20472 ( .A(top_core_KE_new_sboxw_192_4_), .B(n6900), .Y(
        top_core_KE_n1514) );
  XNOR2X1 U20473 ( .A(top_core_KE_new_sboxw_192_3_), .B(n6945), .Y(
        top_core_KE_n1522) );
  XNOR2X1 U20474 ( .A(top_core_KE_new_sboxw_192_28_), .B(n6854), .Y(
        top_core_KE_n1578) );
  XNOR2X1 U20475 ( .A(top_core_KE_new_sboxw_192_27_), .B(n6930), .Y(
        top_core_KE_n1586) );
  XNOR2X1 U20476 ( .A(n6682), .B(top_core_KE_new_sboxw_9_), .Y(
        top_core_KE_n1009) );
  XNOR2X1 U20477 ( .A(n6639), .B(top_core_KE_new_sboxw_11_), .Y(
        top_core_KE_n995) );
  XNOR2X1 U20478 ( .A(n6560), .B(top_core_KE_new_sboxw_12_), .Y(
        top_core_KE_n988) );
  INVX1 U20479 ( .A(top_core_KE_n897), .Y(n7020) );
  XNOR2X1 U20480 ( .A(top_core_KE_n1921), .B(n6463), .Y(top_core_KE_n1666) );
  XNOR2X1 U20481 ( .A(top_core_KE_n1923), .B(n6466), .Y(top_core_KE_n1674) );
  XNOR2X1 U20482 ( .A(top_core_KE_n1919), .B(n6461), .Y(top_core_KE_n1658) );
  XNOR2X1 U20483 ( .A(top_core_KE_n1917), .B(n6458), .Y(top_core_KE_n1650) );
  XNOR2X1 U20484 ( .A(top_core_KE_n1915), .B(n6455), .Y(top_core_KE_n1642) );
  XNOR2X1 U20485 ( .A(top_core_KE_n1913), .B(n6452), .Y(top_core_KE_n1634) );
  XNOR2X1 U20486 ( .A(top_core_KE_n1911), .B(n6449), .Y(top_core_KE_n1626) );
  XNOR2X1 U20487 ( .A(top_core_KE_n1909), .B(n6448), .Y(top_core_KE_n1618) );
  XNOR2X1 U20488 ( .A(n6359), .B(top_core_KE_n1957), .Y(top_core_KE_n1303) );
  XNOR2X1 U20489 ( .A(n6785), .B(top_core_KE_n1941), .Y(top_core_KE_n1247) );
  XNOR2X1 U20490 ( .A(n6735), .B(top_core_KE_n1925), .Y(top_core_KE_n1191) );
  XNOR2X1 U20491 ( .A(n6792), .B(top_core_KE_n1951), .Y(top_core_KE_n1282) );
  XNOR2X1 U20492 ( .A(n6369), .B(top_core_KE_n1967), .Y(top_core_KE_n1338) );
  XNOR2X1 U20493 ( .A(n6787), .B(top_core_KE_n1945), .Y(top_core_KE_n1261) );
  XNOR2X1 U20494 ( .A(n6361), .B(top_core_KE_n1961), .Y(top_core_KE_n1317) );
  XNOR2X1 U20495 ( .A(n6728), .B(top_core_KE_n1935), .Y(top_core_KE_n1226) );
  XNOR2X1 U20496 ( .A(n6722), .B(top_core_KE_n1929), .Y(top_core_KE_n1205) );
  MX2X1 U20497 ( .A(top_core_KE_r343_u_div_PartRem_1__1_), .B(
        top_core_KE_r343_u_div_SumTmp_0__1_), .S0(n7009), .Y(top_core_KE_N1)
         );
  XOR2X1 U20498 ( .A(top_core_KE_round_ctr_reg_0_), .B(
        top_core_KE_r343_u_div_PartRem_1__1_), .Y(
        top_core_KE_r343_u_div_SumTmp_0__1_) );
  XNOR2X1 U20499 ( .A(n6347), .B(top_core_KE_n1959), .Y(top_core_KE_n1310) );
  XNOR2X1 U20500 ( .A(n6797), .B(top_core_KE_n1955), .Y(top_core_KE_n1296) );
  XNOR2X1 U20501 ( .A(n6355), .B(top_core_KE_n1971), .Y(top_core_KE_n1352) );
  XNOR2X1 U20502 ( .A(n6795), .B(top_core_KE_n1953), .Y(top_core_KE_n1289) );
  XNOR2X1 U20503 ( .A(n6374), .B(top_core_KE_n1969), .Y(top_core_KE_n1345) );
  XNOR2X1 U20504 ( .A(n6790), .B(top_core_KE_n1949), .Y(top_core_KE_n1275) );
  XNOR2X1 U20505 ( .A(n6365), .B(top_core_KE_n1965), .Y(top_core_KE_n1331) );
  XNOR2X1 U20506 ( .A(n6788), .B(top_core_KE_n1947), .Y(top_core_KE_n1268) );
  XNOR2X1 U20507 ( .A(n6351), .B(top_core_KE_n1963), .Y(top_core_KE_n1324) );
  XNOR2X1 U20508 ( .A(n6786), .B(top_core_KE_n1943), .Y(top_core_KE_n1254) );
  XNOR2X1 U20509 ( .A(n6721), .B(top_core_KE_n1927), .Y(top_core_KE_n1198) );
  XNOR2X1 U20510 ( .A(n6739), .B(top_core_KE_n1939), .Y(top_core_KE_n1240) );
  XNOR2X1 U20511 ( .A(n6736), .B(top_core_KE_n1937), .Y(top_core_KE_n1233) );
  XNOR2X1 U20512 ( .A(n6732), .B(top_core_KE_n1933), .Y(top_core_KE_n1219) );
  XNOR2X1 U20513 ( .A(n6725), .B(top_core_KE_n1931), .Y(top_core_KE_n1212) );
  XNOR2X1 U20514 ( .A(n1334), .B(top_core_KE_n2729), .Y(top_core_KE_n2723) );
  AOI21X1 U20515 ( .A0(n7023), .A1(n7022), .B0(n7019), .Y(top_core_KE_n2729)
         );
  XNOR2X1 U20516 ( .A(top_core_KE_new_sboxw_23_), .B(top_core_KE_n2599), .Y(
        top_core_KE_n1677) );
  XNOR2X1 U20517 ( .A(top_core_KE_new_sboxw_21_), .B(top_core_KE_n2607), .Y(
        top_core_KE_n1693) );
  XNOR2X1 U20518 ( .A(top_core_KE_new_sboxw_18_), .B(top_core_KE_n2619), .Y(
        top_core_KE_n1717) );
  MXI2X1 U20519 ( .A(top_core_KE_n728), .B(top_core_KE_round_ctr_reg_0_), .S0(
        n7009), .Y(top_core_KE_N0) );
  AOI22X1 U20520 ( .A0(n625), .A1(n11712), .B0(n6731), .B1(n11786), .Y(n11785)
         );
  NAND4X1 U20521 ( .A(n11787), .B(n6922), .C(n11788), .D(n11789), .Y(n11786)
         );
  AOI22X1 U20522 ( .A0(n626), .A1(top_core_KE_sb1_n138), .B0(n6794), .B1(
        top_core_KE_sb1_n214), .Y(top_core_KE_sb1_n213) );
  NAND4X1 U20523 ( .A(top_core_KE_sb1_n215), .B(n6876), .C(
        top_core_KE_sb1_n216), .D(top_core_KE_sb1_n217), .Y(
        top_core_KE_sb1_n214) );
  AOI22X1 U20524 ( .A0(n627), .A1(n12343), .B0(n6439), .B1(n12417), .Y(n12416)
         );
  NAND4X1 U20525 ( .A(n12418), .B(n6629), .C(n12419), .D(n12420), .Y(n12417)
         );
  AOI22X1 U20526 ( .A0(n628), .A1(n12028), .B0(n6495), .B1(n12102), .Y(n12101)
         );
  NAND4X1 U20527 ( .A(n12103), .B(n6582), .C(n12104), .D(n12105), .Y(n12102)
         );
  XNOR2X1 U20528 ( .A(top_core_KE_new_sboxw_14_), .B(top_core_KE_n2635), .Y(
        top_core_KE_n1749) );
  XNOR2X1 U20529 ( .A(top_core_KE_new_sboxw_8_), .B(top_core_KE_n2659), .Y(
        top_core_KE_n1797) );
  XNOR2X1 U20530 ( .A(top_core_KE_new_sboxw_6_), .B(top_core_KE_n2667), .Y(
        top_core_KE_n1813) );
  XNOR2X1 U20531 ( .A(top_core_KE_new_sboxw_0_), .B(top_core_KE_n2691), .Y(
        top_core_KE_n1861) );
  XNOR2X1 U20532 ( .A(top_core_KE_new_sboxw_30_), .B(top_core_KE_n2564), .Y(
        top_core_KE_n1621) );
  XNOR2X1 U20533 ( .A(top_core_KE_new_sboxw_24_), .B(top_core_KE_n2594), .Y(
        top_core_KE_n1669) );
  XNOR2X1 U20534 ( .A(top_core_KE_new_sboxw_9_), .B(top_core_KE_n2655), .Y(
        top_core_KE_n1789) );
  XNOR2X1 U20535 ( .A(top_core_KE_new_sboxw_1_), .B(top_core_KE_n2687), .Y(
        top_core_KE_n1853) );
  XNOR2X1 U20536 ( .A(top_core_KE_new_sboxw_25_), .B(top_core_KE_n2589), .Y(
        top_core_KE_n1661) );
  XNOR2X1 U20537 ( .A(top_core_KE_new_sboxw_12_), .B(top_core_KE_n2643), .Y(
        top_core_KE_n1765) );
  XNOR2X1 U20538 ( .A(top_core_KE_new_sboxw_11_), .B(top_core_KE_n2647), .Y(
        top_core_KE_n1773) );
  XNOR2X1 U20539 ( .A(top_core_KE_new_sboxw_4_), .B(top_core_KE_n2675), .Y(
        top_core_KE_n1829) );
  XNOR2X1 U20540 ( .A(top_core_KE_new_sboxw_3_), .B(top_core_KE_n2679), .Y(
        top_core_KE_n1837) );
  XNOR2X1 U20541 ( .A(top_core_KE_new_sboxw_28_), .B(top_core_KE_n2574), .Y(
        top_core_KE_n1637) );
  XNOR2X1 U20542 ( .A(top_core_KE_new_sboxw_27_), .B(top_core_KE_n2579), .Y(
        top_core_KE_n1645) );
  XNOR2X1 U20543 ( .A(top_core_KE_n2183), .B(top_core_KE_n2559), .Y(
        top_core_KE_n1615) );
  XNOR2X1 U20544 ( .A(n6735), .B(top_core_KE_n2599), .Y(top_core_KE_n1679) );
  XNOR2X1 U20545 ( .A(n6722), .B(top_core_KE_n2607), .Y(top_core_KE_n1695) );
  XNOR2X1 U20546 ( .A(n6728), .B(top_core_KE_n2619), .Y(top_core_KE_n1719) );
  XNOR2X1 U20547 ( .A(n6785), .B(top_core_KE_n2631), .Y(top_core_KE_n1743) );
  XNOR2X1 U20548 ( .A(n6787), .B(top_core_KE_n2639), .Y(top_core_KE_n1759) );
  XNOR2X1 U20549 ( .A(n6792), .B(top_core_KE_n2651), .Y(top_core_KE_n1783) );
  XNOR2X1 U20550 ( .A(n6359), .B(top_core_KE_n2663), .Y(top_core_KE_n1807) );
  XNOR2X1 U20551 ( .A(n6361), .B(top_core_KE_n2671), .Y(top_core_KE_n1823) );
  XNOR2X1 U20552 ( .A(n6369), .B(top_core_KE_n2683), .Y(top_core_KE_n1847) );
  AOI22X1 U20553 ( .A0(n11695), .A1(n11790), .B0(n1354), .B1(n11791), .Y(
        n11784) );
  OAI221XL U20554 ( .A0(n1222), .A1(n185), .B0(n1223), .B1(n50), .C0(n11800), 
        .Y(n11790) );
  OAI222XL U20555 ( .A0(n1798), .A1(n11792), .B0(n11793), .B1(n11674), .C0(
        n11794), .C1(n1795), .Y(n11791) );
  AOI211X1 U20556 ( .A0(n11704), .A1(n1803), .B0(n1202), .C0(n11664), .Y(
        n11800) );
  AOI22X1 U20557 ( .A0(top_core_KE_sb1_n120), .A1(top_core_KE_sb1_n218), .B0(
        n1343), .B1(top_core_KE_sb1_n219), .Y(top_core_KE_sb1_n212) );
  OAI221XL U20558 ( .A0(n1216), .A1(n186), .B0(n1217), .B1(n51), .C0(
        top_core_KE_sb1_n228), .Y(top_core_KE_sb1_n218) );
  OAI222XL U20559 ( .A0(n1819), .A1(top_core_KE_sb1_n220), .B0(
        top_core_KE_sb1_n221), .B1(top_core_KE_sb1_n99), .C0(
        top_core_KE_sb1_n222), .C1(n1816), .Y(top_core_KE_sb1_n219) );
  AOI211X1 U20560 ( .A0(top_core_KE_sb1_n129), .A1(n1824), .B0(n1193), .C0(
        top_core_KE_sb1_n89), .Y(top_core_KE_sb1_n228) );
  AOI22X1 U20561 ( .A0(n12326), .A1(n12421), .B0(n1368), .B1(n12422), .Y(
        n12415) );
  OAI221XL U20562 ( .A0(n1181), .A1(n46), .B0(n1182), .B1(n89), .C0(n12431), 
        .Y(n12421) );
  OAI222XL U20563 ( .A0(n1756), .A1(n12423), .B0(n12424), .B1(n12305), .C0(
        n12425), .C1(n1752), .Y(n12422) );
  AOI211X1 U20564 ( .A0(n12335), .A1(n1761), .B0(n1162), .C0(n12295), .Y(
        n12431) );
  AOI22X1 U20565 ( .A0(n13272), .A1(n13366), .B0(n1356), .B1(n13367), .Y(
        n13360) );
  OAI221XL U20566 ( .A0(n1173), .A1(n187), .B0(n602), .B1(n52), .C0(n13376), 
        .Y(n13366) );
  OAI222XL U20567 ( .A0(n1666), .A1(n13368), .B0(n13369), .B1(n13251), .C0(
        n13370), .C1(n1665), .Y(n13367) );
  AOI211X1 U20568 ( .A0(n13281), .A1(n1681), .B0(n1148), .C0(n13241), .Y(
        n13376) );
  AOI22X1 U20569 ( .A0(n12011), .A1(n12106), .B0(n1357), .B1(n12107), .Y(
        n12100) );
  OAI221XL U20570 ( .A0(n1176), .A1(n188), .B0(n1177), .B1(n53), .C0(n12116), 
        .Y(n12106) );
  OAI222XL U20571 ( .A0(n1777), .A1(n12108), .B0(n12109), .B1(n11990), .C0(
        n12110), .C1(n1774), .Y(n12107) );
  AOI211X1 U20572 ( .A0(n12020), .A1(n1782), .B0(n1153), .C0(n11980), .Y(
        n12116) );
  AOI22X1 U20573 ( .A0(n12642), .A1(n12736), .B0(n1342), .B1(n12737), .Y(
        n12730) );
  OAI221XL U20574 ( .A0(n1213), .A1(n189), .B0(n603), .B1(n54), .C0(n12746), 
        .Y(n12736) );
  OAI222XL U20575 ( .A0(n1724), .A1(n12738), .B0(n12739), .B1(n12621), .C0(
        n12740), .C1(n1723), .Y(n12737) );
  AOI211X1 U20576 ( .A0(n12651), .A1(n1739), .B0(n1188), .C0(n12611), .Y(
        n12746) );
  AOI22X1 U20577 ( .A0(n13587), .A1(n13681), .B0(n1369), .B1(n13682), .Y(
        n13675) );
  OAI221XL U20578 ( .A0(n1178), .A1(n190), .B0(n609), .B1(n55), .C0(n13691), 
        .Y(n13681) );
  OAI222XL U20579 ( .A0(n1638), .A1(n13683), .B0(n13684), .B1(n13566), .C0(
        n13685), .C1(n1635), .Y(n13682) );
  AOI211X1 U20580 ( .A0(n13596), .A1(n1652), .B0(n1157), .C0(n13556), .Y(
        n13691) );
  AOI22X1 U20581 ( .A0(n12957), .A1(n13051), .B0(n1355), .B1(n13052), .Y(
        n13045) );
  OAI221XL U20582 ( .A0(n1219), .A1(n191), .B0(n604), .B1(n56), .C0(n13061), 
        .Y(n13051) );
  OAI222XL U20583 ( .A0(n1695), .A1(n13053), .B0(n13054), .B1(n12936), .C0(
        n13055), .C1(n1694), .Y(n13052) );
  AOI211X1 U20584 ( .A0(n12966), .A1(n1710), .B0(n1197), .C0(n12926), .Y(
        n13061) );
  XNOR2X1 U20585 ( .A(top_core_KE_n2517), .B(top_core_KE_n2569), .Y(
        top_core_KE_n1631) );
  XNOR2X1 U20586 ( .A(top_core_KE_n2526), .B(top_core_KE_n2584), .Y(
        top_core_KE_n1655) );
  XNOR2X1 U20587 ( .A(top_core_KE_n2514), .B(top_core_KE_n2564), .Y(
        top_core_KE_n1623) );
  XNOR2X1 U20588 ( .A(top_core_KE_n2520), .B(top_core_KE_n2574), .Y(
        top_core_KE_n1639) );
  XNOR2X1 U20589 ( .A(top_core_KE_n2523), .B(top_core_KE_n2579), .Y(
        top_core_KE_n1647) );
  XNOR2X1 U20590 ( .A(top_core_KE_n2529), .B(top_core_KE_n2589), .Y(
        top_core_KE_n1663) );
  XNOR2X1 U20591 ( .A(top_core_KE_n2532), .B(top_core_KE_n2594), .Y(
        top_core_KE_n1671) );
  XNOR2X1 U20592 ( .A(n6721), .B(top_core_KE_n2603), .Y(top_core_KE_n1687) );
  XNOR2X1 U20593 ( .A(n6739), .B(top_core_KE_n2627), .Y(top_core_KE_n1735) );
  XNOR2X1 U20594 ( .A(n6786), .B(top_core_KE_n2635), .Y(top_core_KE_n1751) );
  XNOR2X1 U20595 ( .A(n6797), .B(top_core_KE_n2659), .Y(top_core_KE_n1799) );
  XNOR2X1 U20596 ( .A(n6347), .B(top_core_KE_n2667), .Y(top_core_KE_n1815) );
  XNOR2X1 U20597 ( .A(n6355), .B(top_core_KE_n2691), .Y(top_core_KE_n1863) );
  XNOR2X1 U20598 ( .A(n6725), .B(top_core_KE_n2611), .Y(top_core_KE_n1703) );
  XNOR2X1 U20599 ( .A(n6732), .B(top_core_KE_n2615), .Y(top_core_KE_n1711) );
  XNOR2X1 U20600 ( .A(n6736), .B(top_core_KE_n2623), .Y(top_core_KE_n1727) );
  XNOR2X1 U20601 ( .A(n6788), .B(top_core_KE_n2643), .Y(top_core_KE_n1767) );
  XNOR2X1 U20602 ( .A(n6790), .B(top_core_KE_n2647), .Y(top_core_KE_n1775) );
  XNOR2X1 U20603 ( .A(n6795), .B(top_core_KE_n2655), .Y(top_core_KE_n1791) );
  XNOR2X1 U20604 ( .A(n6351), .B(top_core_KE_n2675), .Y(top_core_KE_n1831) );
  XNOR2X1 U20605 ( .A(n6365), .B(top_core_KE_n2679), .Y(top_core_KE_n1839) );
  XNOR2X1 U20606 ( .A(n6374), .B(top_core_KE_n2687), .Y(top_core_KE_n1855) );
  XOR2X1 U20607 ( .A(top_core_KE_n2380), .B(n6496), .Y(top_core_KE_n1179) );
  XOR2X1 U20608 ( .A(top_core_KE_n2344), .B(n6483), .Y(top_core_KE_n1137) );
  XOR2X1 U20609 ( .A(top_core_KE_n2386), .B(n6499), .Y(top_core_KE_n1186) );
  XOR2X1 U20610 ( .A(top_core_KE_n2374), .B(n6492), .Y(top_core_KE_n1172) );
  XOR2X1 U20611 ( .A(top_core_KE_n2368), .B(n6489), .Y(top_core_KE_n1165) );
  XOR2X1 U20612 ( .A(top_core_KE_n2362), .B(n6486), .Y(top_core_KE_n1158) );
  XOR2X1 U20613 ( .A(top_core_KE_n2356), .B(n6485), .Y(top_core_KE_n1151) );
  XOR2X1 U20614 ( .A(top_core_KE_n2350), .B(n6484), .Y(top_core_KE_n1144) );
  XNOR2X1 U20615 ( .A(top_core_KE_new_sboxw_22_), .B(top_core_KE_n2603), .Y(
        top_core_KE_n1685) );
  XNOR2X1 U20616 ( .A(top_core_KE_new_sboxw_16_), .B(top_core_KE_n2627), .Y(
        top_core_KE_n1733) );
  XNOR2X1 U20617 ( .A(n6696), .B(n6499), .Y(top_core_KE_n962) );
  XNOR2X1 U20618 ( .A(n6675), .B(n6492), .Y(top_core_KE_n948) );
  XNOR2X1 U20619 ( .A(n6656), .B(n6489), .Y(top_core_KE_n941) );
  XNOR2X1 U20620 ( .A(n6608), .B(n6486), .Y(top_core_KE_n934) );
  XNOR2X1 U20621 ( .A(n6525), .B(n6485), .Y(top_core_KE_n927) );
  XNOR2X1 U20622 ( .A(n6437), .B(n6484), .Y(top_core_KE_n920) );
  XNOR2X1 U20623 ( .A(n6344), .B(n6483), .Y(top_core_KE_n909) );
  XNOR2X1 U20624 ( .A(n6317), .B(n6496), .Y(top_core_KE_n955) );
  XNOR2X1 U20625 ( .A(top_core_KE_new_sboxw_17_), .B(top_core_KE_n2623), .Y(
        top_core_KE_n1725) );
  XNOR2X1 U20626 ( .A(top_core_KE_new_sboxw_20_), .B(top_core_KE_n2611), .Y(
        top_core_KE_n1701) );
  XNOR2X1 U20627 ( .A(top_core_KE_new_sboxw_19_), .B(top_core_KE_n2615), .Y(
        top_core_KE_n1709) );
  XOR2X1 U20628 ( .A(top_core_KE_new_sboxw_7_), .B(top_core_KE_n1957), .Y(
        top_core_KE_n1301) );
  XOR2X1 U20629 ( .A(top_core_KE_new_sboxw_15_), .B(top_core_KE_n1941), .Y(
        top_core_KE_n1245) );
  XOR2X1 U20630 ( .A(top_core_KE_new_sboxw_10_), .B(top_core_KE_n1951), .Y(
        top_core_KE_n1280) );
  XOR2X1 U20631 ( .A(top_core_KE_new_sboxw_2_), .B(top_core_KE_n1967), .Y(
        top_core_KE_n1336) );
  XOR2X1 U20632 ( .A(top_core_KE_new_sboxw_13_), .B(top_core_KE_n1945), .Y(
        top_core_KE_n1259) );
  XOR2X1 U20633 ( .A(top_core_KE_new_sboxw_5_), .B(top_core_KE_n1961), .Y(
        top_core_KE_n1315) );
  BUFX3 U20634 ( .A(top_core_KE_n745), .Y(n1372) );
  OAI21XL U20635 ( .A0(top_core_KE_n898), .A1(top_core_KE_n899), .B0(n2143), 
        .Y(top_core_KE_n745) );
  OAI221XL U20636 ( .A0(n6342), .A1(top_core_KE_n900), .B0(n6341), .B1(n2228), 
        .C0(top_core_KE_n901), .Y(top_core_KE_n899) );
  OAI221XL U20637 ( .A0(n2149), .A1(n6337), .B0(n2157), .B1(n7245), .C0(
        top_core_KE_n906), .Y(top_core_KE_n898) );
  BUFX3 U20638 ( .A(top_core_KE_n746), .Y(n1373) );
  OAI21XL U20639 ( .A0(top_core_KE_n911), .A1(top_core_KE_n912), .B0(n2138), 
        .Y(top_core_KE_n746) );
  OAI221XL U20640 ( .A0(top_core_KE_n913), .A1(n2193), .B0(top_core_KE_n915), 
        .B1(n7117), .C0(top_core_KE_n916), .Y(top_core_KE_n912) );
  OAI221XL U20641 ( .A0(n2145), .A1(n6405), .B0(n2153), .B1(n7244), .C0(
        top_core_KE_n919), .Y(top_core_KE_n911) );
  BUFX3 U20642 ( .A(top_core_KE_n747), .Y(n1374) );
  OAI21XL U20643 ( .A0(top_core_KE_n921), .A1(top_core_KE_n922), .B0(n2139), 
        .Y(top_core_KE_n747) );
  OAI221XL U20644 ( .A0(top_core_KE_n923), .A1(n2190), .B0(n2208), .B1(n7116), 
        .C0(top_core_KE_n924), .Y(top_core_KE_n922) );
  OAI221XL U20645 ( .A0(n2145), .A1(n6513), .B0(n2153), .B1(n7243), .C0(
        top_core_KE_n926), .Y(top_core_KE_n921) );
  BUFX3 U20646 ( .A(top_core_KE_n748), .Y(n1375) );
  OAI21XL U20647 ( .A0(top_core_KE_n928), .A1(top_core_KE_n929), .B0(n2140), 
        .Y(top_core_KE_n748) );
  OAI221XL U20648 ( .A0(top_core_KE_n930), .A1(n2190), .B0(n2207), .B1(n7115), 
        .C0(top_core_KE_n931), .Y(top_core_KE_n929) );
  OAI221XL U20649 ( .A0(n2145), .A1(n6583), .B0(n2153), .B1(n7242), .C0(
        top_core_KE_n933), .Y(top_core_KE_n928) );
  BUFX3 U20650 ( .A(top_core_KE_n749), .Y(n1376) );
  OAI21XL U20651 ( .A0(top_core_KE_n935), .A1(top_core_KE_n936), .B0(n2137), 
        .Y(top_core_KE_n749) );
  OAI221XL U20652 ( .A0(top_core_KE_n937), .A1(n2190), .B0(n2205), .B1(n7114), 
        .C0(top_core_KE_n938), .Y(top_core_KE_n936) );
  OAI221XL U20653 ( .A0(n2145), .A1(n6647), .B0(n2153), .B1(n7241), .C0(
        top_core_KE_n940), .Y(top_core_KE_n935) );
  BUFX3 U20654 ( .A(top_core_KE_n750), .Y(n1377) );
  OAI21XL U20655 ( .A0(top_core_KE_n942), .A1(top_core_KE_n943), .B0(n2143), 
        .Y(top_core_KE_n750) );
  OAI221XL U20656 ( .A0(top_core_KE_n944), .A1(n2190), .B0(n2210), .B1(n7113), 
        .C0(top_core_KE_n945), .Y(top_core_KE_n943) );
  OAI221XL U20657 ( .A0(n2145), .A1(n6671), .B0(n2153), .B1(n7240), .C0(
        top_core_KE_n947), .Y(top_core_KE_n942) );
  BUFX3 U20658 ( .A(top_core_KE_n751), .Y(n1378) );
  OAI21XL U20659 ( .A0(top_core_KE_n949), .A1(top_core_KE_n950), .B0(n2138), 
        .Y(top_core_KE_n751) );
  OAI221XL U20660 ( .A0(top_core_KE_n951), .A1(n2190), .B0(n2209), .B1(n7112), 
        .C0(top_core_KE_n952), .Y(top_core_KE_n950) );
  OAI221XL U20661 ( .A0(n2145), .A1(n6310), .B0(n2153), .B1(n7239), .C0(
        top_core_KE_n954), .Y(top_core_KE_n949) );
  BUFX3 U20662 ( .A(top_core_KE_n752), .Y(n1379) );
  OAI21XL U20663 ( .A0(top_core_KE_n956), .A1(top_core_KE_n957), .B0(n2139), 
        .Y(top_core_KE_n752) );
  OAI221XL U20664 ( .A0(top_core_KE_n958), .A1(n2190), .B0(n2208), .B1(n7111), 
        .C0(top_core_KE_n959), .Y(top_core_KE_n957) );
  OAI221XL U20665 ( .A0(n2145), .A1(n6692), .B0(n2153), .B1(n7238), .C0(
        top_core_KE_n961), .Y(top_core_KE_n956) );
  BUFX3 U20666 ( .A(top_core_KE_n761), .Y(n1388) );
  OAI21XL U20667 ( .A0(top_core_KE_n1019), .A1(top_core_KE_n1020), .B0(n2141), 
        .Y(top_core_KE_n761) );
  OAI221XL U20668 ( .A0(top_core_KE_n1021), .A1(n2190), .B0(n2208), .B1(n7110), 
        .C0(top_core_KE_n1022), .Y(top_core_KE_n1020) );
  OAI221XL U20669 ( .A0(n2146), .A1(n6323), .B0(n2154), .B1(n7229), .C0(
        top_core_KE_n1024), .Y(top_core_KE_n1019) );
  BUFX3 U20670 ( .A(top_core_KE_n762), .Y(n1389) );
  OAI21XL U20671 ( .A0(top_core_KE_n1026), .A1(top_core_KE_n1027), .B0(n2144), 
        .Y(top_core_KE_n762) );
  OAI221XL U20672 ( .A0(top_core_KE_n1028), .A1(n2190), .B0(n2207), .B1(n7109), 
        .C0(top_core_KE_n1029), .Y(top_core_KE_n1027) );
  OAI221XL U20673 ( .A0(n2146), .A1(n6388), .B0(n2154), .B1(n7228), .C0(
        top_core_KE_n1031), .Y(top_core_KE_n1026) );
  BUFX3 U20674 ( .A(top_core_KE_n763), .Y(n1390) );
  OAI21XL U20675 ( .A0(top_core_KE_n1033), .A1(top_core_KE_n1034), .B0(n2137), 
        .Y(top_core_KE_n763) );
  OAI221XL U20676 ( .A0(top_core_KE_n1035), .A1(n2190), .B0(n2205), .B1(n7108), 
        .C0(top_core_KE_n1036), .Y(top_core_KE_n1034) );
  OAI221XL U20677 ( .A0(n2146), .A1(n6810), .B0(n2154), .B1(n7227), .C0(
        top_core_KE_n1038), .Y(top_core_KE_n1033) );
  BUFX3 U20678 ( .A(top_core_KE_n764), .Y(n1391) );
  OAI21XL U20679 ( .A0(top_core_KE_n1040), .A1(top_core_KE_n1041), .B0(n2138), 
        .Y(top_core_KE_n764) );
  OAI221XL U20680 ( .A0(top_core_KE_n1042), .A1(n2190), .B0(n2210), .B1(n7107), 
        .C0(top_core_KE_n1043), .Y(top_core_KE_n1041) );
  OAI221XL U20681 ( .A0(n2146), .A1(n6877), .B0(n2154), .B1(n7226), .C0(
        top_core_KE_n1045), .Y(top_core_KE_n1040) );
  BUFX3 U20682 ( .A(top_core_KE_n765), .Y(n1392) );
  OAI21XL U20683 ( .A0(top_core_KE_n1047), .A1(top_core_KE_n1048), .B0(n2139), 
        .Y(top_core_KE_n765) );
  OAI221XL U20684 ( .A0(top_core_KE_n1049), .A1(n2190), .B0(n2210), .B1(n7106), 
        .C0(top_core_KE_n1050), .Y(top_core_KE_n1048) );
  OAI221XL U20685 ( .A0(n2146), .A1(n6938), .B0(n2154), .B1(n7225), .C0(
        top_core_KE_n1052), .Y(top_core_KE_n1047) );
  BUFX3 U20686 ( .A(top_core_KE_n766), .Y(n1393) );
  OAI21XL U20687 ( .A0(top_core_KE_n1054), .A1(top_core_KE_n1055), .B0(n2137), 
        .Y(top_core_KE_n766) );
  OAI221XL U20688 ( .A0(top_core_KE_n1056), .A1(n2191), .B0(n2210), .B1(n7105), 
        .C0(top_core_KE_n1057), .Y(top_core_KE_n1055) );
  OAI221XL U20689 ( .A0(n2146), .A1(n6959), .B0(n2154), .B1(n7224), .C0(
        top_core_KE_n1059), .Y(top_core_KE_n1054) );
  BUFX3 U20690 ( .A(top_core_KE_n767), .Y(n1394) );
  OAI21XL U20691 ( .A0(top_core_KE_n1061), .A1(top_core_KE_n1062), .B0(n2137), 
        .Y(top_core_KE_n767) );
  OAI221XL U20692 ( .A0(top_core_KE_n1063), .A1(n2191), .B0(n2210), .B1(n7104), 
        .C0(top_core_KE_n1064), .Y(top_core_KE_n1062) );
  OAI221XL U20693 ( .A0(n2146), .A1(n6970), .B0(n2154), .B1(n7223), .C0(
        top_core_KE_n1066), .Y(top_core_KE_n1061) );
  BUFX3 U20694 ( .A(top_core_KE_n768), .Y(n1395) );
  OAI21XL U20695 ( .A0(top_core_KE_n1068), .A1(top_core_KE_n1069), .B0(n2137), 
        .Y(top_core_KE_n768) );
  OAI221XL U20696 ( .A0(top_core_KE_n1070), .A1(n2191), .B0(n2210), .B1(n7103), 
        .C0(top_core_KE_n1071), .Y(top_core_KE_n1069) );
  OAI221XL U20697 ( .A0(n2146), .A1(n6980), .B0(n2154), .B1(n7222), .C0(
        top_core_KE_n1073), .Y(top_core_KE_n1068) );
  BUFX3 U20698 ( .A(top_core_KE_n769), .Y(n1396) );
  OAI21XL U20699 ( .A0(top_core_KE_n1075), .A1(top_core_KE_n1076), .B0(n2137), 
        .Y(top_core_KE_n769) );
  OAI221XL U20700 ( .A0(top_core_KE_n1077), .A1(n2191), .B0(n2210), .B1(n7102), 
        .C0(top_core_KE_n1078), .Y(top_core_KE_n1076) );
  OAI221XL U20701 ( .A0(n2148), .A1(n6319), .B0(n2155), .B1(n7221), .C0(
        top_core_KE_n1080), .Y(top_core_KE_n1075) );
  BUFX3 U20702 ( .A(top_core_KE_n770), .Y(n1397) );
  OAI21XL U20703 ( .A0(top_core_KE_n1082), .A1(top_core_KE_n1083), .B0(n2137), 
        .Y(top_core_KE_n770) );
  OAI221XL U20704 ( .A0(top_core_KE_n1084), .A1(n2191), .B0(n2210), .B1(n7101), 
        .C0(top_core_KE_n1085), .Y(top_core_KE_n1083) );
  OAI221XL U20705 ( .A0(n2149), .A1(n6380), .B0(n2155), .B1(n7220), .C0(
        top_core_KE_n1087), .Y(top_core_KE_n1082) );
  BUFX3 U20706 ( .A(top_core_KE_n771), .Y(n1398) );
  OAI21XL U20707 ( .A0(top_core_KE_n1089), .A1(top_core_KE_n1090), .B0(n2137), 
        .Y(top_core_KE_n771) );
  OAI221XL U20708 ( .A0(top_core_KE_n1091), .A1(n2191), .B0(n2210), .B1(n7100), 
        .C0(top_core_KE_n1092), .Y(top_core_KE_n1090) );
  OAI221XL U20709 ( .A0(n2145), .A1(n6747), .B0(n2155), .B1(n7219), .C0(
        top_core_KE_n1094), .Y(top_core_KE_n1089) );
  BUFX3 U20710 ( .A(top_core_KE_n772), .Y(n1399) );
  OAI21XL U20711 ( .A0(top_core_KE_n1096), .A1(top_core_KE_n1097), .B0(n2137), 
        .Y(top_core_KE_n772) );
  OAI221XL U20712 ( .A0(top_core_KE_n1098), .A1(n2191), .B0(n2210), .B1(n7099), 
        .C0(top_core_KE_n1099), .Y(top_core_KE_n1097) );
  OAI221XL U20713 ( .A0(n2147), .A1(n6831), .B0(n2155), .B1(n7218), .C0(
        top_core_KE_n1101), .Y(top_core_KE_n1096) );
  BUFX3 U20714 ( .A(top_core_KE_n773), .Y(n1400) );
  OAI21XL U20715 ( .A0(top_core_KE_n1103), .A1(top_core_KE_n1104), .B0(n2137), 
        .Y(top_core_KE_n773) );
  OAI221XL U20716 ( .A0(top_core_KE_n1105), .A1(n2191), .B0(n2210), .B1(n7098), 
        .C0(top_core_KE_n1106), .Y(top_core_KE_n1104) );
  OAI221XL U20717 ( .A0(n2152), .A1(n6923), .B0(n2155), .B1(n7217), .C0(
        top_core_KE_n1108), .Y(top_core_KE_n1103) );
  BUFX3 U20718 ( .A(top_core_KE_n774), .Y(n1401) );
  OAI21XL U20719 ( .A0(top_core_KE_n1110), .A1(top_core_KE_n1111), .B0(n2137), 
        .Y(top_core_KE_n774) );
  OAI221XL U20720 ( .A0(top_core_KE_n1112), .A1(n2191), .B0(n2210), .B1(n7097), 
        .C0(top_core_KE_n1113), .Y(top_core_KE_n1111) );
  OAI221XL U20721 ( .A0(n2150), .A1(n6953), .B0(n2155), .B1(n7216), .C0(
        top_core_KE_n1115), .Y(top_core_KE_n1110) );
  BUFX3 U20722 ( .A(top_core_KE_n775), .Y(n1402) );
  OAI21XL U20723 ( .A0(top_core_KE_n1117), .A1(top_core_KE_n1118), .B0(n2137), 
        .Y(top_core_KE_n775) );
  OAI221XL U20724 ( .A0(top_core_KE_n1119), .A1(n2191), .B0(n2210), .B1(n7096), 
        .C0(top_core_KE_n1120), .Y(top_core_KE_n1118) );
  OAI221XL U20725 ( .A0(n2146), .A1(n6965), .B0(n2155), .B1(n7215), .C0(
        top_core_KE_n1122), .Y(top_core_KE_n1117) );
  BUFX3 U20726 ( .A(top_core_KE_n776), .Y(n1403) );
  OAI21XL U20727 ( .A0(top_core_KE_n1124), .A1(top_core_KE_n1125), .B0(n2140), 
        .Y(top_core_KE_n776) );
  OAI221XL U20728 ( .A0(top_core_KE_n1126), .A1(n2191), .B0(n2209), .B1(n7095), 
        .C0(top_core_KE_n1127), .Y(top_core_KE_n1125) );
  OAI221XL U20729 ( .A0(n2151), .A1(n6975), .B0(n2155), .B1(n7214), .C0(
        top_core_KE_n1129), .Y(top_core_KE_n1124) );
  BUFX3 U20730 ( .A(top_core_KE_n777), .Y(n1404) );
  OAI21XL U20731 ( .A0(top_core_KE_n1131), .A1(top_core_KE_n1132), .B0(n2137), 
        .Y(top_core_KE_n777) );
  OAI221XL U20732 ( .A0(top_core_KE_n1133), .A1(n2191), .B0(n2209), .B1(n7094), 
        .C0(top_core_KE_n1134), .Y(top_core_KE_n1132) );
  OAI221XL U20733 ( .A0(n2148), .A1(n6345), .B0(n2155), .B1(n7213), .C0(
        top_core_KE_n1136), .Y(top_core_KE_n1131) );
  BUFX3 U20734 ( .A(top_core_KE_n778), .Y(n1405) );
  OAI21XL U20735 ( .A0(top_core_KE_n1138), .A1(top_core_KE_n1139), .B0(n2137), 
        .Y(top_core_KE_n778) );
  OAI221XL U20736 ( .A0(top_core_KE_n1140), .A1(n2192), .B0(n2209), .B1(n7093), 
        .C0(top_core_KE_n1141), .Y(top_core_KE_n1139) );
  OAI221XL U20737 ( .A0(n2149), .A1(n6438), .B0(n2155), .B1(n7212), .C0(
        top_core_KE_n1143), .Y(top_core_KE_n1138) );
  BUFX3 U20738 ( .A(top_core_KE_n779), .Y(n1406) );
  OAI21XL U20739 ( .A0(top_core_KE_n1145), .A1(top_core_KE_n1146), .B0(n2137), 
        .Y(top_core_KE_n779) );
  OAI221XL U20740 ( .A0(top_core_KE_n1147), .A1(n2192), .B0(n2209), .B1(n7092), 
        .C0(top_core_KE_n1148), .Y(top_core_KE_n1146) );
  OAI221XL U20741 ( .A0(n2145), .A1(n6526), .B0(n2155), .B1(n7211), .C0(
        top_core_KE_n1150), .Y(top_core_KE_n1145) );
  BUFX3 U20742 ( .A(top_core_KE_n780), .Y(n1407) );
  OAI21XL U20743 ( .A0(top_core_KE_n1152), .A1(top_core_KE_n1153), .B0(n2138), 
        .Y(top_core_KE_n780) );
  OAI221XL U20744 ( .A0(top_core_KE_n1154), .A1(n2192), .B0(n2209), .B1(n7091), 
        .C0(top_core_KE_n1155), .Y(top_core_KE_n1153) );
  OAI221XL U20745 ( .A0(n2147), .A1(n6609), .B0(n2155), .B1(n7210), .C0(
        top_core_KE_n1157), .Y(top_core_KE_n1152) );
  BUFX3 U20746 ( .A(top_core_KE_n781), .Y(n1408) );
  OAI21XL U20747 ( .A0(top_core_KE_n1159), .A1(top_core_KE_n1160), .B0(n2138), 
        .Y(top_core_KE_n781) );
  OAI221XL U20748 ( .A0(top_core_KE_n1161), .A1(n2192), .B0(n2209), .B1(n7090), 
        .C0(top_core_KE_n1162), .Y(top_core_KE_n1160) );
  OAI221XL U20749 ( .A0(n2147), .A1(n6657), .B0(n2156), .B1(n7209), .C0(
        top_core_KE_n1164), .Y(top_core_KE_n1159) );
  BUFX3 U20750 ( .A(top_core_KE_n782), .Y(n1409) );
  OAI21XL U20751 ( .A0(top_core_KE_n1166), .A1(top_core_KE_n1167), .B0(n2138), 
        .Y(top_core_KE_n782) );
  OAI221XL U20752 ( .A0(top_core_KE_n1168), .A1(n2192), .B0(n2209), .B1(n7089), 
        .C0(top_core_KE_n1169), .Y(top_core_KE_n1167) );
  OAI221XL U20753 ( .A0(n2147), .A1(n6676), .B0(n2156), .B1(n7208), .C0(
        top_core_KE_n1171), .Y(top_core_KE_n1166) );
  BUFX3 U20754 ( .A(top_core_KE_n783), .Y(n1410) );
  OAI21XL U20755 ( .A0(top_core_KE_n1173), .A1(top_core_KE_n1174), .B0(n2138), 
        .Y(top_core_KE_n783) );
  OAI221XL U20756 ( .A0(top_core_KE_n1175), .A1(n2192), .B0(n2209), .B1(n7088), 
        .C0(top_core_KE_n1176), .Y(top_core_KE_n1174) );
  OAI221XL U20757 ( .A0(n2147), .A1(n6318), .B0(n2156), .B1(n7207), .C0(
        top_core_KE_n1178), .Y(top_core_KE_n1173) );
  BUFX3 U20758 ( .A(top_core_KE_n784), .Y(n1411) );
  OAI21XL U20759 ( .A0(top_core_KE_n1180), .A1(top_core_KE_n1181), .B0(n2138), 
        .Y(top_core_KE_n784) );
  OAI221XL U20760 ( .A0(top_core_KE_n1182), .A1(n2192), .B0(n2209), .B1(n7087), 
        .C0(top_core_KE_n1183), .Y(top_core_KE_n1181) );
  OAI221XL U20761 ( .A0(n2147), .A1(n6697), .B0(n2156), .B1(n7206), .C0(
        top_core_KE_n1185), .Y(top_core_KE_n1180) );
  BUFX3 U20762 ( .A(top_core_KE_n809), .Y(n1436) );
  OAI21XL U20763 ( .A0(top_core_KE_n1355), .A1(top_core_KE_n1356), .B0(n2140), 
        .Y(top_core_KE_n809) );
  OAI221XL U20764 ( .A0(n6336), .A1(top_core_KE_n900), .B0(n6337), .B1(n2221), 
        .C0(top_core_KE_n1357), .Y(top_core_KE_n1356) );
  OAI221XL U20765 ( .A0(n6344), .A1(n2152), .B0(n7181), .B1(n2154), .C0(
        top_core_KE_n1360), .Y(top_core_KE_n1355) );
  BUFX3 U20766 ( .A(top_core_KE_n810), .Y(n1437) );
  OAI21XL U20767 ( .A0(top_core_KE_n1363), .A1(top_core_KE_n1364), .B0(n2140), 
        .Y(top_core_KE_n810) );
  OAI221XL U20768 ( .A0(top_core_KE_n1365), .A1(n2192), .B0(n2209), .B1(n7086), 
        .C0(top_core_KE_n1366), .Y(top_core_KE_n1364) );
  OAI221XL U20769 ( .A0(n2149), .A1(n6437), .B0(n2157), .B1(n7180), .C0(
        top_core_KE_n1368), .Y(top_core_KE_n1363) );
  BUFX3 U20770 ( .A(top_core_KE_n811), .Y(n1438) );
  OAI21XL U20771 ( .A0(top_core_KE_n1371), .A1(top_core_KE_n1372), .B0(n2140), 
        .Y(top_core_KE_n811) );
  OAI221XL U20772 ( .A0(top_core_KE_n1373), .A1(n2192), .B0(n2209), .B1(n7085), 
        .C0(top_core_KE_n1374), .Y(top_core_KE_n1372) );
  OAI221XL U20773 ( .A0(n2149), .A1(n6525), .B0(n2157), .B1(n7179), .C0(
        top_core_KE_n1376), .Y(top_core_KE_n1371) );
  BUFX3 U20774 ( .A(top_core_KE_n812), .Y(n1439) );
  OAI21XL U20775 ( .A0(top_core_KE_n1379), .A1(top_core_KE_n1380), .B0(n2140), 
        .Y(top_core_KE_n812) );
  OAI221XL U20776 ( .A0(top_core_KE_n1381), .A1(n2192), .B0(n2209), .B1(n7084), 
        .C0(top_core_KE_n1382), .Y(top_core_KE_n1380) );
  OAI221XL U20777 ( .A0(n2149), .A1(n6608), .B0(n2157), .B1(n7178), .C0(
        top_core_KE_n1384), .Y(top_core_KE_n1379) );
  BUFX3 U20778 ( .A(top_core_KE_n813), .Y(n1440) );
  OAI21XL U20779 ( .A0(top_core_KE_n1387), .A1(top_core_KE_n1388), .B0(n2140), 
        .Y(top_core_KE_n813) );
  OAI221XL U20780 ( .A0(top_core_KE_n1389), .A1(n2192), .B0(n2208), .B1(n7083), 
        .C0(top_core_KE_n1390), .Y(top_core_KE_n1388) );
  OAI221XL U20781 ( .A0(n2149), .A1(n6656), .B0(n2157), .B1(n7177), .C0(
        top_core_KE_n1392), .Y(top_core_KE_n1387) );
  BUFX3 U20782 ( .A(top_core_KE_n814), .Y(n1441) );
  OAI21XL U20783 ( .A0(top_core_KE_n1395), .A1(top_core_KE_n1396), .B0(n2140), 
        .Y(top_core_KE_n814) );
  OAI221XL U20784 ( .A0(top_core_KE_n1397), .A1(n2192), .B0(n2208), .B1(n7082), 
        .C0(top_core_KE_n1398), .Y(top_core_KE_n1396) );
  OAI221XL U20785 ( .A0(n2149), .A1(n6675), .B0(n2157), .B1(n7176), .C0(
        top_core_KE_n1400), .Y(top_core_KE_n1395) );
  BUFX3 U20786 ( .A(top_core_KE_n815), .Y(n1442) );
  OAI21XL U20787 ( .A0(top_core_KE_n1403), .A1(top_core_KE_n1404), .B0(n2140), 
        .Y(top_core_KE_n815) );
  OAI221XL U20788 ( .A0(top_core_KE_n1405), .A1(n2193), .B0(n2208), .B1(n7081), 
        .C0(top_core_KE_n1406), .Y(top_core_KE_n1404) );
  OAI221XL U20789 ( .A0(n2149), .A1(n6317), .B0(n2157), .B1(n7175), .C0(
        top_core_KE_n1408), .Y(top_core_KE_n1403) );
  BUFX3 U20790 ( .A(top_core_KE_n816), .Y(n1443) );
  OAI21XL U20791 ( .A0(top_core_KE_n1411), .A1(top_core_KE_n1412), .B0(n2140), 
        .Y(top_core_KE_n816) );
  OAI221XL U20792 ( .A0(top_core_KE_n1413), .A1(n2193), .B0(n2208), .B1(n7080), 
        .C0(top_core_KE_n1414), .Y(top_core_KE_n1412) );
  OAI221XL U20793 ( .A0(n2147), .A1(n6696), .B0(n2158), .B1(n7174), .C0(
        top_core_KE_n1416), .Y(top_core_KE_n1411) );
  BUFX3 U20794 ( .A(top_core_KE_n817), .Y(n1444) );
  OAI21XL U20795 ( .A0(top_core_KE_n1419), .A1(top_core_KE_n1420), .B0(n2140), 
        .Y(top_core_KE_n817) );
  OAI221XL U20796 ( .A0(top_core_KE_n1421), .A1(n2193), .B0(n2208), .B1(n7079), 
        .C0(top_core_KE_n1422), .Y(top_core_KE_n1420) );
  OAI221XL U20797 ( .A0(n2149), .A1(n6395), .B0(n2157), .B1(n7173), .C0(
        top_core_KE_n1424), .Y(top_core_KE_n1419) );
  BUFX3 U20798 ( .A(top_core_KE_n818), .Y(n1445) );
  OAI21XL U20799 ( .A0(top_core_KE_n1427), .A1(top_core_KE_n1428), .B0(n2141), 
        .Y(top_core_KE_n818) );
  OAI221XL U20800 ( .A0(top_core_KE_n1429), .A1(n2193), .B0(n2208), .B1(n7078), 
        .C0(top_core_KE_n1430), .Y(top_core_KE_n1428) );
  OAI221XL U20801 ( .A0(n2152), .A1(n6403), .B0(n2158), .B1(n7172), .C0(
        top_core_KE_n1432), .Y(top_core_KE_n1427) );
  BUFX3 U20802 ( .A(top_core_KE_n819), .Y(n1446) );
  OAI21XL U20803 ( .A0(top_core_KE_n1435), .A1(top_core_KE_n1436), .B0(n2141), 
        .Y(top_core_KE_n819) );
  OAI221XL U20804 ( .A0(top_core_KE_n1437), .A1(n2193), .B0(n2208), .B1(n7077), 
        .C0(top_core_KE_n1438), .Y(top_core_KE_n1436) );
  OAI221XL U20805 ( .A0(n2150), .A1(n6481), .B0(n2158), .B1(n7171), .C0(
        top_core_KE_n1440), .Y(top_core_KE_n1435) );
  BUFX3 U20806 ( .A(top_core_KE_n820), .Y(n1447) );
  OAI21XL U20807 ( .A0(top_core_KE_n1443), .A1(top_core_KE_n1444), .B0(n2141), 
        .Y(top_core_KE_n820) );
  OAI221XL U20808 ( .A0(top_core_KE_n1445), .A1(n2193), .B0(n2208), .B1(n7076), 
        .C0(top_core_KE_n1446), .Y(top_core_KE_n1444) );
  OAI221XL U20809 ( .A0(n2146), .A1(n6561), .B0(n2158), .B1(n7170), .C0(
        top_core_KE_n1448), .Y(top_core_KE_n1443) );
  BUFX3 U20810 ( .A(top_core_KE_n821), .Y(n1448) );
  OAI21XL U20811 ( .A0(top_core_KE_n1451), .A1(top_core_KE_n1452), .B0(n2141), 
        .Y(top_core_KE_n821) );
  OAI221XL U20812 ( .A0(top_core_KE_n1453), .A1(n2193), .B0(n2208), .B1(n7075), 
        .C0(top_core_KE_n1454), .Y(top_core_KE_n1452) );
  OAI221XL U20813 ( .A0(n2146), .A1(n6640), .B0(n2158), .B1(n7169), .C0(
        top_core_KE_n1456), .Y(top_core_KE_n1451) );
  BUFX3 U20814 ( .A(top_core_KE_n822), .Y(n1449) );
  OAI21XL U20815 ( .A0(top_core_KE_n1459), .A1(top_core_KE_n1460), .B0(n2141), 
        .Y(top_core_KE_n822) );
  OAI221XL U20816 ( .A0(top_core_KE_n1461), .A1(n2193), .B0(n2208), .B1(n7074), 
        .C0(top_core_KE_n1462), .Y(top_core_KE_n1460) );
  OAI221XL U20817 ( .A0(n2151), .A1(n6668), .B0(n2158), .B1(n7168), .C0(
        top_core_KE_n1464), .Y(top_core_KE_n1459) );
  BUFX3 U20818 ( .A(top_core_KE_n823), .Y(n1450) );
  OAI21XL U20819 ( .A0(top_core_KE_n1467), .A1(top_core_KE_n1468), .B0(n2141), 
        .Y(top_core_KE_n823) );
  OAI221XL U20820 ( .A0(top_core_KE_n1469), .A1(n2193), .B0(n2208), .B1(n7073), 
        .C0(top_core_KE_n1470), .Y(top_core_KE_n1468) );
  OAI221XL U20821 ( .A0(n2148), .A1(n6683), .B0(n2158), .B1(n7167), .C0(
        top_core_KE_n1472), .Y(top_core_KE_n1467) );
  BUFX3 U20822 ( .A(top_core_KE_n824), .Y(n1451) );
  OAI21XL U20823 ( .A0(top_core_KE_n1475), .A1(top_core_KE_n1476), .B0(n2141), 
        .Y(top_core_KE_n824) );
  OAI221XL U20824 ( .A0(top_core_KE_n1477), .A1(n2193), .B0(n2208), .B1(n7072), 
        .C0(top_core_KE_n1478), .Y(top_core_KE_n1476) );
  OAI221XL U20825 ( .A0(n2149), .A1(n6690), .B0(n2158), .B1(n7166), .C0(
        top_core_KE_n1480), .Y(top_core_KE_n1475) );
  BUFX3 U20826 ( .A(top_core_KE_n825), .Y(n1452) );
  OAI21XL U20827 ( .A0(top_core_KE_n1483), .A1(top_core_KE_n1484), .B0(n2141), 
        .Y(top_core_KE_n825) );
  OAI221XL U20828 ( .A0(top_core_KE_n1485), .A1(n2193), .B0(n2207), .B1(n7071), 
        .C0(top_core_KE_n1486), .Y(top_core_KE_n1484) );
  OAI221XL U20829 ( .A0(n2145), .A1(n6330), .B0(n2158), .B1(n7165), .C0(
        top_core_KE_n1488), .Y(top_core_KE_n1483) );
  BUFX3 U20830 ( .A(top_core_KE_n826), .Y(n1453) );
  OAI21XL U20831 ( .A0(top_core_KE_n1491), .A1(top_core_KE_n1492), .B0(n2141), 
        .Y(top_core_KE_n826) );
  OAI221XL U20832 ( .A0(top_core_KE_n1493), .A1(n2191), .B0(n2207), .B1(n7070), 
        .C0(top_core_KE_n1494), .Y(top_core_KE_n1492) );
  OAI221XL U20833 ( .A0(n2147), .A1(n6719), .B0(n2158), .B1(n7164), .C0(
        top_core_KE_n1496), .Y(top_core_KE_n1491) );
  BUFX3 U20834 ( .A(top_core_KE_n827), .Y(n1454) );
  OAI21XL U20835 ( .A0(top_core_KE_n1499), .A1(top_core_KE_n1500), .B0(n2141), 
        .Y(top_core_KE_n827) );
  OAI221XL U20836 ( .A0(top_core_KE_n1501), .A1(n2192), .B0(n2207), .B1(n7069), 
        .C0(top_core_KE_n1502), .Y(top_core_KE_n1500) );
  OAI221XL U20837 ( .A0(n2152), .A1(n6821), .B0(n2158), .B1(n7163), .C0(
        top_core_KE_n1504), .Y(top_core_KE_n1499) );
  BUFX3 U20838 ( .A(top_core_KE_n828), .Y(n1455) );
  OAI21XL U20839 ( .A0(top_core_KE_n1507), .A1(top_core_KE_n1508), .B0(n2141), 
        .Y(top_core_KE_n828) );
  OAI221XL U20840 ( .A0(top_core_KE_n1509), .A1(n2190), .B0(n2207), .B1(n7068), 
        .C0(top_core_KE_n1510), .Y(top_core_KE_n1508) );
  OAI221XL U20841 ( .A0(n2150), .A1(n6901), .B0(n2159), .B1(n7162), .C0(
        top_core_KE_n1512), .Y(top_core_KE_n1507) );
  BUFX3 U20842 ( .A(top_core_KE_n829), .Y(n1456) );
  OAI21XL U20843 ( .A0(top_core_KE_n1515), .A1(top_core_KE_n1516), .B0(n2141), 
        .Y(top_core_KE_n829) );
  OAI221XL U20844 ( .A0(top_core_KE_n1517), .A1(n2194), .B0(n2207), .B1(n7067), 
        .C0(top_core_KE_n1518), .Y(top_core_KE_n1516) );
  OAI221XL U20845 ( .A0(n2150), .A1(n6946), .B0(n2158), .B1(n7161), .C0(
        top_core_KE_n1520), .Y(top_core_KE_n1515) );
  BUFX3 U20846 ( .A(top_core_KE_n830), .Y(n1457) );
  OAI21XL U20847 ( .A0(top_core_KE_n1523), .A1(top_core_KE_n1524), .B0(n2141), 
        .Y(top_core_KE_n830) );
  OAI221XL U20848 ( .A0(top_core_KE_n1525), .A1(n2193), .B0(n2207), .B1(n7066), 
        .C0(top_core_KE_n1526), .Y(top_core_KE_n1524) );
  OAI221XL U20849 ( .A0(n2150), .A1(n6962), .B0(n2159), .B1(n7160), .C0(
        top_core_KE_n1528), .Y(top_core_KE_n1523) );
  BUFX3 U20850 ( .A(top_core_KE_n831), .Y(n1458) );
  OAI21XL U20851 ( .A0(top_core_KE_n1531), .A1(top_core_KE_n1532), .B0(n2142), 
        .Y(top_core_KE_n831) );
  OAI221XL U20852 ( .A0(top_core_KE_n1533), .A1(n2195), .B0(n2207), .B1(n7065), 
        .C0(top_core_KE_n1534), .Y(top_core_KE_n1532) );
  OAI221XL U20853 ( .A0(n2150), .A1(n6973), .B0(n2159), .B1(n7159), .C0(
        top_core_KE_n1536), .Y(top_core_KE_n1531) );
  BUFX3 U20854 ( .A(top_core_KE_n832), .Y(n1459) );
  OAI21XL U20855 ( .A0(top_core_KE_n1539), .A1(top_core_KE_n1540), .B0(n2142), 
        .Y(top_core_KE_n832) );
  OAI221XL U20856 ( .A0(top_core_KE_n1541), .A1(n2191), .B0(n2207), .B1(n7064), 
        .C0(top_core_KE_n1542), .Y(top_core_KE_n1540) );
  OAI221XL U20857 ( .A0(n2150), .A1(n6983), .B0(n2159), .B1(n7158), .C0(
        top_core_KE_n1544), .Y(top_core_KE_n1539) );
  BUFX3 U20858 ( .A(top_core_KE_n833), .Y(n1460) );
  OAI21XL U20859 ( .A0(top_core_KE_n1547), .A1(top_core_KE_n1548), .B0(n2142), 
        .Y(top_core_KE_n833) );
  OAI221XL U20860 ( .A0(top_core_KE_n1549), .A1(n2192), .B0(n2207), .B1(n7063), 
        .C0(top_core_KE_n1550), .Y(top_core_KE_n1548) );
  OAI221XL U20861 ( .A0(n2150), .A1(n6379), .B0(n2159), .B1(n7157), .C0(
        top_core_KE_n1552), .Y(top_core_KE_n1547) );
  BUFX3 U20862 ( .A(top_core_KE_n834), .Y(n1461) );
  OAI21XL U20863 ( .A0(top_core_KE_n1555), .A1(top_core_KE_n1556), .B0(n2142), 
        .Y(top_core_KE_n834) );
  OAI221XL U20864 ( .A0(top_core_KE_n1557), .A1(n2190), .B0(n2207), .B1(n7062), 
        .C0(top_core_KE_n1558), .Y(top_core_KE_n1556) );
  OAI221XL U20865 ( .A0(n2150), .A1(n6386), .B0(n2159), .B1(n7156), .C0(
        top_core_KE_n1560), .Y(top_core_KE_n1555) );
  BUFX3 U20866 ( .A(top_core_KE_n835), .Y(n1462) );
  OAI21XL U20867 ( .A0(top_core_KE_n1563), .A1(top_core_KE_n1564), .B0(n2142), 
        .Y(top_core_KE_n835) );
  OAI221XL U20868 ( .A0(top_core_KE_n1565), .A1(n2194), .B0(n2207), .B1(n7061), 
        .C0(top_core_KE_n1566), .Y(top_core_KE_n1564) );
  OAI221XL U20869 ( .A0(n2150), .A1(n6783), .B0(n2159), .B1(n7155), .C0(
        top_core_KE_n1568), .Y(top_core_KE_n1563) );
  BUFX3 U20870 ( .A(top_core_KE_n836), .Y(n1463) );
  OAI21XL U20871 ( .A0(top_core_KE_n1571), .A1(top_core_KE_n1572), .B0(n2142), 
        .Y(top_core_KE_n836) );
  OAI221XL U20872 ( .A0(top_core_KE_n1573), .A1(n2193), .B0(n2207), .B1(n7060), 
        .C0(top_core_KE_n1574), .Y(top_core_KE_n1572) );
  OAI221XL U20873 ( .A0(n2150), .A1(n6855), .B0(n2159), .B1(n7154), .C0(
        top_core_KE_n1576), .Y(top_core_KE_n1571) );
  BUFX3 U20874 ( .A(top_core_KE_n837), .Y(n1464) );
  OAI21XL U20875 ( .A0(top_core_KE_n1579), .A1(top_core_KE_n1580), .B0(n2142), 
        .Y(top_core_KE_n837) );
  OAI221XL U20876 ( .A0(top_core_KE_n1581), .A1(n2195), .B0(n2206), .B1(n7059), 
        .C0(top_core_KE_n1582), .Y(top_core_KE_n1580) );
  OAI221XL U20877 ( .A0(n2150), .A1(n6931), .B0(n2159), .B1(n7153), .C0(
        top_core_KE_n1584), .Y(top_core_KE_n1579) );
  BUFX3 U20878 ( .A(top_core_KE_n838), .Y(n1465) );
  OAI21XL U20879 ( .A0(top_core_KE_n1587), .A1(top_core_KE_n1588), .B0(n2142), 
        .Y(top_core_KE_n838) );
  OAI221XL U20880 ( .A0(top_core_KE_n1589), .A1(n2194), .B0(n2206), .B1(n7058), 
        .C0(top_core_KE_n1590), .Y(top_core_KE_n1588) );
  OAI221XL U20881 ( .A0(n2150), .A1(n6956), .B0(n2159), .B1(n7152), .C0(
        top_core_KE_n1592), .Y(top_core_KE_n1587) );
  BUFX3 U20882 ( .A(top_core_KE_n839), .Y(n1466) );
  OAI21XL U20883 ( .A0(top_core_KE_n1595), .A1(top_core_KE_n1596), .B0(n2142), 
        .Y(top_core_KE_n839) );
  OAI221XL U20884 ( .A0(top_core_KE_n1597), .A1(n2194), .B0(n2206), .B1(n7057), 
        .C0(top_core_KE_n1598), .Y(top_core_KE_n1596) );
  OAI221XL U20885 ( .A0(n2150), .A1(n6968), .B0(n2159), .B1(n7151), .C0(
        top_core_KE_n1600), .Y(top_core_KE_n1595) );
  BUFX3 U20886 ( .A(top_core_KE_n840), .Y(n1467) );
  OAI21XL U20887 ( .A0(top_core_KE_n1603), .A1(top_core_KE_n1604), .B0(n2142), 
        .Y(top_core_KE_n840) );
  OAI221XL U20888 ( .A0(top_core_KE_n1605), .A1(n2194), .B0(n2206), .B1(n7056), 
        .C0(top_core_KE_n1606), .Y(top_core_KE_n1604) );
  OAI221XL U20889 ( .A0(n2151), .A1(n6978), .B0(n2160), .B1(n7150), .C0(
        top_core_KE_n1608), .Y(top_core_KE_n1603) );
  BUFX3 U20890 ( .A(top_core_KE_n841), .Y(n1468) );
  OAI21XL U20891 ( .A0(top_core_KE_n1611), .A1(top_core_KE_n1612), .B0(n2142), 
        .Y(top_core_KE_n841) );
  OAI221XL U20892 ( .A0(top_core_KE_n1613), .A1(n2194), .B0(n2206), .B1(n7055), 
        .C0(top_core_KE_n1614), .Y(top_core_KE_n1612) );
  OAI221XL U20893 ( .A0(n2150), .A1(n6989), .B0(n2159), .B1(n7149), .C0(
        top_core_KE_n1616), .Y(top_core_KE_n1611) );
  BUFX3 U20894 ( .A(top_core_KE_n842), .Y(n1469) );
  OAI21XL U20895 ( .A0(top_core_KE_n1619), .A1(top_core_KE_n1620), .B0(n2142), 
        .Y(top_core_KE_n842) );
  OAI221XL U20896 ( .A0(top_core_KE_n1621), .A1(n2194), .B0(n2206), .B1(n7054), 
        .C0(top_core_KE_n1622), .Y(top_core_KE_n1620) );
  OAI221XL U20897 ( .A0(n2151), .A1(n1146), .B0(n2160), .B1(n7148), .C0(
        top_core_KE_n1624), .Y(top_core_KE_n1619) );
  BUFX3 U20898 ( .A(top_core_KE_n843), .Y(n1470) );
  OAI21XL U20899 ( .A0(top_core_KE_n1627), .A1(top_core_KE_n1628), .B0(n2142), 
        .Y(top_core_KE_n843) );
  OAI221XL U20900 ( .A0(top_core_KE_n1629), .A1(n2194), .B0(n2206), .B1(n7053), 
        .C0(top_core_KE_n1630), .Y(top_core_KE_n1628) );
  OAI221XL U20901 ( .A0(n2151), .A1(n1636), .B0(n2160), .B1(n7147), .C0(
        top_core_KE_n1632), .Y(top_core_KE_n1627) );
  BUFX3 U20902 ( .A(top_core_KE_n844), .Y(n1471) );
  OAI21XL U20903 ( .A0(top_core_KE_n1635), .A1(top_core_KE_n1636), .B0(n2143), 
        .Y(top_core_KE_n844) );
  OAI221XL U20904 ( .A0(top_core_KE_n1637), .A1(n2194), .B0(n2206), .B1(n7052), 
        .C0(top_core_KE_n1638), .Y(top_core_KE_n1636) );
  OAI221XL U20905 ( .A0(n2151), .A1(n1159), .B0(n2160), .B1(n7146), .C0(
        top_core_KE_n1640), .Y(top_core_KE_n1635) );
  BUFX3 U20906 ( .A(top_core_KE_n845), .Y(n1472) );
  OAI21XL U20907 ( .A0(top_core_KE_n1643), .A1(top_core_KE_n1644), .B0(n2143), 
        .Y(top_core_KE_n845) );
  OAI221XL U20908 ( .A0(top_core_KE_n1645), .A1(n2194), .B0(n2206), .B1(n7051), 
        .C0(top_core_KE_n1646), .Y(top_core_KE_n1644) );
  OAI221XL U20909 ( .A0(n2151), .A1(n1168), .B0(n2160), .B1(n7145), .C0(
        top_core_KE_n1648), .Y(top_core_KE_n1643) );
  BUFX3 U20910 ( .A(top_core_KE_n846), .Y(n1473) );
  OAI21XL U20911 ( .A0(top_core_KE_n1651), .A1(top_core_KE_n1652), .B0(n2143), 
        .Y(top_core_KE_n846) );
  OAI221XL U20912 ( .A0(top_core_KE_n1653), .A1(n2194), .B0(n2206), .B1(n7050), 
        .C0(top_core_KE_n1654), .Y(top_core_KE_n1652) );
  OAI221XL U20913 ( .A0(n2151), .A1(n1644), .B0(n2160), .B1(n7144), .C0(
        top_core_KE_n1656), .Y(top_core_KE_n1651) );
  BUFX3 U20914 ( .A(top_core_KE_n847), .Y(n1474) );
  OAI21XL U20915 ( .A0(top_core_KE_n1659), .A1(top_core_KE_n1660), .B0(n2143), 
        .Y(top_core_KE_n847) );
  OAI221XL U20916 ( .A0(top_core_KE_n1661), .A1(n2194), .B0(n2206), .B1(n7049), 
        .C0(top_core_KE_n1662), .Y(top_core_KE_n1660) );
  OAI221XL U20917 ( .A0(n2151), .A1(n1656), .B0(n2160), .B1(n7143), .C0(
        top_core_KE_n1664), .Y(top_core_KE_n1659) );
  BUFX3 U20918 ( .A(top_core_KE_n848), .Y(n1475) );
  OAI21XL U20919 ( .A0(top_core_KE_n1667), .A1(top_core_KE_n1668), .B0(n2143), 
        .Y(top_core_KE_n848) );
  OAI221XL U20920 ( .A0(top_core_KE_n1669), .A1(n2194), .B0(n2206), .B1(n7048), 
        .C0(top_core_KE_n1670), .Y(top_core_KE_n1668) );
  OAI221XL U20921 ( .A0(n2151), .A1(n1664), .B0(n2160), .B1(n7142), .C0(
        top_core_KE_n1672), .Y(top_core_KE_n1667) );
  BUFX3 U20922 ( .A(top_core_KE_n849), .Y(n1476) );
  OAI21XL U20923 ( .A0(top_core_KE_n1675), .A1(top_core_KE_n1676), .B0(n2143), 
        .Y(top_core_KE_n849) );
  OAI221XL U20924 ( .A0(top_core_KE_n1677), .A1(n2194), .B0(n2206), .B1(n7047), 
        .C0(top_core_KE_n1678), .Y(top_core_KE_n1676) );
  OAI221XL U20925 ( .A0(n2151), .A1(n6990), .B0(n2160), .B1(n7141), .C0(
        top_core_KE_n1680), .Y(top_core_KE_n1675) );
  BUFX3 U20926 ( .A(top_core_KE_n850), .Y(n1477) );
  OAI21XL U20927 ( .A0(top_core_KE_n1683), .A1(top_core_KE_n1684), .B0(n2143), 
        .Y(top_core_KE_n850) );
  OAI221XL U20928 ( .A0(top_core_KE_n1685), .A1(n2195), .B0(n2206), .B1(n7046), 
        .C0(top_core_KE_n1686), .Y(top_core_KE_n1684) );
  OAI221XL U20929 ( .A0(n2151), .A1(n1185), .B0(n2160), .B1(n7140), .C0(
        top_core_KE_n1688), .Y(top_core_KE_n1683) );
  BUFX3 U20930 ( .A(top_core_KE_n851), .Y(n1478) );
  OAI21XL U20931 ( .A0(top_core_KE_n1691), .A1(top_core_KE_n1692), .B0(n2143), 
        .Y(top_core_KE_n851) );
  OAI221XL U20932 ( .A0(top_core_KE_n1693), .A1(n2195), .B0(n2209), .B1(n7045), 
        .C0(top_core_KE_n1694), .Y(top_core_KE_n1692) );
  OAI221XL U20933 ( .A0(n2151), .A1(n1670), .B0(n2160), .B1(n7139), .C0(
        top_core_KE_n1696), .Y(top_core_KE_n1691) );
  BUFX3 U20934 ( .A(top_core_KE_n852), .Y(n1479) );
  OAI21XL U20935 ( .A0(top_core_KE_n1699), .A1(top_core_KE_n1700), .B0(n2143), 
        .Y(top_core_KE_n852) );
  OAI221XL U20936 ( .A0(top_core_KE_n1701), .A1(n2195), .B0(n2210), .B1(n7044), 
        .C0(top_core_KE_n1702), .Y(top_core_KE_n1700) );
  OAI221XL U20937 ( .A0(n2152), .A1(n1150), .B0(n2159), .B1(n7138), .C0(
        top_core_KE_n1704), .Y(top_core_KE_n1699) );
  BUFX3 U20938 ( .A(top_core_KE_n853), .Y(n1480) );
  OAI21XL U20939 ( .A0(top_core_KE_n1707), .A1(top_core_KE_n1708), .B0(n2143), 
        .Y(top_core_KE_n853) );
  OAI221XL U20940 ( .A0(top_core_KE_n1709), .A1(n2195), .B0(n2208), .B1(n7043), 
        .C0(top_core_KE_n1710), .Y(top_core_KE_n1708) );
  OAI221XL U20941 ( .A0(n2151), .A1(n1166), .B0(n2160), .B1(n7137), .C0(
        top_core_KE_n1712), .Y(top_core_KE_n1707) );
  BUFX3 U20942 ( .A(top_core_KE_n854), .Y(n1481) );
  OAI21XL U20943 ( .A0(top_core_KE_n1715), .A1(top_core_KE_n1716), .B0(n2143), 
        .Y(top_core_KE_n854) );
  OAI221XL U20944 ( .A0(top_core_KE_n1717), .A1(n2195), .B0(n2206), .B1(n7042), 
        .C0(top_core_KE_n1718), .Y(top_core_KE_n1716) );
  OAI221XL U20945 ( .A0(n2152), .A1(n1676), .B0(n2160), .B1(n7136), .C0(
        top_core_KE_n1720), .Y(top_core_KE_n1715) );
  BUFX3 U20946 ( .A(top_core_KE_n855), .Y(n1482) );
  OAI21XL U20947 ( .A0(top_core_KE_n1723), .A1(top_core_KE_n1724), .B0(n2143), 
        .Y(top_core_KE_n855) );
  OAI221XL U20948 ( .A0(top_core_KE_n1725), .A1(n2195), .B0(n2209), .B1(n7041), 
        .C0(top_core_KE_n1726), .Y(top_core_KE_n1724) );
  OAI221XL U20949 ( .A0(n2152), .A1(n1686), .B0(n2155), .B1(n7135), .C0(
        top_core_KE_n1728), .Y(top_core_KE_n1723) );
  BUFX3 U20950 ( .A(top_core_KE_n856), .Y(n1483) );
  OAI21XL U20951 ( .A0(top_core_KE_n1731), .A1(top_core_KE_n1732), .B0(n2143), 
        .Y(top_core_KE_n856) );
  OAI221XL U20952 ( .A0(top_core_KE_n1733), .A1(n2195), .B0(n2210), .B1(n7040), 
        .C0(top_core_KE_n1734), .Y(top_core_KE_n1732) );
  OAI221XL U20953 ( .A0(n2152), .A1(n1692), .B0(n2156), .B1(n7134), .C0(
        top_core_KE_n1736), .Y(top_core_KE_n1731) );
  BUFX3 U20954 ( .A(top_core_KE_n857), .Y(n1484) );
  OAI21XL U20955 ( .A0(top_core_KE_n1739), .A1(top_core_KE_n1740), .B0(n2144), 
        .Y(top_core_KE_n857) );
  OAI221XL U20956 ( .A0(top_core_KE_n1741), .A1(n2195), .B0(n2208), .B1(n7039), 
        .C0(top_core_KE_n1742), .Y(top_core_KE_n1740) );
  OAI221XL U20957 ( .A0(n2152), .A1(n6994), .B0(n2158), .B1(n7133), .C0(
        top_core_KE_n1744), .Y(top_core_KE_n1739) );
  BUFX3 U20958 ( .A(top_core_KE_n858), .Y(n1485) );
  OAI21XL U20959 ( .A0(top_core_KE_n1747), .A1(top_core_KE_n1748), .B0(n2144), 
        .Y(top_core_KE_n858) );
  OAI221XL U20960 ( .A0(top_core_KE_n1749), .A1(n2195), .B0(n2206), .B1(n7038), 
        .C0(top_core_KE_n1750), .Y(top_core_KE_n1748) );
  OAI221XL U20961 ( .A0(n2152), .A1(n1186), .B0(n2159), .B1(n7132), .C0(
        top_core_KE_n1752), .Y(top_core_KE_n1747) );
  BUFX3 U20962 ( .A(top_core_KE_n859), .Y(n1486) );
  OAI21XL U20963 ( .A0(top_core_KE_n1755), .A1(top_core_KE_n1756), .B0(n2144), 
        .Y(top_core_KE_n859) );
  OAI221XL U20964 ( .A0(top_core_KE_n1757), .A1(n2195), .B0(n2209), .B1(n7037), 
        .C0(top_core_KE_n1758), .Y(top_core_KE_n1756) );
  OAI221XL U20965 ( .A0(n2152), .A1(n1699), .B0(n2154), .B1(n7131), .C0(
        top_core_KE_n1760), .Y(top_core_KE_n1755) );
  BUFX3 U20966 ( .A(top_core_KE_n860), .Y(n1487) );
  OAI21XL U20967 ( .A0(top_core_KE_n1763), .A1(top_core_KE_n1764), .B0(n2144), 
        .Y(top_core_KE_n860) );
  OAI221XL U20968 ( .A0(top_core_KE_n1765), .A1(n2195), .B0(n2210), .B1(n7036), 
        .C0(top_core_KE_n1766), .Y(top_core_KE_n1764) );
  OAI221XL U20969 ( .A0(n2152), .A1(n1199), .B0(n2157), .B1(n7130), .C0(
        top_core_KE_n1768), .Y(top_core_KE_n1763) );
  BUFX3 U20970 ( .A(top_core_KE_n861), .Y(n1488) );
  OAI21XL U20971 ( .A0(top_core_KE_n1771), .A1(top_core_KE_n1772), .B0(n2144), 
        .Y(top_core_KE_n861) );
  OAI221XL U20972 ( .A0(top_core_KE_n1773), .A1(n2195), .B0(n2205), .B1(n7035), 
        .C0(top_core_KE_n1774), .Y(top_core_KE_n1772) );
  OAI221XL U20973 ( .A0(n2152), .A1(n1208), .B0(n2153), .B1(n7129), .C0(
        top_core_KE_n1776), .Y(top_core_KE_n1771) );
  BUFX3 U20974 ( .A(top_core_KE_n862), .Y(n1489) );
  OAI21XL U20975 ( .A0(top_core_KE_n1779), .A1(top_core_KE_n1780), .B0(n2144), 
        .Y(top_core_KE_n862) );
  OAI221XL U20976 ( .A0(top_core_KE_n1781), .A1(n2194), .B0(n2205), .B1(n7034), 
        .C0(top_core_KE_n1782), .Y(top_core_KE_n1780) );
  OAI221XL U20977 ( .A0(n2152), .A1(n1706), .B0(n2154), .B1(n7128), .C0(
        top_core_KE_n1784), .Y(top_core_KE_n1779) );
  BUFX3 U20978 ( .A(top_core_KE_n863), .Y(n1490) );
  OAI21XL U20979 ( .A0(top_core_KE_n1787), .A1(top_core_KE_n1788), .B0(n2144), 
        .Y(top_core_KE_n863) );
  OAI221XL U20980 ( .A0(top_core_KE_n1789), .A1(n2192), .B0(n2205), .B1(n7033), 
        .C0(top_core_KE_n1790), .Y(top_core_KE_n1788) );
  OAI221XL U20981 ( .A0(n2152), .A1(n1715), .B0(n2160), .B1(n7127), .C0(
        top_core_KE_n1792), .Y(top_core_KE_n1787) );
  BUFX3 U20982 ( .A(top_core_KE_n864), .Y(n1491) );
  OAI21XL U20983 ( .A0(top_core_KE_n1795), .A1(top_core_KE_n1796), .B0(n2144), 
        .Y(top_core_KE_n864) );
  OAI221XL U20984 ( .A0(top_core_KE_n1797), .A1(n2195), .B0(n2205), .B1(n7032), 
        .C0(top_core_KE_n1798), .Y(top_core_KE_n1796) );
  OAI221XL U20985 ( .A0(n2146), .A1(n1721), .B0(n2160), .B1(n7126), .C0(
        top_core_KE_n1800), .Y(top_core_KE_n1795) );
  BUFX3 U20986 ( .A(top_core_KE_n865), .Y(n1492) );
  OAI21XL U20987 ( .A0(top_core_KE_n1803), .A1(top_core_KE_n1804), .B0(n2144), 
        .Y(top_core_KE_n865) );
  OAI221XL U20988 ( .A0(top_core_KE_n1805), .A1(n2190), .B0(n2205), .B1(n7031), 
        .C0(top_core_KE_n1806), .Y(top_core_KE_n1804) );
  OAI221XL U20989 ( .A0(n2152), .A1(n6995), .B0(n2155), .B1(n7125), .C0(
        top_core_KE_n1808), .Y(top_core_KE_n1803) );
  BUFX3 U20990 ( .A(top_core_KE_n866), .Y(n1493) );
  OAI21XL U20991 ( .A0(top_core_KE_n1811), .A1(top_core_KE_n1812), .B0(n2144), 
        .Y(top_core_KE_n866) );
  OAI221XL U20992 ( .A0(top_core_KE_n1813), .A1(n2191), .B0(n2205), .B1(n7030), 
        .C0(top_core_KE_n1814), .Y(top_core_KE_n1812) );
  OAI221XL U20993 ( .A0(n2150), .A1(n1225), .B0(n2155), .B1(n7124), .C0(
        top_core_KE_n1816), .Y(top_core_KE_n1811) );
  BUFX3 U20994 ( .A(top_core_KE_n867), .Y(n1494) );
  OAI21XL U20995 ( .A0(top_core_KE_n1819), .A1(top_core_KE_n1820), .B0(n2144), 
        .Y(top_core_KE_n867) );
  OAI221XL U20996 ( .A0(top_core_KE_n1821), .A1(n2191), .B0(n2205), .B1(n7029), 
        .C0(top_core_KE_n1822), .Y(top_core_KE_n1820) );
  OAI221XL U20997 ( .A0(n2151), .A1(n1728), .B0(n2156), .B1(n7123), .C0(
        top_core_KE_n1824), .Y(top_core_KE_n1819) );
  BUFX3 U20998 ( .A(top_core_KE_n868), .Y(n1495) );
  OAI21XL U20999 ( .A0(top_core_KE_n1827), .A1(top_core_KE_n1828), .B0(n2144), 
        .Y(top_core_KE_n868) );
  OAI221XL U21000 ( .A0(top_core_KE_n1829), .A1(n2192), .B0(n2205), .B1(n7028), 
        .C0(top_core_KE_n1830), .Y(top_core_KE_n1828) );
  OAI221XL U21001 ( .A0(n2148), .A1(n1190), .B0(n2158), .B1(n7122), .C0(
        top_core_KE_n1832), .Y(top_core_KE_n1827) );
  BUFX3 U21002 ( .A(top_core_KE_n869), .Y(n1496) );
  OAI21XL U21003 ( .A0(top_core_KE_n1835), .A1(top_core_KE_n1836), .B0(n2144), 
        .Y(top_core_KE_n869) );
  OAI221XL U21004 ( .A0(top_core_KE_n1837), .A1(n2194), .B0(n2205), .B1(n7027), 
        .C0(top_core_KE_n1838), .Y(top_core_KE_n1836) );
  OAI221XL U21005 ( .A0(n2149), .A1(n1206), .B0(n2159), .B1(n7121), .C0(
        top_core_KE_n1840), .Y(top_core_KE_n1835) );
  BUFX3 U21006 ( .A(top_core_KE_n870), .Y(n1497) );
  OAI21XL U21007 ( .A0(top_core_KE_n1843), .A1(top_core_KE_n1844), .B0(n2142), 
        .Y(top_core_KE_n870) );
  OAI221XL U21008 ( .A0(top_core_KE_n1845), .A1(n2193), .B0(n2205), .B1(n7026), 
        .C0(top_core_KE_n1846), .Y(top_core_KE_n1844) );
  OAI221XL U21009 ( .A0(n2145), .A1(n1735), .B0(n2157), .B1(n7120), .C0(
        top_core_KE_n1848), .Y(top_core_KE_n1843) );
  BUFX3 U21010 ( .A(top_core_KE_n871), .Y(n1498) );
  OAI21XL U21011 ( .A0(top_core_KE_n1851), .A1(top_core_KE_n1852), .B0(n2143), 
        .Y(top_core_KE_n871) );
  OAI221XL U21012 ( .A0(top_core_KE_n1853), .A1(n2195), .B0(n2205), .B1(n7025), 
        .C0(top_core_KE_n1854), .Y(top_core_KE_n1852) );
  OAI221XL U21013 ( .A0(n2151), .A1(n1744), .B0(n2153), .B1(n7119), .C0(
        top_core_KE_n1856), .Y(top_core_KE_n1851) );
  BUFX3 U21014 ( .A(top_core_KE_n872), .Y(n1499) );
  OAI21XL U21015 ( .A0(top_core_KE_n1859), .A1(top_core_KE_n1860), .B0(n2142), 
        .Y(top_core_KE_n872) );
  OAI221XL U21016 ( .A0(top_core_KE_n1861), .A1(n2190), .B0(n2205), .B1(n7024), 
        .C0(top_core_KE_n1862), .Y(top_core_KE_n1860) );
  OAI221XL U21017 ( .A0(n2145), .A1(n1750), .B0(n2153), .B1(n7118), .C0(
        top_core_KE_n1867), .Y(top_core_KE_n1859) );
  BUFX3 U21018 ( .A(top_core_KE_n753), .Y(n1380) );
  OAI21XL U21019 ( .A0(top_core_KE_n963), .A1(n6392), .B0(n2137), .Y(
        top_core_KE_n753) );
  INVX1 U21020 ( .A(top_core_KE_n964), .Y(n6392) );
  OAI221XL U21021 ( .A0(n2145), .A1(n6332), .B0(n2153), .B1(n7237), .C0(
        top_core_KE_n968), .Y(top_core_KE_n963) );
  BUFX3 U21022 ( .A(top_core_KE_n754), .Y(n1381) );
  OAI21XL U21023 ( .A0(top_core_KE_n970), .A1(n6400), .B0(n2141), .Y(
        top_core_KE_n754) );
  INVX1 U21024 ( .A(top_core_KE_n971), .Y(n6400) );
  OAI221XL U21025 ( .A0(n2145), .A1(n6396), .B0(n2153), .B1(n7236), .C0(
        top_core_KE_n975), .Y(top_core_KE_n970) );
  BUFX3 U21026 ( .A(top_core_KE_n755), .Y(n1382) );
  OAI21XL U21027 ( .A0(top_core_KE_n977), .A1(n6478), .B0(n2144), .Y(
        top_core_KE_n755) );
  INVX1 U21028 ( .A(top_core_KE_n978), .Y(n6478) );
  OAI221XL U21029 ( .A0(n2145), .A1(n6444), .B0(n2153), .B1(n7235), .C0(
        top_core_KE_n982), .Y(top_core_KE_n977) );
  BUFX3 U21030 ( .A(top_core_KE_n756), .Y(n1383) );
  OAI21XL U21031 ( .A0(top_core_KE_n984), .A1(n6488), .B0(n2142), .Y(
        top_core_KE_n756) );
  INVX1 U21032 ( .A(top_core_KE_n985), .Y(n6488) );
  OAI221XL U21033 ( .A0(n2145), .A1(n6535), .B0(n2153), .B1(n7234), .C0(
        top_core_KE_n989), .Y(top_core_KE_n984) );
  BUFX3 U21034 ( .A(top_core_KE_n757), .Y(n1384) );
  OAI21XL U21035 ( .A0(top_core_KE_n991), .A1(n6491), .B0(n2137), .Y(
        top_core_KE_n757) );
  INVX1 U21036 ( .A(top_core_KE_n992), .Y(n6491) );
  OAI221XL U21037 ( .A0(n2146), .A1(n6630), .B0(n2154), .B1(n7233), .C0(
        top_core_KE_n996), .Y(top_core_KE_n991) );
  BUFX3 U21038 ( .A(top_core_KE_n758), .Y(n1385) );
  OAI21XL U21039 ( .A0(top_core_KE_n998), .A1(n6494), .B0(n2143), .Y(
        top_core_KE_n758) );
  INVX1 U21040 ( .A(top_core_KE_n999), .Y(n6494) );
  OAI221XL U21041 ( .A0(n2146), .A1(n6663), .B0(n2154), .B1(n7232), .C0(
        top_core_KE_n1003), .Y(top_core_KE_n998) );
  BUFX3 U21042 ( .A(top_core_KE_n759), .Y(n1386) );
  OAI21XL U21043 ( .A0(top_core_KE_n1005), .A1(n6498), .B0(n2138), .Y(
        top_core_KE_n759) );
  INVX1 U21044 ( .A(top_core_KE_n1006), .Y(n6498) );
  OAI221XL U21045 ( .A0(n2146), .A1(n6678), .B0(n2154), .B1(n7231), .C0(
        top_core_KE_n1010), .Y(top_core_KE_n1005) );
  BUFX3 U21046 ( .A(top_core_KE_n760), .Y(n1387) );
  OAI21XL U21047 ( .A0(top_core_KE_n1012), .A1(n6501), .B0(n2139), .Y(
        top_core_KE_n760) );
  INVX1 U21048 ( .A(top_core_KE_n1013), .Y(n6501) );
  OAI221XL U21049 ( .A0(n2146), .A1(n6685), .B0(n2154), .B1(n7230), .C0(
        top_core_KE_n1017), .Y(top_core_KE_n1012) );
  BUFX3 U21050 ( .A(top_core_KE_n785), .Y(n1412) );
  OAI21XL U21051 ( .A0(top_core_KE_n1187), .A1(n6334), .B0(n2138), .Y(
        top_core_KE_n785) );
  INVX1 U21052 ( .A(top_core_KE_n1188), .Y(n6334) );
  OAI221XL U21053 ( .A0(n2147), .A1(n6991), .B0(n2156), .B1(n7205), .C0(
        top_core_KE_n1192), .Y(top_core_KE_n1187) );
  BUFX3 U21054 ( .A(top_core_KE_n786), .Y(n1413) );
  OAI21XL U21055 ( .A0(top_core_KE_n1194), .A1(n6398), .B0(n2138), .Y(
        top_core_KE_n786) );
  INVX1 U21056 ( .A(top_core_KE_n1195), .Y(n6398) );
  OAI221XL U21057 ( .A0(n2147), .A1(n6404), .B0(n2156), .B1(n7204), .C0(
        top_core_KE_n1199), .Y(top_core_KE_n1194) );
  BUFX3 U21058 ( .A(top_core_KE_n787), .Y(n1414) );
  OAI21XL U21059 ( .A0(top_core_KE_n1201), .A1(n6446), .B0(n2138), .Y(
        top_core_KE_n787) );
  INVX1 U21060 ( .A(top_core_KE_n1202), .Y(n6446) );
  OAI221XL U21061 ( .A0(n2147), .A1(n6482), .B0(n2156), .B1(n7203), .C0(
        top_core_KE_n1206), .Y(top_core_KE_n1201) );
  BUFX3 U21062 ( .A(top_core_KE_n788), .Y(n1415) );
  OAI21XL U21063 ( .A0(top_core_KE_n1208), .A1(n6487), .B0(n2138), .Y(
        top_core_KE_n788) );
  INVX1 U21064 ( .A(top_core_KE_n1209), .Y(n6487) );
  OAI221XL U21065 ( .A0(n2147), .A1(n6562), .B0(n2156), .B1(n7202), .C0(
        top_core_KE_n1213), .Y(top_core_KE_n1208) );
  BUFX3 U21066 ( .A(top_core_KE_n789), .Y(n1416) );
  OAI21XL U21067 ( .A0(top_core_KE_n1215), .A1(n6490), .B0(n2138), .Y(
        top_core_KE_n789) );
  INVX1 U21068 ( .A(top_core_KE_n1216), .Y(n6490) );
  OAI221XL U21069 ( .A0(n2147), .A1(n6641), .B0(n2156), .B1(n7201), .C0(
        top_core_KE_n1220), .Y(top_core_KE_n1215) );
  BUFX3 U21070 ( .A(top_core_KE_n790), .Y(n1417) );
  OAI21XL U21071 ( .A0(top_core_KE_n1222), .A1(n6493), .B0(n2138), .Y(
        top_core_KE_n790) );
  INVX1 U21072 ( .A(top_core_KE_n1223), .Y(n6493) );
  OAI221XL U21073 ( .A0(n2147), .A1(n6669), .B0(n2156), .B1(n7200), .C0(
        top_core_KE_n1227), .Y(top_core_KE_n1222) );
  BUFX3 U21074 ( .A(top_core_KE_n791), .Y(n1418) );
  OAI21XL U21075 ( .A0(top_core_KE_n1229), .A1(n6497), .B0(n2138), .Y(
        top_core_KE_n791) );
  INVX1 U21076 ( .A(top_core_KE_n1230), .Y(n6497) );
  OAI221XL U21077 ( .A0(n2147), .A1(n6684), .B0(n2156), .B1(n7199), .C0(
        top_core_KE_n1234), .Y(top_core_KE_n1229) );
  BUFX3 U21078 ( .A(top_core_KE_n792), .Y(n1419) );
  OAI21XL U21079 ( .A0(top_core_KE_n1236), .A1(n6500), .B0(n2138), .Y(
        top_core_KE_n792) );
  INVX1 U21080 ( .A(top_core_KE_n1237), .Y(n6500) );
  OAI221XL U21081 ( .A0(n2147), .A1(n6691), .B0(n2156), .B1(n7198), .C0(
        top_core_KE_n1241), .Y(top_core_KE_n1236) );
  BUFX3 U21082 ( .A(top_core_KE_n793), .Y(n1420) );
  OAI21XL U21083 ( .A0(top_core_KE_n1243), .A1(n6325), .B0(n2139), .Y(
        top_core_KE_n793) );
  INVX1 U21084 ( .A(top_core_KE_n1244), .Y(n6325) );
  OAI221XL U21085 ( .A0(n2148), .A1(n6331), .B0(n2157), .B1(n7197), .C0(
        top_core_KE_n1248), .Y(top_core_KE_n1243) );
  BUFX3 U21086 ( .A(top_core_KE_n794), .Y(n1421) );
  OAI21XL U21087 ( .A0(top_core_KE_n1250), .A1(n6390), .B0(n2139), .Y(
        top_core_KE_n794) );
  INVX1 U21088 ( .A(top_core_KE_n1251), .Y(n6390) );
  OAI221XL U21089 ( .A0(n2148), .A1(n6720), .B0(n2153), .B1(n7196), .C0(
        top_core_KE_n1255), .Y(top_core_KE_n1250) );
  BUFX3 U21090 ( .A(top_core_KE_n795), .Y(n1422) );
  OAI21XL U21091 ( .A0(top_core_KE_n1257), .A1(n6723), .B0(n2139), .Y(
        top_core_KE_n795) );
  INVX1 U21092 ( .A(top_core_KE_n1258), .Y(n6723) );
  OAI221XL U21093 ( .A0(n2148), .A1(n6822), .B0(n2156), .B1(n7195), .C0(
        top_core_KE_n1262), .Y(top_core_KE_n1257) );
  BUFX3 U21094 ( .A(top_core_KE_n796), .Y(n1423) );
  OAI21XL U21095 ( .A0(top_core_KE_n1264), .A1(n6726), .B0(n2139), .Y(
        top_core_KE_n796) );
  INVX1 U21096 ( .A(top_core_KE_n1265), .Y(n6726) );
  OAI221XL U21097 ( .A0(n2148), .A1(n6902), .B0(n2158), .B1(n7194), .C0(
        top_core_KE_n1269), .Y(top_core_KE_n1264) );
  BUFX3 U21098 ( .A(top_core_KE_n797), .Y(n1424) );
  OAI21XL U21099 ( .A0(top_core_KE_n1271), .A1(n6733), .B0(n2139), .Y(
        top_core_KE_n797) );
  INVX1 U21100 ( .A(top_core_KE_n1272), .Y(n6733) );
  OAI221XL U21101 ( .A0(n2148), .A1(n6947), .B0(n2154), .B1(n7193), .C0(
        top_core_KE_n1276), .Y(top_core_KE_n1271) );
  BUFX3 U21102 ( .A(top_core_KE_n798), .Y(n1425) );
  OAI21XL U21103 ( .A0(top_core_KE_n1278), .A1(n6729), .B0(n2139), .Y(
        top_core_KE_n798) );
  INVX1 U21104 ( .A(top_core_KE_n1279), .Y(n6729) );
  OAI221XL U21105 ( .A0(n2148), .A1(n6963), .B0(n2159), .B1(n7192), .C0(
        top_core_KE_n1283), .Y(top_core_KE_n1278) );
  BUFX3 U21106 ( .A(top_core_KE_n799), .Y(n1426) );
  OAI21XL U21107 ( .A0(top_core_KE_n1285), .A1(n6737), .B0(n2139), .Y(
        top_core_KE_n799) );
  INVX1 U21108 ( .A(top_core_KE_n1286), .Y(n6737) );
  OAI221XL U21109 ( .A0(n2148), .A1(n6974), .B0(n2157), .B1(n7191), .C0(
        top_core_KE_n1290), .Y(top_core_KE_n1285) );
  BUFX3 U21110 ( .A(top_core_KE_n800), .Y(n1427) );
  OAI21XL U21111 ( .A0(top_core_KE_n1292), .A1(n6740), .B0(n2139), .Y(
        top_core_KE_n800) );
  INVX1 U21112 ( .A(top_core_KE_n1293), .Y(n6740) );
  OAI221XL U21113 ( .A0(n2148), .A1(n6984), .B0(n2153), .B1(n7190), .C0(
        top_core_KE_n1297), .Y(top_core_KE_n1292) );
  BUFX3 U21114 ( .A(top_core_KE_n801), .Y(n1428) );
  OAI21XL U21115 ( .A0(top_core_KE_n1299), .A1(n6321), .B0(n2139), .Y(
        top_core_KE_n801) );
  INVX1 U21116 ( .A(top_core_KE_n1300), .Y(n6321) );
  OAI221XL U21117 ( .A0(n2148), .A1(n6996), .B0(n2160), .B1(n7189), .C0(
        top_core_KE_n1304), .Y(top_core_KE_n1299) );
  BUFX3 U21118 ( .A(top_core_KE_n802), .Y(n1429) );
  OAI21XL U21119 ( .A0(top_core_KE_n1306), .A1(n6346), .B0(n2139), .Y(
        top_core_KE_n802) );
  INVX1 U21120 ( .A(top_core_KE_n1307), .Y(n6346) );
  OAI221XL U21121 ( .A0(n2148), .A1(n6387), .B0(n2155), .B1(n7188), .C0(
        top_core_KE_n1311), .Y(top_core_KE_n1306) );
  BUFX3 U21122 ( .A(top_core_KE_n803), .Y(n1430) );
  OAI21XL U21123 ( .A0(top_core_KE_n1313), .A1(n6360), .B0(n2139), .Y(
        top_core_KE_n803) );
  INVX1 U21124 ( .A(top_core_KE_n1314), .Y(n6360) );
  OAI221XL U21125 ( .A0(n2148), .A1(n6784), .B0(n2156), .B1(n7187), .C0(
        top_core_KE_n1318), .Y(top_core_KE_n1313) );
  BUFX3 U21126 ( .A(top_core_KE_n804), .Y(n1431) );
  OAI21XL U21127 ( .A0(top_core_KE_n1320), .A1(n6350), .B0(n2139), .Y(
        top_core_KE_n804) );
  INVX1 U21128 ( .A(top_core_KE_n1321), .Y(n6350) );
  OAI221XL U21129 ( .A0(n2148), .A1(n6856), .B0(n2158), .B1(n7186), .C0(
        top_core_KE_n1325), .Y(top_core_KE_n1320) );
  BUFX3 U21130 ( .A(top_core_KE_n805), .Y(n1432) );
  OAI21XL U21131 ( .A0(top_core_KE_n1327), .A1(n6364), .B0(n2139), .Y(
        top_core_KE_n805) );
  INVX1 U21132 ( .A(top_core_KE_n1328), .Y(n6364) );
  OAI221XL U21133 ( .A0(n2149), .A1(n6932), .B0(n2157), .B1(n7185), .C0(
        top_core_KE_n1332), .Y(top_core_KE_n1327) );
  BUFX3 U21134 ( .A(top_core_KE_n806), .Y(n1433) );
  OAI21XL U21135 ( .A0(top_core_KE_n1334), .A1(n6368), .B0(n2140), .Y(
        top_core_KE_n806) );
  INVX1 U21136 ( .A(top_core_KE_n1335), .Y(n6368) );
  OAI221XL U21137 ( .A0(n2149), .A1(n6957), .B0(n2157), .B1(n7184), .C0(
        top_core_KE_n1339), .Y(top_core_KE_n1334) );
  BUFX3 U21138 ( .A(top_core_KE_n807), .Y(n1434) );
  OAI21XL U21139 ( .A0(top_core_KE_n1341), .A1(n6373), .B0(n2140), .Y(
        top_core_KE_n807) );
  INVX1 U21140 ( .A(top_core_KE_n1342), .Y(n6373) );
  OAI221XL U21141 ( .A0(n2149), .A1(n6969), .B0(n2157), .B1(n7183), .C0(
        top_core_KE_n1346), .Y(top_core_KE_n1341) );
  BUFX3 U21142 ( .A(top_core_KE_n808), .Y(n1435) );
  OAI21XL U21143 ( .A0(top_core_KE_n1348), .A1(n6354), .B0(n2140), .Y(
        top_core_KE_n808) );
  INVX1 U21144 ( .A(top_core_KE_n1349), .Y(n6354) );
  OAI221XL U21145 ( .A0(n2149), .A1(n6979), .B0(n2157), .B1(n7182), .C0(
        top_core_KE_n1353), .Y(top_core_KE_n1348) );
  BUFX3 U21146 ( .A(top_core_KE_n744), .Y(n1371) );
  NAND2BX1 U21147 ( .AN(top_core_KE_n892), .B(n2144), .Y(top_core_KE_n744) );
  AOI211X1 U21148 ( .A0(top_core_KE_n894), .A1(top_core_KE_n895), .B0(
        top_core_KE_n896), .C0(top_core_KE_n897), .Y(top_core_KE_n892) );
  OAI2BB2X1 U21149 ( .B0(n1332), .B1(top_core_KE_n2716), .A0N(
        top_core_KE_n2718), .A1N(n1332), .Y(top_core_KE_n4931) );
  XOR2X1 U21150 ( .A(top_core_KE_new_sboxw_23_), .B(top_core_KE_n1925), .Y(
        top_core_KE_n1189) );
  XOR2X1 U21151 ( .A(top_core_KE_new_sboxw_18_), .B(top_core_KE_n1935), .Y(
        top_core_KE_n1224) );
  XOR2X1 U21152 ( .A(top_core_KE_new_sboxw_21_), .B(top_core_KE_n1929), .Y(
        top_core_KE_n1203) );
  NAND4X1 U21153 ( .A(n11756), .B(n11757), .C(n11758), .D(n11759), .Y(n11755)
         );
  AOI21X1 U21154 ( .A0(n6826), .A1(n11765), .B0(n6824), .Y(n11758) );
  OAI22X1 U21155 ( .A0(n11762), .A1(n1795), .B0(n1800), .B1(n11763), .Y(n11760) );
  NAND4X1 U21156 ( .A(top_core_KE_sb1_n184), .B(top_core_KE_sb1_n185), .C(
        top_core_KE_sb1_n186), .D(top_core_KE_sb1_n187), .Y(
        top_core_KE_sb1_n183) );
  AOI21X1 U21157 ( .A0(n6804), .A1(top_core_KE_sb1_n193), .B0(n6802), .Y(
        top_core_KE_sb1_n186) );
  OAI22X1 U21158 ( .A0(top_core_KE_sb1_n190), .A1(n1816), .B0(n1821), .B1(
        top_core_KE_sb1_n191), .Y(top_core_KE_sb1_n188) );
  NAND4X1 U21159 ( .A(n12072), .B(n12073), .C(n12074), .D(n12075), .Y(n12071)
         );
  AOI21X1 U21160 ( .A0(n6507), .A1(n12081), .B0(n6505), .Y(n12074) );
  OAI22X1 U21161 ( .A0(n12078), .A1(n1774), .B0(n1779), .B1(n12079), .Y(n12076) );
  XNOR2X1 U21162 ( .A(top_core_KE_new_sboxw_18_), .B(n6667), .Y(
        top_core_KE_n1000) );
  XNOR2X1 U21163 ( .A(top_core_KE_new_sboxw_21_), .B(n6480), .Y(
        top_core_KE_n979) );
  XNOR2X1 U21164 ( .A(top_core_KE_new_sboxw_23_), .B(n6394), .Y(
        top_core_KE_n965) );
  XOR2X1 U21165 ( .A(top_core_KE_new_sboxw_6_), .B(top_core_KE_n1959), .Y(
        top_core_KE_n1308) );
  XOR2X1 U21166 ( .A(top_core_KE_new_sboxw_8_), .B(top_core_KE_n1955), .Y(
        top_core_KE_n1294) );
  XOR2X1 U21167 ( .A(top_core_KE_new_sboxw_0_), .B(top_core_KE_n1971), .Y(
        top_core_KE_n1350) );
  XOR2X1 U21168 ( .A(top_core_KE_new_sboxw_14_), .B(top_core_KE_n1943), .Y(
        top_core_KE_n1252) );
  XOR2X1 U21169 ( .A(top_core_KE_new_sboxw_9_), .B(top_core_KE_n1953), .Y(
        top_core_KE_n1287) );
  XOR2X1 U21170 ( .A(top_core_KE_new_sboxw_1_), .B(top_core_KE_n1969), .Y(
        top_core_KE_n1343) );
  XOR2X1 U21171 ( .A(top_core_KE_new_sboxw_11_), .B(top_core_KE_n1949), .Y(
        top_core_KE_n1273) );
  XOR2X1 U21172 ( .A(top_core_KE_new_sboxw_3_), .B(top_core_KE_n1965), .Y(
        top_core_KE_n1329) );
  XOR2X1 U21173 ( .A(top_core_KE_new_sboxw_12_), .B(top_core_KE_n1947), .Y(
        top_core_KE_n1266) );
  XOR2X1 U21174 ( .A(top_core_KE_new_sboxw_4_), .B(top_core_KE_n1963), .Y(
        top_core_KE_n1322) );
  AND2X2 U21175 ( .A(n1333), .B(n1334), .Y(top_core_KE_r343_quotient_2_) );
  XOR2X1 U21176 ( .A(top_core_KE_new_sboxw_22_), .B(top_core_KE_n1927), .Y(
        top_core_KE_n1196) );
  XOR2X1 U21177 ( .A(top_core_KE_new_sboxw_16_), .B(top_core_KE_n1939), .Y(
        top_core_KE_n1238) );
  XOR2X1 U21178 ( .A(top_core_KE_new_sboxw_17_), .B(top_core_KE_n1937), .Y(
        top_core_KE_n1231) );
  XOR2X1 U21179 ( .A(top_core_KE_new_sboxw_19_), .B(top_core_KE_n1933), .Y(
        top_core_KE_n1217) );
  XOR2X1 U21180 ( .A(top_core_KE_new_sboxw_20_), .B(top_core_KE_n1931), .Y(
        top_core_KE_n1210) );
  XNOR2X1 U21181 ( .A(top_core_KE_new_sboxw_16_), .B(n6689), .Y(
        top_core_KE_n1014) );
  XNOR2X1 U21182 ( .A(top_core_KE_new_sboxw_22_), .B(n6402), .Y(
        top_core_KE_n972) );
  XNOR2X1 U21183 ( .A(top_core_KE_new_sboxw_17_), .B(n6682), .Y(
        top_core_KE_n1007) );
  XNOR2X1 U21184 ( .A(top_core_KE_new_sboxw_19_), .B(n6639), .Y(
        top_core_KE_n993) );
  XNOR2X1 U21185 ( .A(top_core_KE_new_sboxw_20_), .B(n6560), .Y(
        top_core_KE_n986) );
  AOI21X1 U21186 ( .A0(n4262), .A1(n4261), .B0(top_core_io_n653), .Y(
        top_core_io_N127) );
  XNOR2X1 U21187 ( .A(n6992), .B(top_core_KE_n1425), .Y(top_core_KE_n1681) );
  XNOR2X1 U21188 ( .A(n6993), .B(top_core_KE_n1489), .Y(top_core_KE_n1745) );
  XNOR2X1 U21189 ( .A(n6997), .B(top_core_KE_n1553), .Y(top_core_KE_n1809) );
  XNOR2X1 U21190 ( .A(n1774), .B(top_core_KE_n1441), .Y(top_core_KE_n1697) );
  XNOR2X1 U21191 ( .A(n1795), .B(top_core_KE_n1505), .Y(top_core_KE_n1761) );
  XNOR2X1 U21192 ( .A(n1816), .B(top_core_KE_n1569), .Y(top_core_KE_n1825) );
  XNOR2X1 U21193 ( .A(n1167), .B(top_core_KE_n1457), .Y(top_core_KE_n1713) );
  XNOR2X1 U21194 ( .A(n1209), .B(top_core_KE_n1521), .Y(top_core_KE_n1777) );
  XNOR2X1 U21195 ( .A(n1207), .B(top_core_KE_n1585), .Y(top_core_KE_n1841) );
  XNOR2X1 U21196 ( .A(top_core_KE_n2512), .B(top_core_KE_n2344), .Y(
        top_core_KE_n1361) );
  XNOR2X1 U21197 ( .A(n6338), .B(top_core_KE_n2183), .Y(top_core_KE_n2512) );
  XNOR2X1 U21198 ( .A(n1184), .B(top_core_KE_n1433), .Y(top_core_KE_n1689) );
  XNOR2X1 U21199 ( .A(n1155), .B(top_core_KE_n1449), .Y(top_core_KE_n1705) );
  XNOR2X1 U21200 ( .A(n1170), .B(top_core_KE_n1465), .Y(top_core_KE_n1721) );
  XNOR2X1 U21201 ( .A(n1187), .B(top_core_KE_n1497), .Y(top_core_KE_n1753) );
  XNOR2X1 U21202 ( .A(n1204), .B(top_core_KE_n1513), .Y(top_core_KE_n1769) );
  XNOR2X1 U21203 ( .A(n1211), .B(top_core_KE_n1529), .Y(top_core_KE_n1785) );
  XNOR2X1 U21204 ( .A(n1224), .B(top_core_KE_n1561), .Y(top_core_KE_n1817) );
  XNOR2X1 U21205 ( .A(n1195), .B(top_core_KE_n1577), .Y(top_core_KE_n1833) );
  XNOR2X1 U21206 ( .A(n1210), .B(top_core_KE_n1593), .Y(top_core_KE_n1849) );
  XNOR2X1 U21207 ( .A(n1784), .B(top_core_KE_n1473), .Y(top_core_KE_n1729) );
  XNOR2X1 U21208 ( .A(n1791), .B(top_core_KE_n1481), .Y(top_core_KE_n1737) );
  XNOR2X1 U21209 ( .A(n1805), .B(top_core_KE_n1537), .Y(top_core_KE_n1793) );
  XNOR2X1 U21210 ( .A(n1812), .B(top_core_KE_n1545), .Y(top_core_KE_n1801) );
  XNOR2X1 U21211 ( .A(n1826), .B(top_core_KE_n1601), .Y(top_core_KE_n1857) );
  XNOR2X1 U21212 ( .A(n1833), .B(top_core_KE_n1609), .Y(top_core_KE_n1868) );
  OAI21XL U21213 ( .A0(n1350), .A1(n11684), .B0(n11685), .Y(n11683) );
  OAI21XL U21214 ( .A0(n1352), .A1(top_core_KE_sb1_n109), .B0(
        top_core_KE_sb1_n110), .Y(top_core_KE_sb1_n108) );
  OAI21XL U21215 ( .A0(n1364), .A1(n12315), .B0(n12316), .Y(n12314) );
  OAI21XL U21216 ( .A0(n1367), .A1(n13261), .B0(n13262), .Y(n13260) );
  OAI21XL U21217 ( .A0(n1366), .A1(n12000), .B0(n12001), .Y(n11999) );
  OAI21XL U21218 ( .A0(n1351), .A1(n12946), .B0(n12947), .Y(n12945) );
  OAI21XL U21219 ( .A0(n1365), .A1(n13576), .B0(n13577), .Y(n13575) );
  OAI21XL U21220 ( .A0(n1353), .A1(n12631), .B0(n12632), .Y(n12630) );
  AOI21X1 U21221 ( .A0(n1350), .A1(n6826), .B0(n11656), .Y(n11655) );
  AOI21X1 U21222 ( .A0(n1352), .A1(n6804), .B0(top_core_KE_sb1_n81), .Y(
        top_core_KE_sb1_n80) );
  AOI21X1 U21223 ( .A0(n1364), .A1(n6530), .B0(n12288), .Y(n12287) );
  AOI21X1 U21224 ( .A0(n1367), .A1(n6472), .B0(n13233), .Y(n13232) );
  AOI21X1 U21225 ( .A0(n1366), .A1(n6507), .B0(n11972), .Y(n11971) );
  AOI21X1 U21226 ( .A0(n1351), .A1(n6815), .B0(n12918), .Y(n12917) );
  AOI21X1 U21227 ( .A0(n1365), .A1(n6519), .B0(n13548), .Y(n13547) );
  AOI21X1 U21228 ( .A0(n1353), .A1(n6775), .B0(n12603), .Y(n12602) );
  AND2X2 U21229 ( .A(top_core_KE_n2700), .B(top_core_KE_n2506), .Y(
        top_core_KE_n2699) );
  BUFX3 U21230 ( .A(top_core_EC_ss_in[83]), .Y(n1505) );
  OAI22X1 U21231 ( .A0(n2385), .A1(n6221), .B0(n2422), .B1(n855), .Y(
        top_core_EC_ss_in[83]) );
  BUFX3 U21232 ( .A(top_core_EC_ss_in[3]), .Y(n1517) );
  OAI22X1 U21233 ( .A0(n2389), .A1(n6301), .B0(n2406), .B1(n856), .Y(
        top_core_EC_ss_in[3]) );
  BUFX3 U21234 ( .A(top_core_EC_ss_in[115]), .Y(n1529) );
  OAI22X1 U21235 ( .A0(n2392), .A1(n6189), .B0(n2474), .B1(n860), .Y(
        top_core_EC_ss_in[115]) );
  BUFX3 U21236 ( .A(top_core_EC_ss_in[35]), .Y(n1519) );
  OAI22X1 U21237 ( .A0(n2389), .A1(n6269), .B0(n2404), .B1(n861), .Y(
        top_core_EC_ss_in[35]) );
  BUFX3 U21238 ( .A(top_core_EC_ss_in[43]), .Y(n1516) );
  OAI22X1 U21239 ( .A0(n2384), .A1(n6261), .B0(n2407), .B1(n868), .Y(
        top_core_EC_ss_in[43]) );
  BUFX3 U21240 ( .A(top_core_EC_ss_in[75]), .Y(n1508) );
  OAI22X1 U21241 ( .A0(n2386), .A1(n6229), .B0(n2419), .B1(n869), .Y(
        top_core_EC_ss_in[75]) );
  BUFX3 U21242 ( .A(top_core_EC_ss_in[123]), .Y(n1526) );
  OAI22X1 U21243 ( .A0(n2391), .A1(n6181), .B0(n2440), .B1(n870), .Y(
        top_core_EC_ss_in[123]) );
  BUFX3 U21244 ( .A(top_core_EC_ss_in[27]), .Y(n1521) );
  OAI22X1 U21245 ( .A0(n2390), .A1(n6277), .B0(n2401), .B1(n871), .Y(
        top_core_EC_ss_in[27]) );
  BUFX3 U21246 ( .A(top_core_EC_ss_in[67]), .Y(n1510) );
  OAI22X1 U21247 ( .A0(n2386), .A1(n6237), .B0(n2416), .B1(n872), .Y(
        top_core_EC_ss_in[67]) );
  BUFX3 U21248 ( .A(top_core_EC_ss_in[107]), .Y(n1531) );
  OAI22X1 U21249 ( .A0(n2392), .A1(n6197), .B0(n2398), .B1(n873), .Y(
        top_core_EC_ss_in[107]) );
  BUFX3 U21250 ( .A(top_core_EC_ss_in[19]), .Y(n1523) );
  OAI22X1 U21251 ( .A0(n2390), .A1(n6285), .B0(n2432), .B1(n874), .Y(
        top_core_EC_ss_in[19]) );
  BUFX3 U21252 ( .A(top_core_EC_ss_in[59]), .Y(n1512) );
  OAI22X1 U21253 ( .A0(n2387), .A1(n6245), .B0(n2413), .B1(n875), .Y(
        top_core_EC_ss_in[59]) );
  BUFX3 U21254 ( .A(top_core_EC_ss_in[99]), .Y(n1501) );
  OAI22X1 U21255 ( .A0(n2384), .A1(n6205), .B0(n2406), .B1(n876), .Y(
        top_core_EC_ss_in[99]) );
  BUFX3 U21256 ( .A(top_core_EC_ss_in[11]), .Y(n1527) );
  OAI22X1 U21257 ( .A0(n2391), .A1(n6293), .B0(n2487), .B1(n877), .Y(
        top_core_EC_ss_in[11]) );
  BUFX3 U21258 ( .A(top_core_EC_ss_in[51]), .Y(n1514) );
  OAI22X1 U21259 ( .A0(n2388), .A1(n6253), .B0(n2410), .B1(n878), .Y(
        top_core_EC_ss_in[51]) );
  BUFX3 U21260 ( .A(top_core_EC_ss_in[91]), .Y(n1503) );
  OAI22X1 U21261 ( .A0(n2384), .A1(n6213), .B0(n2425), .B1(n879), .Y(
        top_core_EC_ss_in[91]) );
  INVX1 U21262 ( .A(n1334), .Y(n7007) );
  NAND4BXL U21263 ( .AN(n11703), .B(n11734), .C(n11870), .D(n11871), .Y(n11857) );
  AOI22X1 U21264 ( .A0(n11797), .A1(n577), .B0(n6951), .B1(n1344), .Y(n11870)
         );
  NAND4BXL U21265 ( .AN(top_core_KE_sb1_n128), .B(top_core_KE_sb1_n161), .C(
        top_core_KE_sb1_n299), .D(top_core_KE_sb1_n300), .Y(
        top_core_KE_sb1_n286) );
  AOI22X1 U21266 ( .A0(top_core_KE_sb1_n225), .A1(n578), .B0(n6936), .B1(n1345), .Y(top_core_KE_sb1_n299) );
  NAND4BXL U21267 ( .AN(n12334), .B(n12365), .C(n12501), .D(n12502), .Y(n12488) );
  AOI22X1 U21268 ( .A0(n12428), .A1(n579), .B0(n6661), .B1(n1358), .Y(n12501)
         );
  NAND4BXL U21269 ( .AN(n12019), .B(n12050), .C(n12186), .D(n12187), .Y(n12173) );
  AOI22X1 U21270 ( .A0(n12113), .A1(n581), .B0(n6645), .B1(n1359), .Y(n12186)
         );
  OAI22X1 U21271 ( .A0(n3584), .A1(n6246), .B0(top_core_EC_ss_n176), .B1(n3592), .Y(top_core_EC_add_in_r[58]) );
  OAI22X1 U21272 ( .A0(n3584), .A1(n6245), .B0(top_core_EC_ss_n175), .B1(n3591), .Y(top_core_EC_add_in_r[59]) );
  OAI22X1 U21273 ( .A0(n3585), .A1(n6244), .B0(top_core_EC_ss_n173), .B1(n3600), .Y(top_core_EC_add_in_r[60]) );
  OAI22X1 U21274 ( .A0(n3582), .A1(n6243), .B0(top_core_EC_ss_n172), .B1(n3611), .Y(top_core_EC_add_in_r[61]) );
  OAI22X1 U21275 ( .A0(n3583), .A1(n6242), .B0(top_core_EC_ss_n171), .B1(n3602), .Y(top_core_EC_add_in_r[62]) );
  OAI22X1 U21276 ( .A0(n3585), .A1(n6241), .B0(top_core_EC_ss_n170), .B1(n3601), .Y(top_core_EC_add_in_r[63]) );
  OAI22X1 U21277 ( .A0(n3586), .A1(n6240), .B0(top_core_EC_ss_n169), .B1(n3595), .Y(top_core_EC_add_in_r[64]) );
  OAI22X1 U21278 ( .A0(n3584), .A1(n6239), .B0(top_core_EC_ss_n168), .B1(n3613), .Y(top_core_EC_add_in_r[65]) );
  OAI22X1 U21279 ( .A0(n3582), .A1(n6238), .B0(top_core_EC_ss_n167), .B1(n3627), .Y(top_core_EC_add_in_r[66]) );
  OAI22X1 U21280 ( .A0(n3583), .A1(n6237), .B0(top_core_EC_ss_n166), .B1(n3591), .Y(top_core_EC_add_in_r[67]) );
  OAI22X1 U21281 ( .A0(n3587), .A1(n6236), .B0(top_core_EC_ss_n165), .B1(n3594), .Y(top_core_EC_add_in_r[68]) );
  OAI22X1 U21282 ( .A0(n3585), .A1(n6235), .B0(top_core_EC_ss_n164), .B1(n3589), .Y(top_core_EC_add_in_r[69]) );
  OAI22X1 U21283 ( .A0(n3587), .A1(n6234), .B0(top_core_EC_ss_n162), .B1(n3603), .Y(top_core_EC_add_in_r[70]) );
  OAI22X1 U21284 ( .A0(n3585), .A1(n6233), .B0(top_core_EC_ss_n161), .B1(n3613), .Y(top_core_EC_add_in_r[71]) );
  OAI22X1 U21285 ( .A0(n3585), .A1(n6232), .B0(top_core_EC_ss_n160), .B1(n3612), .Y(top_core_EC_add_in_r[72]) );
  OAI22X1 U21286 ( .A0(n3585), .A1(n6231), .B0(top_core_EC_ss_n159), .B1(n3607), .Y(top_core_EC_add_in_r[73]) );
  OAI22X1 U21287 ( .A0(n3585), .A1(n6230), .B0(top_core_EC_ss_n158), .B1(n3597), .Y(top_core_EC_add_in_r[74]) );
  OAI22X1 U21288 ( .A0(n3585), .A1(n6229), .B0(top_core_EC_ss_n157), .B1(n3589), .Y(top_core_EC_add_in_r[75]) );
  OAI22X1 U21289 ( .A0(n3585), .A1(n6228), .B0(top_core_EC_ss_n156), .B1(n3590), .Y(top_core_EC_add_in_r[76]) );
  OAI22X1 U21290 ( .A0(n3585), .A1(n6227), .B0(top_core_EC_ss_n155), .B1(n3590), .Y(top_core_EC_add_in_r[77]) );
  OAI22X1 U21291 ( .A0(n3585), .A1(n6226), .B0(top_core_EC_ss_n154), .B1(n3590), .Y(top_core_EC_add_in_r[78]) );
  OAI22X1 U21292 ( .A0(n3585), .A1(n6225), .B0(top_core_EC_ss_n153), .B1(n3589), .Y(top_core_EC_add_in_r[79]) );
  OAI22X1 U21293 ( .A0(n3585), .A1(n6224), .B0(top_core_EC_ss_n151), .B1(n3588), .Y(top_core_EC_add_in_r[80]) );
  OAI22X1 U21294 ( .A0(n3585), .A1(n6223), .B0(top_core_EC_ss_n150), .B1(n3588), .Y(top_core_EC_add_in_r[81]) );
  OAI22X1 U21295 ( .A0(n3586), .A1(n6222), .B0(top_core_EC_ss_n149), .B1(n3594), .Y(top_core_EC_add_in_r[82]) );
  OAI22X1 U21296 ( .A0(n3586), .A1(n6221), .B0(top_core_EC_ss_n148), .B1(n3595), .Y(top_core_EC_add_in_r[83]) );
  OAI22X1 U21297 ( .A0(n3586), .A1(n6220), .B0(top_core_EC_ss_n147), .B1(n3597), .Y(top_core_EC_add_in_r[84]) );
  OAI22X1 U21298 ( .A0(n3586), .A1(n6219), .B0(top_core_EC_ss_n146), .B1(n3598), .Y(top_core_EC_add_in_r[85]) );
  OAI22X1 U21299 ( .A0(n3586), .A1(n6218), .B0(top_core_EC_ss_n145), .B1(n3610), .Y(top_core_EC_add_in_r[86]) );
  OAI22X1 U21300 ( .A0(n3586), .A1(n6217), .B0(top_core_EC_ss_n144), .B1(n3609), .Y(top_core_EC_add_in_r[87]) );
  OAI22X1 U21301 ( .A0(n3586), .A1(n6216), .B0(top_core_EC_ss_n143), .B1(n3589), .Y(top_core_EC_add_in_r[88]) );
  OAI22X1 U21302 ( .A0(n3586), .A1(n6215), .B0(top_core_EC_ss_n142), .B1(n3590), .Y(top_core_EC_add_in_r[89]) );
  OAI22X1 U21303 ( .A0(n3586), .A1(n6214), .B0(top_core_EC_ss_n140), .B1(n3606), .Y(top_core_EC_add_in_r[90]) );
  OAI22X1 U21304 ( .A0(n3586), .A1(n6213), .B0(top_core_EC_ss_n139), .B1(n3605), .Y(top_core_EC_add_in_r[91]) );
  OAI22X1 U21305 ( .A0(n3586), .A1(n6212), .B0(top_core_EC_ss_n138), .B1(n3590), .Y(top_core_EC_add_in_r[92]) );
  OAI22X1 U21306 ( .A0(n3587), .A1(n6211), .B0(top_core_EC_ss_n137), .B1(n3596), .Y(top_core_EC_add_in_r[93]) );
  OAI22X1 U21307 ( .A0(n3587), .A1(n6210), .B0(top_core_EC_ss_n136), .B1(n3605), .Y(top_core_EC_add_in_r[94]) );
  OAI22X1 U21308 ( .A0(n3587), .A1(n6209), .B0(top_core_EC_ss_n135), .B1(n3624), .Y(top_core_EC_add_in_r[95]) );
  OAI22X1 U21309 ( .A0(n3587), .A1(n6208), .B0(top_core_EC_ss_n134), .B1(n3602), .Y(top_core_EC_add_in_r[96]) );
  OAI22X1 U21310 ( .A0(n3587), .A1(n6207), .B0(top_core_EC_ss_n133), .B1(n3604), .Y(top_core_EC_add_in_r[97]) );
  OAI22X1 U21311 ( .A0(n3587), .A1(n6206), .B0(top_core_EC_ss_n132), .B1(n3612), .Y(top_core_EC_add_in_r[98]) );
  OAI22X1 U21312 ( .A0(n3587), .A1(n6205), .B0(top_core_EC_ss_n131), .B1(n3605), .Y(top_core_EC_add_in_r[99]) );
  OAI22X1 U21313 ( .A0(n237), .A1(n6204), .B0(top_core_EC_ss_n256), .B1(n3613), 
        .Y(top_core_EC_add_in_r[100]) );
  OAI22X1 U21314 ( .A0(n3586), .A1(n6203), .B0(top_core_EC_ss_n255), .B1(n3603), .Y(top_core_EC_add_in_r[101]) );
  OAI22X1 U21315 ( .A0(n3584), .A1(n6202), .B0(top_core_EC_ss_n254), .B1(n3604), .Y(top_core_EC_add_in_r[102]) );
  OAI22X1 U21316 ( .A0(n3623), .A1(n6201), .B0(top_core_EC_ss_n253), .B1(n3607), .Y(top_core_EC_add_in_r[103]) );
  OAI22X1 U21317 ( .A0(n3586), .A1(n6200), .B0(top_core_EC_ss_n252), .B1(n3598), .Y(top_core_EC_add_in_r[104]) );
  OAI22X1 U21318 ( .A0(n3615), .A1(n6199), .B0(top_core_EC_ss_n251), .B1(n3613), .Y(top_core_EC_add_in_r[105]) );
  OAI22X1 U21319 ( .A0(n3626), .A1(n6198), .B0(top_core_EC_ss_n250), .B1(n3613), .Y(top_core_EC_add_in_r[106]) );
  OAI22X1 U21320 ( .A0(n3615), .A1(n6197), .B0(top_core_EC_ss_n249), .B1(n3612), .Y(top_core_EC_add_in_r[107]) );
  OAI22X1 U21321 ( .A0(n3617), .A1(n6196), .B0(top_core_EC_ss_n248), .B1(n3612), .Y(top_core_EC_add_in_r[108]) );
  OAI22X1 U21322 ( .A0(n3616), .A1(n6195), .B0(top_core_EC_ss_n247), .B1(n3611), .Y(top_core_EC_add_in_r[109]) );
  OAI22X1 U21323 ( .A0(n3615), .A1(n6194), .B0(top_core_EC_ss_n245), .B1(n3601), .Y(top_core_EC_add_in_r[110]) );
  OAI22X1 U21324 ( .A0(n3626), .A1(n6193), .B0(top_core_EC_ss_n244), .B1(n3610), .Y(top_core_EC_add_in_r[111]) );
  OAI22X1 U21325 ( .A0(n3615), .A1(n6192), .B0(top_core_EC_ss_n243), .B1(n3625), .Y(top_core_EC_add_in_r[112]) );
  OAI22X1 U21326 ( .A0(n3617), .A1(n6191), .B0(top_core_EC_ss_n242), .B1(n3606), .Y(top_core_EC_add_in_r[113]) );
  OAI22X1 U21327 ( .A0(n3616), .A1(n6190), .B0(top_core_EC_ss_n241), .B1(n3594), .Y(top_core_EC_add_in_r[114]) );
  OAI22X1 U21328 ( .A0(n3619), .A1(n6189), .B0(top_core_EC_ss_n240), .B1(n3593), .Y(top_core_EC_add_in_r[115]) );
  OAI22X1 U21329 ( .A0(n3618), .A1(n6188), .B0(top_core_EC_ss_n239), .B1(n3603), .Y(top_core_EC_add_in_r[116]) );
  OAI22X1 U21330 ( .A0(n3614), .A1(n6187), .B0(top_core_EC_ss_n238), .B1(n3604), .Y(top_core_EC_add_in_r[117]) );
  OAI22X1 U21331 ( .A0(n3620), .A1(n6186), .B0(top_core_EC_ss_n237), .B1(n3588), .Y(top_core_EC_add_in_r[118]) );
  OAI22X1 U21332 ( .A0(n3621), .A1(n6185), .B0(top_core_EC_ss_n236), .B1(n3607), .Y(top_core_EC_add_in_r[119]) );
  OAI22X1 U21333 ( .A0(n3587), .A1(n6184), .B0(top_core_EC_ss_n234), .B1(n3596), .Y(top_core_EC_add_in_r[120]) );
  OAI22X1 U21334 ( .A0(n3585), .A1(n6183), .B0(top_core_EC_ss_n233), .B1(n3610), .Y(top_core_EC_add_in_r[121]) );
  OAI22X1 U21335 ( .A0(n3586), .A1(n6182), .B0(top_core_EC_ss_n232), .B1(n3610), .Y(top_core_EC_add_in_r[122]) );
  OAI22X1 U21336 ( .A0(n3582), .A1(n6181), .B0(top_core_EC_ss_n231), .B1(n3609), .Y(top_core_EC_add_in_r[123]) );
  OAI22X1 U21337 ( .A0(n3583), .A1(n6180), .B0(top_core_EC_ss_n230), .B1(n3609), .Y(top_core_EC_add_in_r[124]) );
  OAI22X1 U21338 ( .A0(n3587), .A1(n6179), .B0(top_core_EC_ss_n229), .B1(n3608), .Y(top_core_EC_add_in_r[125]) );
  OAI22X1 U21339 ( .A0(n3584), .A1(n6178), .B0(top_core_EC_ss_n228), .B1(n3608), .Y(top_core_EC_add_in_r[126]) );
  OAI22X1 U21340 ( .A0(n3583), .A1(n6177), .B0(top_core_EC_ss_n227), .B1(n3611), .Y(top_core_EC_add_in_r[127]) );
  NOR2X1 U21341 ( .A(n4761), .B(n1582), .Y(top_core_io_N141) );
  NOR2X1 U21342 ( .A(n4760), .B(n1582), .Y(top_core_io_N140) );
  NOR2X1 U21343 ( .A(n4759), .B(n1582), .Y(top_core_io_N139) );
  NOR2X1 U21344 ( .A(n4774), .B(n1582), .Y(top_core_io_N138) );
  NOR2X1 U21345 ( .A(n4773), .B(n1582), .Y(top_core_io_N137) );
  NOR2X1 U21346 ( .A(n4772), .B(n1582), .Y(top_core_io_N136) );
  NOR2X1 U21347 ( .A(n4771), .B(n1582), .Y(top_core_io_N135) );
  NOR2X1 U21348 ( .A(n4770), .B(n1582), .Y(top_core_io_N134) );
  NOR2X1 U21349 ( .A(n4769), .B(n1582), .Y(top_core_io_N133) );
  NOR2X1 U21350 ( .A(n4768), .B(n1582), .Y(top_core_io_N132) );
  NOR2X1 U21351 ( .A(n4767), .B(n1582), .Y(top_core_io_N131) );
  NOR2X1 U21352 ( .A(n4277), .B(n1603), .Y(top_core_io_N505) );
  NOR2X1 U21353 ( .A(n4276), .B(n1603), .Y(top_core_io_N504) );
  NOR2X1 U21354 ( .A(n4275), .B(n1603), .Y(top_core_io_N503) );
  NOR2X1 U21355 ( .A(n4274), .B(n1603), .Y(top_core_io_N502) );
  NOR2X1 U21356 ( .A(n4273), .B(n1603), .Y(top_core_io_N501) );
  NOR2X1 U21357 ( .A(n4272), .B(n1603), .Y(top_core_io_N500) );
  NOR2X1 U21358 ( .A(n4271), .B(n1603), .Y(top_core_io_N499) );
  NOR2X1 U21359 ( .A(n4286), .B(n1603), .Y(top_core_io_N498) );
  NOR2X1 U21360 ( .A(n4285), .B(n1603), .Y(top_core_io_N497) );
  NOR2X1 U21361 ( .A(n4284), .B(n1603), .Y(top_core_io_N496) );
  NOR2X1 U21362 ( .A(n4283), .B(n1603), .Y(top_core_io_N495) );
  NOR2X1 U21363 ( .A(n4282), .B(n1603), .Y(top_core_io_N494) );
  NOR2X1 U21364 ( .A(n4281), .B(n1603), .Y(top_core_io_N493) );
  NOR2X1 U21365 ( .A(n4280), .B(n1602), .Y(top_core_io_N492) );
  NOR2X1 U21366 ( .A(n4279), .B(n1602), .Y(top_core_io_N491) );
  NOR2X1 U21367 ( .A(n4294), .B(n1602), .Y(top_core_io_N490) );
  NOR2X1 U21368 ( .A(n4293), .B(n1602), .Y(top_core_io_N489) );
  NOR2X1 U21369 ( .A(n4292), .B(n1602), .Y(top_core_io_N488) );
  NOR2X1 U21370 ( .A(n4291), .B(n1602), .Y(top_core_io_N487) );
  NOR2X1 U21371 ( .A(n4290), .B(n1602), .Y(top_core_io_N486) );
  NOR2X1 U21372 ( .A(n4289), .B(n1602), .Y(top_core_io_N485) );
  NOR2X1 U21373 ( .A(n4288), .B(n1602), .Y(top_core_io_N484) );
  NOR2X1 U21374 ( .A(n4287), .B(n1602), .Y(top_core_io_N483) );
  NOR2X1 U21375 ( .A(n4302), .B(n1602), .Y(top_core_io_N482) );
  NOR2X1 U21376 ( .A(n4301), .B(n1602), .Y(top_core_io_N481) );
  NOR2X1 U21377 ( .A(n4300), .B(n1602), .Y(top_core_io_N480) );
  NOR2X1 U21378 ( .A(n4299), .B(n1601), .Y(top_core_io_N479) );
  NOR2X1 U21379 ( .A(n4298), .B(n1601), .Y(top_core_io_N478) );
  NOR2X1 U21380 ( .A(n4297), .B(n1601), .Y(top_core_io_N477) );
  NOR2X1 U21381 ( .A(n4296), .B(n1601), .Y(top_core_io_N476) );
  NOR2X1 U21382 ( .A(n4295), .B(n1601), .Y(top_core_io_N475) );
  NOR2X1 U21383 ( .A(n4310), .B(n1601), .Y(top_core_io_N474) );
  NOR2X1 U21384 ( .A(n4309), .B(n1601), .Y(top_core_io_N473) );
  NOR2X1 U21385 ( .A(n4308), .B(n1601), .Y(top_core_io_N472) );
  NOR2X1 U21386 ( .A(n4307), .B(n1601), .Y(top_core_io_N471) );
  NOR2X1 U21387 ( .A(n4306), .B(n1601), .Y(top_core_io_N470) );
  NOR2X1 U21388 ( .A(n4305), .B(n1601), .Y(top_core_io_N469) );
  NOR2X1 U21389 ( .A(n4304), .B(n1601), .Y(top_core_io_N468) );
  NOR2X1 U21390 ( .A(n4303), .B(n1601), .Y(top_core_io_N467) );
  NOR2X1 U21391 ( .A(n4318), .B(n1592), .Y(top_core_io_N466) );
  NOR2X1 U21392 ( .A(n4317), .B(n1586), .Y(top_core_io_N465) );
  NOR2X1 U21393 ( .A(n4316), .B(n1583), .Y(top_core_io_N464) );
  NOR2X1 U21394 ( .A(n4315), .B(n1601), .Y(top_core_io_N463) );
  NOR2X1 U21395 ( .A(n4314), .B(n1588), .Y(top_core_io_N462) );
  NOR2X1 U21396 ( .A(n4313), .B(n1591), .Y(top_core_io_N461) );
  NOR2X1 U21397 ( .A(n4312), .B(n1590), .Y(top_core_io_N460) );
  NOR2X1 U21398 ( .A(n4311), .B(n1599), .Y(top_core_io_N459) );
  NOR2X1 U21399 ( .A(n4326), .B(n1597), .Y(top_core_io_N458) );
  NOR2X1 U21400 ( .A(n4325), .B(n1596), .Y(top_core_io_N457) );
  NOR2X1 U21401 ( .A(n4324), .B(n1598), .Y(top_core_io_N456) );
  NOR2X1 U21402 ( .A(n4323), .B(n1595), .Y(top_core_io_N455) );
  NOR2X1 U21403 ( .A(n4322), .B(n1594), .Y(top_core_io_N454) );
  NOR2X1 U21404 ( .A(n4321), .B(n1600), .Y(top_core_io_N453) );
  NOR2X1 U21405 ( .A(n4320), .B(n1600), .Y(top_core_io_N452) );
  NOR2X1 U21406 ( .A(n4319), .B(n1600), .Y(top_core_io_N451) );
  NOR2X1 U21407 ( .A(n4334), .B(n1600), .Y(top_core_io_N450) );
  NOR2X1 U21408 ( .A(n4333), .B(n1600), .Y(top_core_io_N449) );
  NOR2X1 U21409 ( .A(n4332), .B(n1600), .Y(top_core_io_N448) );
  NOR2X1 U21410 ( .A(n4331), .B(n1600), .Y(top_core_io_N447) );
  NOR2X1 U21411 ( .A(n4330), .B(n1600), .Y(top_core_io_N446) );
  NOR2X1 U21412 ( .A(n4329), .B(n1600), .Y(top_core_io_N445) );
  NOR2X1 U21413 ( .A(n4328), .B(n1600), .Y(top_core_io_N444) );
  NOR2X1 U21414 ( .A(n4327), .B(n1600), .Y(top_core_io_N443) );
  NOR2X1 U21415 ( .A(n4342), .B(n1600), .Y(top_core_io_N442) );
  NOR2X1 U21416 ( .A(n4341), .B(n1600), .Y(top_core_io_N441) );
  NOR2X1 U21417 ( .A(n4340), .B(n1599), .Y(top_core_io_N440) );
  NOR2X1 U21418 ( .A(n4339), .B(n1599), .Y(top_core_io_N439) );
  NOR2X1 U21419 ( .A(n4338), .B(n1599), .Y(top_core_io_N438) );
  NOR2X1 U21420 ( .A(n4337), .B(n1599), .Y(top_core_io_N437) );
  NOR2X1 U21421 ( .A(n4336), .B(n1599), .Y(top_core_io_N436) );
  NOR2X1 U21422 ( .A(n4335), .B(n1599), .Y(top_core_io_N435) );
  NOR2X1 U21423 ( .A(n4350), .B(n1599), .Y(top_core_io_N434) );
  NOR2X1 U21424 ( .A(n4349), .B(n1599), .Y(top_core_io_N433) );
  NOR2X1 U21425 ( .A(n4348), .B(n1599), .Y(top_core_io_N432) );
  NOR2X1 U21426 ( .A(n4347), .B(n1599), .Y(top_core_io_N431) );
  NOR2X1 U21427 ( .A(n4346), .B(n1599), .Y(top_core_io_N430) );
  NOR2X1 U21428 ( .A(n4345), .B(n1599), .Y(top_core_io_N429) );
  NOR2X1 U21429 ( .A(n4344), .B(n1599), .Y(top_core_io_N428) );
  NOR2X1 U21430 ( .A(n4343), .B(n1598), .Y(top_core_io_N427) );
  NOR2X1 U21431 ( .A(n4358), .B(n1598), .Y(top_core_io_N426) );
  NOR2X1 U21432 ( .A(n4357), .B(n1598), .Y(top_core_io_N425) );
  NOR2X1 U21433 ( .A(n4356), .B(n1598), .Y(top_core_io_N424) );
  NOR2X1 U21434 ( .A(n4355), .B(n1598), .Y(top_core_io_N423) );
  NOR2X1 U21435 ( .A(n4354), .B(n1598), .Y(top_core_io_N422) );
  NOR2X1 U21436 ( .A(n4353), .B(n1598), .Y(top_core_io_N421) );
  NOR2X1 U21437 ( .A(n4352), .B(n1598), .Y(top_core_io_N420) );
  NOR2X1 U21438 ( .A(n4351), .B(n1598), .Y(top_core_io_N419) );
  NOR2X1 U21439 ( .A(n4366), .B(n1598), .Y(top_core_io_N418) );
  NOR2X1 U21440 ( .A(n4365), .B(n1598), .Y(top_core_io_N417) );
  NOR2X1 U21441 ( .A(n4364), .B(n1598), .Y(top_core_io_N416) );
  NOR2X1 U21442 ( .A(n4363), .B(n1598), .Y(top_core_io_N415) );
  NOR2X1 U21443 ( .A(n4362), .B(n1597), .Y(top_core_io_N414) );
  NOR2X1 U21444 ( .A(n4361), .B(n1597), .Y(top_core_io_N413) );
  NOR2X1 U21445 ( .A(n4360), .B(n1597), .Y(top_core_io_N412) );
  NOR2X1 U21446 ( .A(n4359), .B(n1597), .Y(top_core_io_N411) );
  NOR2X1 U21447 ( .A(n4374), .B(n1597), .Y(top_core_io_N410) );
  NOR2X1 U21448 ( .A(n4373), .B(n1597), .Y(top_core_io_N409) );
  NOR2X1 U21449 ( .A(n4372), .B(n1597), .Y(top_core_io_N408) );
  NOR2X1 U21450 ( .A(n4371), .B(n1597), .Y(top_core_io_N407) );
  NOR2X1 U21451 ( .A(n4370), .B(n1597), .Y(top_core_io_N406) );
  NOR2X1 U21452 ( .A(n4369), .B(n1597), .Y(top_core_io_N405) );
  NOR2X1 U21453 ( .A(n4368), .B(n1597), .Y(top_core_io_N404) );
  NOR2X1 U21454 ( .A(n4367), .B(n1597), .Y(top_core_io_N403) );
  NOR2X1 U21455 ( .A(n4382), .B(n1597), .Y(top_core_io_N402) );
  NOR2X1 U21456 ( .A(n4381), .B(n1596), .Y(top_core_io_N401) );
  NOR2X1 U21457 ( .A(n4380), .B(n1596), .Y(top_core_io_N400) );
  NOR2X1 U21458 ( .A(n4379), .B(n1596), .Y(top_core_io_N399) );
  NOR2X1 U21459 ( .A(n4378), .B(n1596), .Y(top_core_io_N398) );
  NOR2X1 U21460 ( .A(n4377), .B(n1596), .Y(top_core_io_N397) );
  NOR2X1 U21461 ( .A(n4376), .B(n1596), .Y(top_core_io_N396) );
  NOR2X1 U21462 ( .A(n4375), .B(n1596), .Y(top_core_io_N395) );
  NOR2X1 U21463 ( .A(n4390), .B(n1596), .Y(top_core_io_N394) );
  NOR2X1 U21464 ( .A(n4389), .B(n1596), .Y(top_core_io_N393) );
  NOR2X1 U21465 ( .A(n4388), .B(n1596), .Y(top_core_io_N392) );
  NOR2X1 U21466 ( .A(n4387), .B(n1596), .Y(top_core_io_N391) );
  NOR2X1 U21467 ( .A(n4386), .B(n1596), .Y(top_core_io_N390) );
  NOR2X1 U21468 ( .A(n4385), .B(n1596), .Y(top_core_io_N389) );
  NOR2X1 U21469 ( .A(n4384), .B(n1595), .Y(top_core_io_N388) );
  NOR2X1 U21470 ( .A(n4383), .B(n1595), .Y(top_core_io_N387) );
  NOR2X1 U21471 ( .A(n4398), .B(n1595), .Y(top_core_io_N386) );
  NOR2X1 U21472 ( .A(n4397), .B(n1595), .Y(top_core_io_N385) );
  NOR2X1 U21473 ( .A(n4396), .B(n1595), .Y(top_core_io_N384) );
  NOR2X1 U21474 ( .A(n4395), .B(n1595), .Y(top_core_io_N383) );
  NOR2X1 U21475 ( .A(n4394), .B(n1595), .Y(top_core_io_N382) );
  NOR2X1 U21476 ( .A(n4393), .B(n1595), .Y(top_core_io_N381) );
  NOR2X1 U21477 ( .A(n4392), .B(n1595), .Y(top_core_io_N380) );
  NOR2X1 U21478 ( .A(n4391), .B(n1595), .Y(top_core_io_N379) );
  NOR2X1 U21479 ( .A(n4406), .B(n1595), .Y(top_core_io_N378) );
  NOR2X1 U21480 ( .A(n4405), .B(n1595), .Y(top_core_io_N377) );
  NOR2X1 U21481 ( .A(n4404), .B(n1595), .Y(top_core_io_N376) );
  NOR2X1 U21482 ( .A(n4403), .B(n1594), .Y(top_core_io_N375) );
  NOR2X1 U21483 ( .A(n4402), .B(n1594), .Y(top_core_io_N374) );
  NOR2X1 U21484 ( .A(n4401), .B(n1594), .Y(top_core_io_N373) );
  NOR2X1 U21485 ( .A(n4400), .B(n1594), .Y(top_core_io_N372) );
  NOR2X1 U21486 ( .A(n4399), .B(n1594), .Y(top_core_io_N371) );
  NOR2X1 U21487 ( .A(n4414), .B(n1594), .Y(top_core_io_N370) );
  NOR2X1 U21488 ( .A(n4413), .B(n1594), .Y(top_core_io_N369) );
  NOR2X1 U21489 ( .A(n4412), .B(n1594), .Y(top_core_io_N368) );
  NOR2X1 U21490 ( .A(n4411), .B(n1594), .Y(top_core_io_N367) );
  NOR2X1 U21491 ( .A(n4410), .B(n1594), .Y(top_core_io_N366) );
  NOR2X1 U21492 ( .A(n4409), .B(n1594), .Y(top_core_io_N365) );
  NOR2X1 U21493 ( .A(n4408), .B(n1594), .Y(top_core_io_N364) );
  NOR2X1 U21494 ( .A(n4407), .B(n1594), .Y(top_core_io_N363) );
  NOR2X1 U21495 ( .A(n4422), .B(n1587), .Y(top_core_io_N362) );
  NOR2X1 U21496 ( .A(n4421), .B(n1603), .Y(top_core_io_N361) );
  NOR2X1 U21497 ( .A(n4420), .B(n1602), .Y(top_core_io_N360) );
  NOR2X1 U21498 ( .A(n4419), .B(n4257), .Y(top_core_io_N359) );
  NOR2X1 U21499 ( .A(n4418), .B(n1600), .Y(top_core_io_N358) );
  NOR2X1 U21500 ( .A(n4417), .B(n1586), .Y(top_core_io_N357) );
  NOR2X1 U21501 ( .A(n4416), .B(n1583), .Y(top_core_io_N356) );
  NOR2X1 U21502 ( .A(n4415), .B(n1601), .Y(top_core_io_N355) );
  NOR2X1 U21503 ( .A(n4430), .B(n1588), .Y(top_core_io_N354) );
  NOR2X1 U21504 ( .A(n4429), .B(n1591), .Y(top_core_io_N353) );
  NOR2X1 U21505 ( .A(n4428), .B(n1590), .Y(top_core_io_N352) );
  NOR2X1 U21506 ( .A(n4427), .B(n1599), .Y(top_core_io_N351) );
  NOR2X1 U21507 ( .A(n4426), .B(n1597), .Y(top_core_io_N350) );
  NOR2X1 U21508 ( .A(n4425), .B(n4257), .Y(top_core_io_N349) );
  NOR2X1 U21509 ( .A(n4424), .B(n1598), .Y(top_core_io_N348) );
  NOR2X1 U21510 ( .A(n4423), .B(n1595), .Y(top_core_io_N347) );
  NOR2X1 U21511 ( .A(n4438), .B(n1594), .Y(top_core_io_N346) );
  NOR2X1 U21512 ( .A(n4437), .B(n1585), .Y(top_core_io_N345) );
  NOR2X1 U21513 ( .A(n4436), .B(n1584), .Y(top_core_io_N344) );
  NOR2X1 U21514 ( .A(n4435), .B(n1582), .Y(top_core_io_N343) );
  NOR2X1 U21515 ( .A(n4434), .B(n1604), .Y(top_core_io_N342) );
  NOR2X1 U21516 ( .A(n4433), .B(n1584), .Y(top_core_io_N341) );
  NOR2X1 U21517 ( .A(n4432), .B(n1604), .Y(top_core_io_N340) );
  NOR2X1 U21518 ( .A(n4431), .B(n1596), .Y(top_core_io_N339) );
  NOR2X1 U21519 ( .A(n4446), .B(n1593), .Y(top_core_io_N338) );
  NOR2X1 U21520 ( .A(n4445), .B(n1592), .Y(top_core_io_N337) );
  NOR2X1 U21521 ( .A(n4444), .B(n1593), .Y(top_core_io_N336) );
  NOR2X1 U21522 ( .A(n4443), .B(n1593), .Y(top_core_io_N335) );
  NOR2X1 U21523 ( .A(n4442), .B(n1593), .Y(top_core_io_N334) );
  NOR2X1 U21524 ( .A(n4441), .B(n1593), .Y(top_core_io_N333) );
  NOR2X1 U21525 ( .A(n4440), .B(n1593), .Y(top_core_io_N332) );
  NOR2X1 U21526 ( .A(n4439), .B(n1593), .Y(top_core_io_N331) );
  NOR2X1 U21527 ( .A(n4454), .B(n1593), .Y(top_core_io_N330) );
  NOR2X1 U21528 ( .A(n4453), .B(n1593), .Y(top_core_io_N329) );
  NOR2X1 U21529 ( .A(n4452), .B(n1593), .Y(top_core_io_N328) );
  NOR2X1 U21530 ( .A(n4451), .B(n1593), .Y(top_core_io_N327) );
  NOR2X1 U21531 ( .A(n4450), .B(n1593), .Y(top_core_io_N326) );
  NOR2X1 U21532 ( .A(n4449), .B(n1593), .Y(top_core_io_N325) );
  NOR2X1 U21533 ( .A(n4448), .B(n1593), .Y(top_core_io_N324) );
  NOR2X1 U21534 ( .A(n4447), .B(n1592), .Y(top_core_io_N323) );
  NOR2X1 U21535 ( .A(n4462), .B(n1592), .Y(top_core_io_N322) );
  NOR2X1 U21536 ( .A(n4461), .B(n1592), .Y(top_core_io_N321) );
  NOR2X1 U21537 ( .A(n4460), .B(n1592), .Y(top_core_io_N320) );
  NOR2X1 U21538 ( .A(n4459), .B(n1592), .Y(top_core_io_N319) );
  NOR2X1 U21539 ( .A(n4458), .B(n1592), .Y(top_core_io_N318) );
  NOR2X1 U21540 ( .A(n4457), .B(n1592), .Y(top_core_io_N317) );
  NOR2X1 U21541 ( .A(n4456), .B(n1592), .Y(top_core_io_N316) );
  NOR2X1 U21542 ( .A(n4455), .B(n1592), .Y(top_core_io_N315) );
  NOR2X1 U21543 ( .A(n4470), .B(n1592), .Y(top_core_io_N314) );
  NOR2X1 U21544 ( .A(n4469), .B(n1592), .Y(top_core_io_N313) );
  NOR2X1 U21545 ( .A(n4468), .B(n1592), .Y(top_core_io_N312) );
  NOR2X1 U21546 ( .A(n4467), .B(n1592), .Y(top_core_io_N311) );
  NOR2X1 U21547 ( .A(n4466), .B(n1591), .Y(top_core_io_N310) );
  NOR2X1 U21548 ( .A(n4465), .B(n1591), .Y(top_core_io_N309) );
  NOR2X1 U21549 ( .A(n4464), .B(n1591), .Y(top_core_io_N308) );
  NOR2X1 U21550 ( .A(n4463), .B(n1591), .Y(top_core_io_N307) );
  NOR2X1 U21551 ( .A(n4478), .B(n1591), .Y(top_core_io_N306) );
  NOR2X1 U21552 ( .A(n4477), .B(n1591), .Y(top_core_io_N305) );
  NOR2X1 U21553 ( .A(n4476), .B(n1591), .Y(top_core_io_N304) );
  NOR2X1 U21554 ( .A(n4475), .B(n1591), .Y(top_core_io_N303) );
  NOR2X1 U21555 ( .A(n4474), .B(n1591), .Y(top_core_io_N302) );
  NOR2X1 U21556 ( .A(n4473), .B(n1591), .Y(top_core_io_N301) );
  NOR2X1 U21557 ( .A(n4472), .B(n1591), .Y(top_core_io_N300) );
  NOR2X1 U21558 ( .A(n4471), .B(n1591), .Y(top_core_io_N299) );
  NOR2X1 U21559 ( .A(n4486), .B(n1591), .Y(top_core_io_N298) );
  NOR2X1 U21560 ( .A(n4485), .B(n1590), .Y(top_core_io_N297) );
  NOR2X1 U21561 ( .A(n4484), .B(n1590), .Y(top_core_io_N296) );
  NOR2X1 U21562 ( .A(n4483), .B(n1590), .Y(top_core_io_N295) );
  NOR2X1 U21563 ( .A(n4482), .B(n1590), .Y(top_core_io_N294) );
  NOR2X1 U21564 ( .A(n4481), .B(n1590), .Y(top_core_io_N293) );
  NOR2X1 U21565 ( .A(n4480), .B(n1590), .Y(top_core_io_N292) );
  NOR2X1 U21566 ( .A(n4479), .B(n1590), .Y(top_core_io_N291) );
  NOR2X1 U21567 ( .A(n4494), .B(n1590), .Y(top_core_io_N290) );
  NOR2X1 U21568 ( .A(n4493), .B(n1590), .Y(top_core_io_N289) );
  NOR2X1 U21569 ( .A(n4492), .B(n1590), .Y(top_core_io_N288) );
  NOR2X1 U21570 ( .A(n4491), .B(n1590), .Y(top_core_io_N287) );
  NOR2X1 U21571 ( .A(n4490), .B(n1590), .Y(top_core_io_N286) );
  NOR2X1 U21572 ( .A(n4489), .B(n1590), .Y(top_core_io_N285) );
  NOR2X1 U21573 ( .A(n4488), .B(n1587), .Y(top_core_io_N284) );
  NOR2X1 U21574 ( .A(n4487), .B(n1603), .Y(top_core_io_N283) );
  NOR2X1 U21575 ( .A(n4502), .B(n1602), .Y(top_core_io_N282) );
  NOR2X1 U21576 ( .A(n4501), .B(n1593), .Y(top_core_io_N281) );
  NOR2X1 U21577 ( .A(n4500), .B(n1600), .Y(top_core_io_N280) );
  NOR2X1 U21578 ( .A(n4499), .B(n1586), .Y(top_core_io_N279) );
  NOR2X1 U21579 ( .A(n4498), .B(n1583), .Y(top_core_io_N278) );
  NOR2X1 U21580 ( .A(n4497), .B(n1601), .Y(top_core_io_N277) );
  NOR2X1 U21581 ( .A(n4496), .B(n1588), .Y(top_core_io_N276) );
  NOR2X1 U21582 ( .A(n4495), .B(n1591), .Y(top_core_io_N275) );
  NOR2X1 U21583 ( .A(n4510), .B(n1590), .Y(top_core_io_N274) );
  NOR2X1 U21584 ( .A(n4509), .B(n1599), .Y(top_core_io_N273) );
  NOR2X1 U21585 ( .A(n4508), .B(n1597), .Y(top_core_io_N272) );
  NOR2X1 U21586 ( .A(n4507), .B(n1589), .Y(top_core_io_N271) );
  NOR2X1 U21587 ( .A(n4506), .B(n1589), .Y(top_core_io_N270) );
  NOR2X1 U21588 ( .A(n4505), .B(n1589), .Y(top_core_io_N269) );
  NOR2X1 U21589 ( .A(n4504), .B(n1589), .Y(top_core_io_N268) );
  NOR2X1 U21590 ( .A(n4503), .B(n1589), .Y(top_core_io_N267) );
  NOR2X1 U21591 ( .A(n4518), .B(n1589), .Y(top_core_io_N266) );
  NOR2X1 U21592 ( .A(n4517), .B(n1589), .Y(top_core_io_N265) );
  NOR2X1 U21593 ( .A(n4516), .B(n1589), .Y(top_core_io_N264) );
  NOR2X1 U21594 ( .A(n4515), .B(n1589), .Y(top_core_io_N263) );
  NOR2X1 U21595 ( .A(n4514), .B(n1589), .Y(top_core_io_N262) );
  NOR2X1 U21596 ( .A(n4513), .B(n1589), .Y(top_core_io_N261) );
  NOR2X1 U21597 ( .A(n4512), .B(n1589), .Y(top_core_io_N260) );
  NOR2X1 U21598 ( .A(n4511), .B(n1589), .Y(top_core_io_N259) );
  NOR2X1 U21599 ( .A(n4654), .B(n1588), .Y(top_core_io_N258) );
  NOR2X1 U21600 ( .A(n4653), .B(n1588), .Y(top_core_io_N257) );
  NOR2X1 U21601 ( .A(n4652), .B(n1588), .Y(top_core_io_N256) );
  NOR2X1 U21602 ( .A(n4651), .B(n1588), .Y(top_core_io_N255) );
  NOR2X1 U21603 ( .A(n4650), .B(n1588), .Y(top_core_io_N254) );
  NOR2X1 U21604 ( .A(n4649), .B(n1588), .Y(top_core_io_N253) );
  NOR2X1 U21605 ( .A(n4648), .B(n1588), .Y(top_core_io_N252) );
  NOR2X1 U21606 ( .A(n4647), .B(n1588), .Y(top_core_io_N251) );
  NOR2X1 U21607 ( .A(n4662), .B(n1588), .Y(top_core_io_N250) );
  NOR2X1 U21608 ( .A(n4661), .B(n1588), .Y(top_core_io_N249) );
  NOR2X1 U21609 ( .A(n4660), .B(n1588), .Y(top_core_io_N248) );
  NOR2X1 U21610 ( .A(n4659), .B(n1588), .Y(top_core_io_N247) );
  NOR2X1 U21611 ( .A(n4658), .B(n1588), .Y(top_core_io_N246) );
  NOR2X1 U21612 ( .A(n4657), .B(n4257), .Y(top_core_io_N245) );
  NOR2X1 U21613 ( .A(n4656), .B(n1586), .Y(top_core_io_N244) );
  NOR2X1 U21614 ( .A(n4655), .B(n1583), .Y(top_core_io_N243) );
  NOR2X1 U21615 ( .A(n4670), .B(n1601), .Y(top_core_io_N242) );
  NOR2X1 U21616 ( .A(n4669), .B(n1588), .Y(top_core_io_N241) );
  NOR2X1 U21617 ( .A(n4668), .B(n1591), .Y(top_core_io_N240) );
  NOR2X1 U21618 ( .A(n4667), .B(n1590), .Y(top_core_io_N239) );
  NOR2X1 U21619 ( .A(n4666), .B(n1599), .Y(top_core_io_N238) );
  NOR2X1 U21620 ( .A(n4665), .B(n1597), .Y(top_core_io_N237) );
  NOR2X1 U21621 ( .A(n4664), .B(n1596), .Y(top_core_io_N236) );
  NOR2X1 U21622 ( .A(n4663), .B(n1598), .Y(top_core_io_N235) );
  NOR2X1 U21623 ( .A(n4678), .B(n1595), .Y(top_core_io_N234) );
  NOR2X1 U21624 ( .A(n4677), .B(n1594), .Y(top_core_io_N233) );
  NOR2X1 U21625 ( .A(n4676), .B(n1587), .Y(top_core_io_N232) );
  NOR2X1 U21626 ( .A(n4675), .B(n1587), .Y(top_core_io_N231) );
  NOR2X1 U21627 ( .A(n4674), .B(n1587), .Y(top_core_io_N230) );
  NOR2X1 U21628 ( .A(n4673), .B(n1587), .Y(top_core_io_N229) );
  NOR2X1 U21629 ( .A(n4672), .B(n1587), .Y(top_core_io_N228) );
  NOR2X1 U21630 ( .A(n4671), .B(n1587), .Y(top_core_io_N227) );
  NOR2X1 U21631 ( .A(n4686), .B(n1587), .Y(top_core_io_N226) );
  NOR2X1 U21632 ( .A(n4685), .B(n1587), .Y(top_core_io_N225) );
  NOR2X1 U21633 ( .A(n4684), .B(n1587), .Y(top_core_io_N224) );
  NOR2X1 U21634 ( .A(n4683), .B(n1587), .Y(top_core_io_N223) );
  NOR2X1 U21635 ( .A(n4682), .B(n1587), .Y(top_core_io_N222) );
  NOR2X1 U21636 ( .A(n4681), .B(n1587), .Y(top_core_io_N221) );
  NOR2X1 U21637 ( .A(n4680), .B(n1587), .Y(top_core_io_N220) );
  NOR2X1 U21638 ( .A(n4679), .B(n1586), .Y(top_core_io_N219) );
  NOR2X1 U21639 ( .A(n4694), .B(n1586), .Y(top_core_io_N218) );
  NOR2X1 U21640 ( .A(n4693), .B(n1586), .Y(top_core_io_N217) );
  NOR2X1 U21641 ( .A(n4692), .B(n1586), .Y(top_core_io_N216) );
  NOR2X1 U21642 ( .A(n4691), .B(n1586), .Y(top_core_io_N215) );
  NOR2X1 U21643 ( .A(n4690), .B(n1586), .Y(top_core_io_N214) );
  NOR2X1 U21644 ( .A(n4689), .B(n1586), .Y(top_core_io_N213) );
  NOR2X1 U21645 ( .A(n4688), .B(n1586), .Y(top_core_io_N212) );
  NOR2X1 U21646 ( .A(n4687), .B(n1586), .Y(top_core_io_N211) );
  NOR2X1 U21647 ( .A(n4702), .B(n1586), .Y(top_core_io_N210) );
  NOR2X1 U21648 ( .A(n4701), .B(n1586), .Y(top_core_io_N209) );
  NOR2X1 U21649 ( .A(n4700), .B(n1586), .Y(top_core_io_N208) );
  NOR2X1 U21650 ( .A(n4699), .B(n1586), .Y(top_core_io_N207) );
  NOR2X1 U21651 ( .A(n4698), .B(n1585), .Y(top_core_io_N206) );
  NOR2X1 U21652 ( .A(n4697), .B(n1585), .Y(top_core_io_N205) );
  NOR2X1 U21653 ( .A(n4696), .B(n1585), .Y(top_core_io_N204) );
  NOR2X1 U21654 ( .A(n4695), .B(n1585), .Y(top_core_io_N203) );
  NOR2X1 U21655 ( .A(n4710), .B(n1585), .Y(top_core_io_N202) );
  NOR2X1 U21656 ( .A(n4709), .B(n1585), .Y(top_core_io_N201) );
  NOR2X1 U21657 ( .A(n4708), .B(n1585), .Y(top_core_io_N200) );
  NOR2X1 U21658 ( .A(n4707), .B(n1585), .Y(top_core_io_N199) );
  NOR2X1 U21659 ( .A(n4706), .B(n1585), .Y(top_core_io_N198) );
  NOR2X1 U21660 ( .A(n4705), .B(n1585), .Y(top_core_io_N197) );
  NOR2X1 U21661 ( .A(n4704), .B(n1585), .Y(top_core_io_N196) );
  NOR2X1 U21662 ( .A(n4703), .B(n1585), .Y(top_core_io_N195) );
  NOR2X1 U21663 ( .A(n4718), .B(n1585), .Y(top_core_io_N194) );
  NOR2X1 U21664 ( .A(n4717), .B(n1584), .Y(top_core_io_N193) );
  NOR2X1 U21665 ( .A(n4716), .B(n1584), .Y(top_core_io_N192) );
  NOR2X1 U21666 ( .A(n4715), .B(n1584), .Y(top_core_io_N191) );
  NOR2X1 U21667 ( .A(n4714), .B(n1584), .Y(top_core_io_N190) );
  NOR2X1 U21668 ( .A(n4713), .B(n1584), .Y(top_core_io_N189) );
  NOR2X1 U21669 ( .A(n4712), .B(n1584), .Y(top_core_io_N188) );
  NOR2X1 U21670 ( .A(n4711), .B(n1584), .Y(top_core_io_N187) );
  NOR2X1 U21671 ( .A(n4726), .B(n1584), .Y(top_core_io_N186) );
  NOR2X1 U21672 ( .A(n4725), .B(n1584), .Y(top_core_io_N185) );
  NOR2X1 U21673 ( .A(n4724), .B(n1584), .Y(top_core_io_N184) );
  NOR2X1 U21674 ( .A(n4723), .B(n1584), .Y(top_core_io_N183) );
  NOR2X1 U21675 ( .A(n4722), .B(n1584), .Y(top_core_io_N182) );
  NOR2X1 U21676 ( .A(n4721), .B(n1584), .Y(top_core_io_N181) );
  NOR2X1 U21677 ( .A(n4720), .B(n1595), .Y(top_core_io_N180) );
  NOR2X1 U21678 ( .A(n4719), .B(n1594), .Y(top_core_io_N179) );
  NOR2X1 U21679 ( .A(n4734), .B(n1585), .Y(top_core_io_N178) );
  NOR2X1 U21680 ( .A(n4733), .B(n1584), .Y(top_core_io_N177) );
  NOR2X1 U21681 ( .A(n4732), .B(n1582), .Y(top_core_io_N176) );
  NOR2X1 U21682 ( .A(n4731), .B(n1604), .Y(top_core_io_N175) );
  NOR2X1 U21683 ( .A(n4730), .B(n1585), .Y(top_core_io_N174) );
  NOR2X1 U21684 ( .A(n4729), .B(n1593), .Y(top_core_io_N173) );
  NOR2X1 U21685 ( .A(n4728), .B(n1592), .Y(top_core_io_N172) );
  NOR2X1 U21686 ( .A(n4727), .B(n1589), .Y(top_core_io_N171) );
  NOR2X1 U21687 ( .A(n4742), .B(n1587), .Y(top_core_io_N170) );
  NOR2X1 U21688 ( .A(n4741), .B(n1603), .Y(top_core_io_N169) );
  NOR2X1 U21689 ( .A(n4740), .B(n1602), .Y(top_core_io_N168) );
  NOR2X1 U21690 ( .A(n4739), .B(n4257), .Y(top_core_io_N167) );
  NOR2X1 U21691 ( .A(n4738), .B(n4257), .Y(top_core_io_N166) );
  NOR2X1 U21692 ( .A(n4737), .B(n1604), .Y(top_core_io_N165) );
  NOR2X1 U21693 ( .A(n4736), .B(n1604), .Y(top_core_io_N164) );
  NOR2X1 U21694 ( .A(n4735), .B(n1604), .Y(top_core_io_N163) );
  NOR2X1 U21695 ( .A(n4750), .B(n1582), .Y(top_core_io_N162) );
  NOR2X1 U21696 ( .A(n4749), .B(n1600), .Y(top_core_io_N161) );
  NOR2X1 U21697 ( .A(n4748), .B(n1598), .Y(top_core_io_N160) );
  NOR2X1 U21698 ( .A(n4747), .B(n1589), .Y(top_core_io_N159) );
  NOR2X1 U21699 ( .A(n4746), .B(n1596), .Y(top_core_io_N158) );
  NOR2X1 U21700 ( .A(n4745), .B(n1593), .Y(top_core_io_N157) );
  NOR2X1 U21701 ( .A(n4744), .B(n1592), .Y(top_core_io_N156) );
  NOR2X1 U21702 ( .A(n4743), .B(n1589), .Y(top_core_io_N155) );
  NOR2X1 U21703 ( .A(n4758), .B(n1583), .Y(top_core_io_N154) );
  NOR2X1 U21704 ( .A(n4757), .B(n1583), .Y(top_core_io_N153) );
  NOR2X1 U21705 ( .A(n4756), .B(n1583), .Y(top_core_io_N152) );
  NOR2X1 U21706 ( .A(n4755), .B(n1583), .Y(top_core_io_N151) );
  NOR2X1 U21707 ( .A(n4754), .B(n1583), .Y(top_core_io_N150) );
  NOR2X1 U21708 ( .A(n4753), .B(n1583), .Y(top_core_io_N149) );
  NOR2X1 U21709 ( .A(n4752), .B(n1583), .Y(top_core_io_N148) );
  NOR2X1 U21710 ( .A(n4751), .B(n1583), .Y(top_core_io_N147) );
  NOR2X1 U21711 ( .A(n4766), .B(n1583), .Y(top_core_io_N146) );
  NOR2X1 U21712 ( .A(n4765), .B(n1583), .Y(top_core_io_N145) );
  NOR2X1 U21713 ( .A(n4764), .B(n1583), .Y(top_core_io_N144) );
  NOR2X1 U21714 ( .A(n4763), .B(n1583), .Y(top_core_io_N143) );
  NOR2X1 U21715 ( .A(n4762), .B(n1583), .Y(top_core_io_N142) );
  NOR2X1 U21716 ( .A(n4278), .B(n1604), .Y(top_core_io_N506) );
  NOR2X1 U21717 ( .A(n4270), .B(n1604), .Y(top_core_io_N514) );
  NOR2X1 U21718 ( .A(n4269), .B(n1604), .Y(top_core_io_N513) );
  NOR2X1 U21719 ( .A(n4268), .B(n1604), .Y(top_core_io_N512) );
  NOR2X1 U21720 ( .A(n4267), .B(n1604), .Y(top_core_io_N511) );
  NOR2X1 U21721 ( .A(n4266), .B(n1604), .Y(top_core_io_N510) );
  NOR2X1 U21722 ( .A(n4265), .B(n1604), .Y(top_core_io_N509) );
  NOR2X1 U21723 ( .A(n4264), .B(n1604), .Y(top_core_io_N508) );
  NOR2X1 U21724 ( .A(n4263), .B(n1604), .Y(top_core_io_N507) );
  NOR2X1 U21725 ( .A(n4260), .B(n1604), .Y(top_core_io_N515) );
  INVX1 U21726 ( .A(n1344), .Y(n6964) );
  INVX1 U21727 ( .A(n1345), .Y(n6958) );
  INVX1 U21728 ( .A(n1359), .Y(n6670) );
  BUFX3 U21729 ( .A(n6651), .Y(n1168) );
  INVX1 U21730 ( .A(n1361), .Y(n6651) );
  BUFX3 U21731 ( .A(n6634), .Y(n1166) );
  INVX1 U21732 ( .A(n1363), .Y(n6634) );
  BUFX3 U21733 ( .A(n6941), .Y(n1208) );
  INVX1 U21734 ( .A(n1347), .Y(n6941) );
  BUFX3 U21735 ( .A(n6926), .Y(n1206) );
  INVX1 U21736 ( .A(n1349), .Y(n6926) );
  BUFX3 U21737 ( .A(n6949), .Y(n1209) );
  INVX1 U21738 ( .A(n1346), .Y(n6949) );
  BUFX3 U21739 ( .A(n6934), .Y(n1207) );
  INVX1 U21740 ( .A(n1348), .Y(n6934) );
  BUFX3 U21741 ( .A(n6643), .Y(n1167) );
  INVX1 U21742 ( .A(n1362), .Y(n6643) );
  OR3XL U21743 ( .A(top_core_KE_round_ctr_reg_0_), .B(n1334), .C(n7013), .Y(
        n743) );
  BUFX3 U21744 ( .A(n6659), .Y(n1169) );
  INVX1 U21745 ( .A(n1360), .Y(n6659) );
  AND2X2 U21746 ( .A(n1358), .B(n752), .Y(n744) );
  AND2X2 U21747 ( .A(n1344), .B(n753), .Y(n745) );
  AND2X2 U21748 ( .A(n1345), .B(n754), .Y(n746) );
  AND2X2 U21749 ( .A(n1359), .B(n755), .Y(n747) );
  BUFX3 U21750 ( .A(n6599), .Y(n1159) );
  INVX1 U21751 ( .A(n1365), .Y(n6599) );
  BUFX3 U21752 ( .A(n6430), .Y(n1146) );
  INVX1 U21753 ( .A(n1369), .Y(n6430) );
  BUFX3 U21754 ( .A(n6551), .Y(n1150) );
  INVX1 U21755 ( .A(n1367), .Y(n6551) );
  BUFX3 U21756 ( .A(n6892), .Y(n1199) );
  INVX1 U21757 ( .A(n1351), .Y(n6892) );
  BUFX3 U21758 ( .A(n6846), .Y(n1190) );
  INVX1 U21759 ( .A(n1353), .Y(n6846) );
  BUFX3 U21760 ( .A(n6700), .Y(n1185) );
  INVX1 U21761 ( .A(n1356), .Y(n6700) );
  BUFX3 U21762 ( .A(n6711), .Y(n1186) );
  INVX1 U21763 ( .A(n1355), .Y(n6711) );
  BUFX3 U21764 ( .A(n6987), .Y(n1225) );
  INVX1 U21765 ( .A(n1342), .Y(n6987) );
  BUFX3 U21766 ( .A(n6742), .Y(n1187) );
  INVX1 U21767 ( .A(n1354), .Y(n6742) );
  BUFX3 U21768 ( .A(n6985), .Y(n1224) );
  INVX1 U21769 ( .A(n1343), .Y(n6985) );
  BUFX3 U21770 ( .A(n6698), .Y(n1184) );
  INVX1 U21771 ( .A(n1357), .Y(n6698) );
  BUFX3 U21772 ( .A(n6916), .Y(n1204) );
  INVX1 U21773 ( .A(n1350), .Y(n6916) );
  BUFX3 U21774 ( .A(n6870), .Y(n1195) );
  INVX1 U21775 ( .A(n1352), .Y(n6870) );
  BUFX3 U21776 ( .A(n6576), .Y(n1155) );
  INVX1 U21777 ( .A(n1366), .Y(n6576) );
  XNOR2X1 U21778 ( .A(top_core_KE_n1974), .B(top_core_KE_n2180), .Y(
        top_core_KE_n2178) );
  XNOR2X1 U21779 ( .A(top_core_KE_n2002), .B(top_core_KE_n2218), .Y(
        top_core_KE_n2217) );
  XNOR2X1 U21780 ( .A(top_core_KE_n1994), .B(top_core_KE_n2208), .Y(
        top_core_KE_n2207) );
  XNOR2X1 U21781 ( .A(top_core_KE_n1990), .B(top_core_KE_n2203), .Y(
        top_core_KE_n2202) );
  XNOR2X1 U21782 ( .A(top_core_KE_n1986), .B(top_core_KE_n2198), .Y(
        top_core_KE_n2197) );
  XNOR2X1 U21783 ( .A(top_core_KE_n1982), .B(top_core_KE_n2193), .Y(
        top_core_KE_n2192) );
  XNOR2X1 U21784 ( .A(top_core_KE_n1978), .B(top_core_KE_n2188), .Y(
        top_core_KE_n2187) );
  XNOR2X1 U21785 ( .A(top_core_KE_n1998), .B(top_core_KE_n2213), .Y(
        top_core_KE_n2212) );
  XOR2X1 U21786 ( .A(top_core_KE_n2213), .B(top_core_KE_n2379), .Y(
        top_core_KE_n2378) );
  XNOR2X1 U21787 ( .A(n1651), .B(top_core_KE_n1998), .Y(top_core_KE_n2379) );
  XOR2X1 U21788 ( .A(top_core_KE_n2303), .B(top_core_KE_n2471), .Y(
        top_core_KE_n2470) );
  XNOR2X1 U21789 ( .A(top_core_KE_new_sboxw_192_31_), .B(n1336), .Y(
        top_core_KE_n2471) );
  XOR2X1 U21790 ( .A(top_core_KE_n2263), .B(top_core_KE_n2431), .Y(
        top_core_KE_n2430) );
  XNOR2X1 U21791 ( .A(top_core_KE_new_sboxw_192_7_), .B(n1337), .Y(
        top_core_KE_n2431) );
  XOR2X1 U21792 ( .A(top_core_KE_n2223), .B(top_core_KE_n2391), .Y(
        top_core_KE_n2390) );
  XNOR2X1 U21793 ( .A(top_core_KE_new_sboxw_192_15_), .B(n1340), .Y(
        top_core_KE_n2391) );
  XOR2X1 U21794 ( .A(top_core_KE_n2180), .B(top_core_KE_n2343), .Y(
        top_core_KE_n2342) );
  XNOR2X1 U21795 ( .A(n1341), .B(top_core_KE_n1974), .Y(top_core_KE_n2343) );
  XOR2X1 U21796 ( .A(top_core_KE_n2308), .B(top_core_KE_n2476), .Y(
        top_core_KE_n2475) );
  XNOR2X1 U21797 ( .A(top_core_KE_new_sboxw_192_30_), .B(n1342), .Y(
        top_core_KE_n2476) );
  XOR2X1 U21798 ( .A(top_core_KE_n2283), .B(top_core_KE_n2451), .Y(
        top_core_KE_n2450) );
  XNOR2X1 U21799 ( .A(top_core_KE_new_sboxw_192_3_), .B(n1347), .Y(
        top_core_KE_n2451) );
  XOR2X1 U21800 ( .A(top_core_KE_n2323), .B(top_core_KE_n2491), .Y(
        top_core_KE_n2490) );
  XNOR2X1 U21801 ( .A(top_core_KE_new_sboxw_192_27_), .B(n1349), .Y(
        top_core_KE_n2491) );
  XOR2X1 U21802 ( .A(top_core_KE_n2278), .B(top_core_KE_n2446), .Y(
        top_core_KE_n2445) );
  XNOR2X1 U21803 ( .A(top_core_KE_new_sboxw_192_4_), .B(n1351), .Y(
        top_core_KE_n2446) );
  XOR2X1 U21804 ( .A(top_core_KE_n2318), .B(top_core_KE_n2486), .Y(
        top_core_KE_n2485) );
  XNOR2X1 U21805 ( .A(top_core_KE_new_sboxw_192_28_), .B(n1353), .Y(
        top_core_KE_n2486) );
  XOR2X1 U21806 ( .A(top_core_KE_n2268), .B(top_core_KE_n2436), .Y(
        top_core_KE_n2435) );
  XNOR2X1 U21807 ( .A(top_core_KE_new_sboxw_192_6_), .B(n1355), .Y(
        top_core_KE_n2436) );
  XOR2X1 U21808 ( .A(top_core_KE_n2228), .B(top_core_KE_n2396), .Y(
        top_core_KE_n2395) );
  XNOR2X1 U21809 ( .A(top_core_KE_new_sboxw_192_14_), .B(n1356), .Y(
        top_core_KE_n2396) );
  XOR2X1 U21810 ( .A(top_core_KE_n2218), .B(top_core_KE_n2385), .Y(
        top_core_KE_n2384) );
  XNOR2X1 U21811 ( .A(n1658), .B(top_core_KE_n2002), .Y(top_core_KE_n2385) );
  XOR2X1 U21812 ( .A(top_core_KE_n2208), .B(top_core_KE_n2373), .Y(
        top_core_KE_n2372) );
  XNOR2X1 U21813 ( .A(n1648), .B(top_core_KE_n1994), .Y(top_core_KE_n2373) );
  XOR2X1 U21814 ( .A(top_core_KE_n2203), .B(top_core_KE_n2367), .Y(
        top_core_KE_n2366) );
  XNOR2X1 U21815 ( .A(n1361), .B(top_core_KE_n1990), .Y(top_core_KE_n2367) );
  XOR2X1 U21816 ( .A(top_core_KE_n2243), .B(top_core_KE_n2411), .Y(
        top_core_KE_n2410) );
  XNOR2X1 U21817 ( .A(top_core_KE_new_sboxw_192_11_), .B(n1363), .Y(
        top_core_KE_n2411) );
  XOR2X1 U21818 ( .A(top_core_KE_n2198), .B(top_core_KE_n2361), .Y(
        top_core_KE_n2360) );
  XNOR2X1 U21819 ( .A(n1365), .B(top_core_KE_n1986), .Y(top_core_KE_n2361) );
  XOR2X1 U21820 ( .A(top_core_KE_n2238), .B(top_core_KE_n2406), .Y(
        top_core_KE_n2405) );
  XNOR2X1 U21821 ( .A(top_core_KE_new_sboxw_192_12_), .B(n1367), .Y(
        top_core_KE_n2406) );
  XOR2X1 U21822 ( .A(top_core_KE_n2193), .B(top_core_KE_n2355), .Y(
        top_core_KE_n2354) );
  XNOR2X1 U21823 ( .A(n1637), .B(top_core_KE_n1982), .Y(top_core_KE_n2355) );
  XOR2X1 U21824 ( .A(top_core_KE_n2188), .B(top_core_KE_n2349), .Y(
        top_core_KE_n2348) );
  XNOR2X1 U21825 ( .A(n1369), .B(top_core_KE_n1978), .Y(top_core_KE_n2349) );
  INVXL U21826 ( .A(n2), .Y(n4259) );
  INVX1 U21827 ( .A(n18877), .Y(n7009) );
  AOI21X1 U21828 ( .A0(top_core_KE_r343_u_div_PartRem_1__1_), .A1(
        top_core_KE_round_ctr_reg_0_), .B0(
        top_core_KE_r343_u_div_PartRem_1__2_), .Y(n18877) );
  MX2X1 U21829 ( .A(top_core_KE_r343_u_div_PartRem_2__1_), .B(
        top_core_KE_r343_u_div_SumTmp_1__1_), .S0(n7010), .Y(
        top_core_KE_r343_u_div_PartRem_1__2_) );
  XOR2X1 U21830 ( .A(n1332), .B(top_core_KE_r343_u_div_PartRem_2__1_), .Y(
        top_core_KE_r343_u_div_SumTmp_1__1_) );
  INVX1 U21831 ( .A(n18876), .Y(n7010) );
  AOI21X1 U21832 ( .A0(top_core_KE_r343_u_div_PartRem_2__1_), .A1(n1332), .B0(
        top_core_KE_r343_u_div_PartRem_2__2_), .Y(n18876) );
  MX2X1 U21833 ( .A(n1334), .B(top_core_KE_r343_u_div_SumTmp_2__1_), .S0(
        top_core_KE_r343_quotient_2_), .Y(top_core_KE_r343_u_div_PartRem_2__2_) );
  XOR2X1 U21834 ( .A(n1333), .B(n1334), .Y(top_core_KE_r343_u_div_SumTmp_2__1_) );
  AND2X2 U21835 ( .A(n1367), .B(n1166), .Y(n748) );
  AND2X2 U21836 ( .A(n1353), .B(n1206), .Y(n749) );
  AND2X2 U21837 ( .A(n1351), .B(n1208), .Y(n750) );
  AND2X2 U21838 ( .A(n1365), .B(n1168), .Y(n751) );
  AND2X2 U21839 ( .A(n1364), .B(n1169), .Y(n752) );
  AND2X2 U21840 ( .A(n1350), .B(n1209), .Y(n753) );
  AND2X2 U21841 ( .A(n1352), .B(n1207), .Y(n754) );
  AND2X2 U21842 ( .A(n1366), .B(n1167), .Y(n755) );
  AND2X2 U21843 ( .A(n1367), .B(n1363), .Y(n756) );
  AND2X2 U21844 ( .A(n1353), .B(n1349), .Y(n757) );
  AND2X2 U21845 ( .A(n1351), .B(n1347), .Y(n758) );
  AND2X2 U21846 ( .A(n1365), .B(n1361), .Y(n759) );
  AND2X2 U21847 ( .A(n1364), .B(n1360), .Y(n760) );
  AND2X2 U21848 ( .A(n1350), .B(n1346), .Y(n761) );
  AND2X2 U21849 ( .A(n1352), .B(n1348), .Y(n762) );
  AND2X2 U21850 ( .A(n1366), .B(n1362), .Y(n763) );
  BUFX3 U21851 ( .A(n7012), .Y(n1226) );
  INVX1 U21852 ( .A(n1333), .Y(n7012) );
  AOI211X1 U21853 ( .A0(n6919), .A1(n1814), .B0(n11731), .C0(n11732), .Y(
        n11729) );
  OAI21XL U21854 ( .A0(n11661), .A1(n11733), .B0(n11734), .Y(n11732) );
  AOI211X1 U21855 ( .A0(n6873), .A1(n1835), .B0(top_core_KE_sb1_n158), .C0(
        top_core_KE_sb1_n159), .Y(top_core_KE_sb1_n156) );
  OAI21XL U21856 ( .A0(top_core_KE_sb1_n86), .A1(top_core_KE_sb1_n160), .B0(
        top_core_KE_sb1_n161), .Y(top_core_KE_sb1_n159) );
  AOI211X1 U21857 ( .A0(n6626), .A1(n1773), .B0(n12362), .C0(n12363), .Y(
        n12360) );
  OAI21XL U21858 ( .A0(n1264), .A1(n12364), .B0(n12365), .Y(n12363) );
  AOI211X1 U21859 ( .A0(n6579), .A1(n1793), .B0(n12047), .C0(n12048), .Y(
        n12045) );
  OAI21XL U21860 ( .A0(n11977), .A1(n12049), .B0(n12050), .Y(n12048) );
  AOI211X1 U21861 ( .A0(n6849), .A1(n1748), .B0(n12678), .C0(n12679), .Y(
        n12676) );
  OAI21XL U21862 ( .A0(n12608), .A1(n12680), .B0(n12681), .Y(n12679) );
  AOI211X1 U21863 ( .A0(n6895), .A1(n1719), .B0(n12993), .C0(n12994), .Y(
        n12991) );
  OAI21XL U21864 ( .A0(n12923), .A1(n12995), .B0(n12996), .Y(n12994) );
  AOI211X1 U21865 ( .A0(n6602), .A1(n1660), .B0(n13623), .C0(n13624), .Y(
        n13621) );
  OAI21XL U21866 ( .A0(n13553), .A1(n13625), .B0(n13626), .Y(n13624) );
  BUFX3 U21867 ( .A(n6440), .Y(n1147) );
  INVX1 U21868 ( .A(n1368), .Y(n6440) );
  BUFX3 U21869 ( .A(n6623), .Y(n1164) );
  INVX1 U21870 ( .A(n1364), .Y(n6623) );
  OAI2BB1X1 U21871 ( .A0N(top_core_KE_n2714), .A1N(n1334), .B0(
        top_core_KE_n2715), .Y(top_core_KE_n4929) );
  OR4X2 U21872 ( .A(top_core_KE_n2716), .B(n1226), .C(n7014), .D(n1334), .Y(
        top_core_KE_n2715) );
  OAI21XL U21873 ( .A0(n7016), .A1(n1333), .B0(top_core_KE_n2717), .Y(
        top_core_KE_n2714) );
  AOI222X1 U21874 ( .A0(n6951), .A1(n1344), .B0(n11663), .B1(n681), .C0(n6917), 
        .C1(n1808), .Y(n11898) );
  AOI222X1 U21875 ( .A0(n6936), .A1(n1345), .B0(top_core_KE_sb1_n88), .B1(n682), .C0(n6871), .C1(n1829), .Y(top_core_KE_sb1_n327) );
  AOI222X1 U21876 ( .A0(n6661), .A1(n1358), .B0(n12294), .B1(n683), .C0(n6624), 
        .C1(n1765), .Y(n12529) );
  AOI222X1 U21877 ( .A0(n6645), .A1(n1359), .B0(n11979), .B1(n684), .C0(n6577), 
        .C1(n1787), .Y(n12214) );
  OAI32X1 U21878 ( .A0(top_core_KE_n2716), .A1(n1333), .A2(n7014), .B0(
        top_core_KE_n2717), .B1(n1226), .Y(top_core_KE_n4930) );
  OAI21XL U21879 ( .A0(n6587), .A1(n1160), .B0(n1663), .Y(n13607) );
  OAI21XL U21880 ( .A0(n6539), .A1(n1151), .B0(n1689), .Y(n13292) );
  OAI21XL U21881 ( .A0(n6834), .A1(n1191), .B0(n1747), .Y(n12662) );
  OAI21XL U21882 ( .A0(n6880), .A1(n1200), .B0(n1718), .Y(n12977) );
  OAI21XL U21883 ( .A0(n6904), .A1(n745), .B0(n1813), .Y(n11715) );
  OAI21XL U21884 ( .A0(n6858), .A1(n746), .B0(n1834), .Y(top_core_KE_sb1_n141)
         );
  OAI21XL U21885 ( .A0(n6564), .A1(n747), .B0(n1792), .Y(n12031) );
  OAI21XL U21886 ( .A0(n6611), .A1(n744), .B0(n1769), .Y(n12346) );
  INVX1 U21887 ( .A(top_core_io_n653), .Y(n4258) );
  INVX1 U21888 ( .A(top_core_KE_n903), .Y(n6342) );
  INVX1 U21889 ( .A(top_core_KE_n1056), .Y(n6730) );
  INVX1 U21890 ( .A(top_core_KE_n1112), .Y(n6793) );
  INVX1 U21891 ( .A(top_core_KE_n1035), .Y(n6724) );
  INVX1 U21892 ( .A(top_core_KE_n1091), .Y(n6782) );
  INVX1 U21893 ( .A(top_core_KE_n1077), .Y(n6378) );
  INVX1 U21894 ( .A(top_core_KE_n1021), .Y(n6329) );
  INVX1 U21895 ( .A(top_core_KE_n944), .Y(n6371) );
  INVX1 U21896 ( .A(top_core_KE_n923), .Y(n6363) );
  INVX1 U21897 ( .A(top_core_KE_n1070), .Y(n6741) );
  INVX1 U21898 ( .A(top_core_KE_n1126), .Y(n6798) );
  INVX1 U21899 ( .A(top_core_KE_n1028), .Y(n6718) );
  INVX1 U21900 ( .A(top_core_KE_n958), .Y(n6357) );
  INVX1 U21901 ( .A(top_core_KE_n913), .Y(n6349) );
  INVX1 U21902 ( .A(top_core_KE_n1084), .Y(n6385) );
  INVX1 U21903 ( .A(top_core_KE_n1063), .Y(n6738) );
  INVX1 U21904 ( .A(top_core_KE_n1119), .Y(n6796) );
  INVX1 U21905 ( .A(top_core_KE_n1049), .Y(n6734) );
  INVX1 U21906 ( .A(top_core_KE_n1105), .Y(n6791) );
  INVX1 U21907 ( .A(top_core_KE_n1042), .Y(n6727) );
  INVX1 U21908 ( .A(top_core_KE_n1098), .Y(n6789) );
  INVX1 U21909 ( .A(top_core_KE_n951), .Y(n6315) );
  INVX1 U21910 ( .A(top_core_KE_n937), .Y(n6367) );
  INVX1 U21911 ( .A(top_core_KE_n930), .Y(n6353) );
  INVX1 U21912 ( .A(top_core_KE_prev_key1_reg_85_), .Y(n1668) );
  INVX1 U21913 ( .A(top_core_KE_prev_key1_reg_69_), .Y(n1726) );
  INVX1 U21914 ( .A(top_core_KE_prev_key1_reg_77_), .Y(n1697) );
  INVX1 U21915 ( .A(n1650), .Y(n1645) );
  INVX1 U21916 ( .A(top_core_KE_prev_key1_reg_85_), .Y(n1669) );
  INVX1 U21917 ( .A(top_core_KE_prev_key1_reg_69_), .Y(n1727) );
  INVX1 U21918 ( .A(top_core_KE_prev_key1_reg_77_), .Y(n1698) );
  INVX1 U21919 ( .A(n1644), .Y(n1646) );
  INVX1 U21920 ( .A(top_core_KE_prev_key1_reg_85_), .Y(n1670) );
  INVX1 U21921 ( .A(top_core_KE_prev_key1_reg_69_), .Y(n1728) );
  INVX1 U21922 ( .A(top_core_KE_prev_key1_reg_77_), .Y(n1699) );
  INVX1 U21923 ( .A(n1796), .Y(n1797) );
  INVX1 U21924 ( .A(n1817), .Y(n1818) );
  INVX1 U21925 ( .A(n1775), .Y(n1776) );
  INVX1 U21926 ( .A(n1650), .Y(n1647) );
  INVX1 U21927 ( .A(n1753), .Y(n1754) );
  INVX1 U21928 ( .A(n1796), .Y(n1798) );
  INVX1 U21929 ( .A(n1817), .Y(n1819) );
  INVX1 U21930 ( .A(n1775), .Y(n1777) );
  INVX1 U21931 ( .A(n1650), .Y(n1648) );
  INVX1 U21932 ( .A(n1752), .Y(n1755) );
  INVX1 U21933 ( .A(n1642), .Y(n1637) );
  AND3X2 U21934 ( .A(n7015), .B(n7008), .C(top_core_KE_n2700), .Y(n764) );
  AND2X2 U21935 ( .A(top_core_KE_n1871), .B(top_core_KE_n894), .Y(n765) );
  AND2X2 U21936 ( .A(top_core_EC_n862), .B(top_core_EC_n861), .Y(n766) );
  NAND2BX1 U21937 ( .AN(top_core_EC_n861), .B(top_core_EC_n862), .Y(
        top_core_EC_n730) );
  INVX1 U21938 ( .A(top_core_KE_n2175), .Y(n2286) );
  INVX1 U21939 ( .A(top_core_EC_operation), .Y(n2540) );
  INVX1 U21940 ( .A(n1759), .Y(n1756) );
  INVX1 U21941 ( .A(n1650), .Y(n1649) );
  INVX1 U21942 ( .A(n1642), .Y(n1638) );
  INVX1 U21943 ( .A(n1759), .Y(n1757) );
  INVX1 U21944 ( .A(n1642), .Y(n1639) );
  INVX1 U21945 ( .A(n1795), .Y(n1799) );
  INVX1 U21946 ( .A(n1816), .Y(n1820) );
  INVX1 U21947 ( .A(n1774), .Y(n1778) );
  INVX1 U21948 ( .A(n1642), .Y(n1640) );
  INVX1 U21949 ( .A(n1795), .Y(n1800) );
  INVX1 U21950 ( .A(n1816), .Y(n1821) );
  INVX1 U21951 ( .A(n1774), .Y(n1779) );
  INVX1 U21952 ( .A(n4034), .Y(n4033) );
  INVX1 U21953 ( .A(n4095), .Y(n4031) );
  INVX1 U21954 ( .A(n4034), .Y(n4032) );
  INVX1 U21955 ( .A(n1795), .Y(n1801) );
  INVX1 U21956 ( .A(n1816), .Y(n1822) );
  INVX1 U21957 ( .A(n1774), .Y(n1780) );
  INVX1 U21958 ( .A(top_core_KE_n2175), .Y(n2285) );
  INVX1 U21959 ( .A(top_core_KE_n2181), .Y(n2335) );
  INVX1 U21960 ( .A(top_core_KE_n2181), .Y(n2336) );
  INVX1 U21961 ( .A(top_core_EC_n872), .Y(n3558) );
  INVX1 U21962 ( .A(n1753), .Y(n1758) );
  INVX1 U21963 ( .A(n1642), .Y(n1641) );
  INVX1 U21964 ( .A(n4028), .Y(n3988) );
  INVX1 U21965 ( .A(n2366), .Y(n2365) );
  OAI22X1 U21966 ( .A0(n2388), .A1(n6262), .B0(n2407), .B1(n770), .Y(
        top_core_EC_ss_in[42]) );
  OAI22X1 U21967 ( .A0(n2386), .A1(n6230), .B0(n2419), .B1(n776), .Y(
        top_core_EC_ss_in[74]) );
  OAI22X1 U21968 ( .A0(n2391), .A1(n6182), .B0(n2428), .B1(n779), .Y(
        top_core_EC_ss_in[122]) );
  OAI22X1 U21969 ( .A0(n2389), .A1(n6302), .B0(n2402), .B1(n780), .Y(
        top_core_EC_ss_in[2]) );
  OAI22X1 U21970 ( .A0(n2385), .A1(n6222), .B0(n2422), .B1(n782), .Y(
        top_core_EC_ss_in[82]) );
  OAI22X1 U21971 ( .A0(n2392), .A1(n6190), .B0(n2473), .B1(n783), .Y(
        top_core_EC_ss_in[114]) );
  OAI22X1 U21972 ( .A0(n2389), .A1(n6270), .B0(n2404), .B1(n784), .Y(
        top_core_EC_ss_in[34]) );
  OAI22X1 U21973 ( .A0(n2390), .A1(n6278), .B0(n2401), .B1(n785), .Y(
        top_core_EC_ss_in[26]) );
  OAI22X1 U21974 ( .A0(n2386), .A1(n6238), .B0(n2416), .B1(n787), .Y(
        top_core_EC_ss_in[66]) );
  OAI22X1 U21975 ( .A0(n2390), .A1(n6286), .B0(n2438), .B1(n789), .Y(
        top_core_EC_ss_in[18]) );
  OAI22X1 U21976 ( .A0(n2388), .A1(n6206), .B0(n2449), .B1(n792), .Y(
        top_core_EC_ss_in[98]) );
  OAI22X1 U21977 ( .A0(n2388), .A1(n6254), .B0(n2410), .B1(n794), .Y(
        top_core_EC_ss_in[50]) );
  OAI22X1 U21978 ( .A0(n2385), .A1(n6214), .B0(n2425), .B1(n796), .Y(
        top_core_EC_ss_in[90]) );
  OAI22X1 U21979 ( .A0(n2392), .A1(n6198), .B0(n2398), .B1(n821), .Y(
        top_core_EC_ss_in[106]) );
  OAI22X1 U21980 ( .A0(n2387), .A1(n6246), .B0(n2413), .B1(n824), .Y(
        top_core_EC_ss_in[58]) );
  OAI22X1 U21981 ( .A0(n2392), .A1(n6294), .B0(n2399), .B1(n825), .Y(
        top_core_EC_ss_in[10]) );
  OAI22X1 U21982 ( .A0(n2385), .A1(n6219), .B0(n2423), .B1(n801), .Y(
        top_core_EC_ss_in[85]) );
  OAI22X1 U21983 ( .A0(n2385), .A1(n6220), .B0(n2422), .B1(n802), .Y(
        top_core_EC_ss_in[84]) );
  OAI22X1 U21984 ( .A0(n2387), .A1(n6299), .B0(n2413), .B1(n805), .Y(
        top_core_EC_ss_in[5]) );
  OAI22X1 U21985 ( .A0(n2388), .A1(n6300), .B0(n2410), .B1(n806), .Y(
        top_core_EC_ss_in[4]) );
  OAI22X1 U21986 ( .A0(n2391), .A1(n6187), .B0(n2456), .B1(n811), .Y(
        top_core_EC_ss_in[117]) );
  OAI22X1 U21987 ( .A0(n2392), .A1(n6188), .B0(n2406), .B1(n812), .Y(
        top_core_EC_ss_in[116]) );
  OAI22X1 U21988 ( .A0(n2389), .A1(n6267), .B0(n2405), .B1(n813), .Y(
        top_core_EC_ss_in[37]) );
  OAI22X1 U21989 ( .A0(n2389), .A1(n6268), .B0(n2404), .B1(n814), .Y(
        top_core_EC_ss_in[36]) );
  OAI22X1 U21990 ( .A0(n2388), .A1(n6259), .B0(n2408), .B1(n822), .Y(
        top_core_EC_ss_in[45]) );
  OAI22X1 U21991 ( .A0(n2388), .A1(n6260), .B0(n2408), .B1(n823), .Y(
        top_core_EC_ss_in[44]) );
  OAI22X1 U21992 ( .A0(n2391), .A1(n6180), .B0(n2490), .B1(n827), .Y(
        top_core_EC_ss_in[124]) );
  OAI22X1 U21993 ( .A0(n2386), .A1(n6227), .B0(n2420), .B1(n828), .Y(
        top_core_EC_ss_in[77]) );
  OAI22X1 U21994 ( .A0(n2386), .A1(n6228), .B0(n2419), .B1(n829), .Y(
        top_core_EC_ss_in[76]) );
  OAI22X1 U21995 ( .A0(n2391), .A1(n6179), .B0(n2423), .B1(n830), .Y(
        top_core_EC_ss_in[125]) );
  OAI22X1 U21996 ( .A0(n2392), .A1(n6195), .B0(n2399), .B1(n831), .Y(
        top_core_EC_ss_in[109]) );
  OAI22X1 U21997 ( .A0(n2392), .A1(n6196), .B0(n2398), .B1(n832), .Y(
        top_core_EC_ss_in[108]) );
  OAI22X1 U21998 ( .A0(n2387), .A1(n6243), .B0(n2414), .B1(n834), .Y(
        top_core_EC_ss_in[61]) );
  OAI22X1 U21999 ( .A0(n2391), .A1(n6291), .B0(n2441), .B1(n835), .Y(
        top_core_EC_ss_in[13]) );
  OAI22X1 U22000 ( .A0(n2386), .A1(n6236), .B0(n2416), .B1(n838), .Y(
        top_core_EC_ss_in[68]) );
  OAI22X1 U22001 ( .A0(n2386), .A1(n6235), .B0(n2417), .B1(n839), .Y(
        top_core_EC_ss_in[69]) );
  OAI22X1 U22002 ( .A0(n2390), .A1(n6284), .B0(n2527), .B1(n840), .Y(
        top_core_EC_ss_in[20]) );
  OAI22X1 U22003 ( .A0(n2390), .A1(n6283), .B0(n2525), .B1(n841), .Y(
        top_core_EC_ss_in[21]) );
  OAI22X1 U22004 ( .A0(n2393), .A1(n6204), .B0(n2396), .B1(n842), .Y(
        top_core_EC_ss_in[100]) );
  OAI22X1 U22005 ( .A0(n2393), .A1(n6203), .B0(n2396), .B1(n843), .Y(
        top_core_EC_ss_in[101]) );
  OAI22X1 U22006 ( .A0(n2388), .A1(n6252), .B0(n2411), .B1(n844), .Y(
        top_core_EC_ss_in[52]) );
  OAI22X1 U22007 ( .A0(n2387), .A1(n6251), .B0(n2411), .B1(n845), .Y(
        top_core_EC_ss_in[53]) );
  OAI22X1 U22008 ( .A0(n2384), .A1(n6212), .B0(n2425), .B1(n846), .Y(
        top_core_EC_ss_in[92]) );
  OAI22X1 U22009 ( .A0(n2387), .A1(n6244), .B0(n2414), .B1(n848), .Y(
        top_core_EC_ss_in[60]) );
  OAI22X1 U22010 ( .A0(n2389), .A1(n6275), .B0(n2402), .B1(n849), .Y(
        top_core_EC_ss_in[29]) );
  OAI22X1 U22011 ( .A0(n2389), .A1(n6276), .B0(n2401), .B1(n850), .Y(
        top_core_EC_ss_in[28]) );
  OAI22X1 U22012 ( .A0(n2384), .A1(n6211), .B0(n2540), .B1(n851), .Y(
        top_core_EC_ss_in[93]) );
  OAI22X1 U22013 ( .A0(n2393), .A1(n6292), .B0(n2443), .B1(n852), .Y(
        top_core_EC_ss_in[12]) );
  OAI22X1 U22014 ( .A0(n2386), .A1(n6298), .B0(n2417), .B1(n826), .Y(
        top_core_EC_ss_in[6]) );
  OAI22X1 U22015 ( .A0(n2385), .A1(n6218), .B0(n2423), .B1(n833), .Y(
        top_core_EC_ss_in[86]) );
  OAI22X1 U22016 ( .A0(n2391), .A1(n6186), .B0(n2457), .B1(n836), .Y(
        top_core_EC_ss_in[118]) );
  OAI22X1 U22017 ( .A0(n2389), .A1(n6266), .B0(n2405), .B1(n837), .Y(
        top_core_EC_ss_in[38]) );
  OAI22X1 U22018 ( .A0(n2388), .A1(n6258), .B0(n2408), .B1(n847), .Y(
        top_core_EC_ss_in[46]) );
  OAI22X1 U22019 ( .A0(n2386), .A1(n6226), .B0(n2420), .B1(n853), .Y(
        top_core_EC_ss_in[78]) );
  OAI22X1 U22020 ( .A0(n2392), .A1(n6194), .B0(n2399), .B1(n854), .Y(
        top_core_EC_ss_in[110]) );
  OAI22X1 U22021 ( .A0(n2387), .A1(n6242), .B0(n2414), .B1(n857), .Y(
        top_core_EC_ss_in[62]) );
  OAI22X1 U22022 ( .A0(n2391), .A1(n6178), .B0(n2425), .B1(n858), .Y(
        top_core_EC_ss_in[126]) );
  OAI22X1 U22023 ( .A0(n2391), .A1(n6290), .B0(n2450), .B1(n859), .Y(
        top_core_EC_ss_in[14]) );
  OAI22X1 U22024 ( .A0(n2386), .A1(n6234), .B0(n2417), .B1(n862), .Y(
        top_core_EC_ss_in[70]) );
  OAI22X1 U22025 ( .A0(n2390), .A1(n6282), .B0(n2527), .B1(n863), .Y(
        top_core_EC_ss_in[22]) );
  OAI22X1 U22026 ( .A0(n2393), .A1(n6202), .B0(n2396), .B1(n864), .Y(
        top_core_EC_ss_in[102]) );
  OAI22X1 U22027 ( .A0(n2387), .A1(n6250), .B0(n2411), .B1(n865), .Y(
        top_core_EC_ss_in[54]) );
  OAI22X1 U22028 ( .A0(n2384), .A1(n6210), .B0(n2421), .B1(n866), .Y(
        top_core_EC_ss_in[94]) );
  OAI22X1 U22029 ( .A0(n2389), .A1(n6274), .B0(n2402), .B1(n867), .Y(
        top_core_EC_ss_in[30]) );
  AND2X2 U22030 ( .A(top_core_KE_n2692), .B(top_core_KE_round_ctr_reg_0_), .Y(
        n767) );
  INVX1 U22031 ( .A(top_core_KE_n918), .Y(n2221) );
  NOR2BX1 U22032 ( .AN(top_core_KE_n894), .B(top_core_KE_n2701), .Y(
        top_core_KE_n918) );
  INVX1 U22033 ( .A(top_core_EC_ss_in[0]), .Y(n3507) );
  OAI22X1 U22034 ( .A0(n2393), .A1(n6304), .B0(n2395), .B1(n769), .Y(
        top_core_EC_ss_in[0]) );
  INVX1 U22035 ( .A(top_core_EC_ss_in[1]), .Y(n3492) );
  OAI22X1 U22036 ( .A0(n2390), .A1(n6303), .B0(n2480), .B1(n771), .Y(
        top_core_EC_ss_in[1]) );
  INVX1 U22037 ( .A(top_core_EC_ss_in[81]), .Y(n2891) );
  OAI22X1 U22038 ( .A0(n2385), .A1(n6223), .B0(n2421), .B1(n772), .Y(
        top_core_EC_ss_in[81]) );
  INVX1 U22039 ( .A(top_core_EC_ss_in[113]), .Y(n2649) );
  OAI22X1 U22040 ( .A0(n2392), .A1(n6191), .B0(n2531), .B1(n773), .Y(
        top_core_EC_ss_in[113]) );
  INVX1 U22041 ( .A(top_core_EC_ss_in[33]), .Y(n3251) );
  OAI22X1 U22042 ( .A0(n2389), .A1(n6271), .B0(n2403), .B1(n774), .Y(
        top_core_EC_ss_in[33]) );
  OAI22X1 U22043 ( .A0(n2385), .A1(n6224), .B0(n2421), .B1(n775), .Y(
        top_core_EC_ss_in[80]) );
  INVX1 U22044 ( .A(top_core_EC_ss_in[112]), .Y(n2664) );
  OAI22X1 U22045 ( .A0(n2392), .A1(n6192), .B0(n2528), .B1(n777), .Y(
        top_core_EC_ss_in[112]) );
  OAI22X1 U22046 ( .A0(n2389), .A1(n6272), .B0(n2403), .B1(n778), .Y(
        top_core_EC_ss_in[32]) );
  INVX1 U22047 ( .A(top_core_EC_ss_in[57]), .Y(n3071) );
  OAI22X1 U22048 ( .A0(n2387), .A1(n6247), .B0(n2412), .B1(n781), .Y(
        top_core_EC_ss_in[57]) );
  INVX1 U22049 ( .A(top_core_EC_ss_in[9]), .Y(n3431) );
  OAI22X1 U22050 ( .A0(n2393), .A1(n6295), .B0(n768), .B1(n2449), .Y(
        top_core_EC_ss_in[9]) );
  INVX1 U22051 ( .A(top_core_EC_ss_in[89]), .Y(n2831) );
  OAI22X1 U22052 ( .A0(n2385), .A1(n6215), .B0(n2424), .B1(n786), .Y(
        top_core_EC_ss_in[89]) );
  INVX1 U22053 ( .A(top_core_EC_ss_in[65]), .Y(n3013) );
  OAI22X1 U22054 ( .A0(n2387), .A1(n6239), .B0(n2415), .B1(n788), .Y(
        top_core_EC_ss_in[65]) );
  OAI22X1 U22055 ( .A0(n2390), .A1(n6287), .B0(n2435), .B1(n790), .Y(
        top_core_EC_ss_in[17]) );
  OAI22X1 U22056 ( .A0(n2391), .A1(n6183), .B0(n2488), .B1(n791), .Y(
        top_core_EC_ss_in[121]) );
  OAI22X1 U22057 ( .A0(n2384), .A1(n6207), .B0(n2524), .B1(n793), .Y(
        top_core_EC_ss_in[97]) );
  OAI22X1 U22058 ( .A0(n2388), .A1(n6255), .B0(n2409), .B1(n795), .Y(
        top_core_EC_ss_in[49]) );
  INVX1 U22059 ( .A(top_core_EC_ss_in[25]), .Y(n3312) );
  OAI22X1 U22060 ( .A0(n2390), .A1(n6279), .B0(n2400), .B1(n797), .Y(
        top_core_EC_ss_in[25]) );
  OAI22X1 U22061 ( .A0(n2392), .A1(n6200), .B0(n2397), .B1(n798), .Y(
        top_core_EC_ss_in[104]) );
  OAI22X1 U22062 ( .A0(n2388), .A1(n6264), .B0(n2406), .B1(n799), .Y(
        top_core_EC_ss_in[40]) );
  OAI22X1 U22063 ( .A0(n2392), .A1(n6199), .B0(n2397), .B1(n800), .Y(
        top_core_EC_ss_in[105]) );
  INVX1 U22064 ( .A(top_core_EC_ss_in[56]), .Y(n3086) );
  OAI22X1 U22065 ( .A0(n2387), .A1(n6248), .B0(n2412), .B1(n803), .Y(
        top_core_EC_ss_in[56]) );
  OAI22X1 U22066 ( .A0(n2388), .A1(n6263), .B0(n2407), .B1(n804), .Y(
        top_core_EC_ss_in[41]) );
  INVX1 U22067 ( .A(top_core_EC_ss_in[120]), .Y(n2603) );
  OAI22X1 U22068 ( .A0(n2391), .A1(n6184), .B0(n2492), .B1(n807), .Y(
        top_core_EC_ss_in[120]) );
  OAI22X1 U22069 ( .A0(n2385), .A1(n6296), .B0(n2424), .B1(n808), .Y(
        top_core_EC_ss_in[8]) );
  OAI22X1 U22070 ( .A0(n2386), .A1(n6232), .B0(n2418), .B1(n809), .Y(
        top_core_EC_ss_in[72]) );
  INVX1 U22071 ( .A(top_core_EC_ss_in[73]), .Y(n2952) );
  OAI22X1 U22072 ( .A0(n2386), .A1(n6231), .B0(n2418), .B1(n810), .Y(
        top_core_EC_ss_in[73]) );
  INVX1 U22073 ( .A(top_core_EC_ss_in[24]), .Y(n3327) );
  OAI22X1 U22074 ( .A0(n2390), .A1(n6280), .B0(n2400), .B1(n815), .Y(
        top_core_EC_ss_in[24]) );
  INVX1 U22075 ( .A(top_core_EC_ss_in[64]), .Y(n3025) );
  OAI22X1 U22076 ( .A0(n2387), .A1(n6240), .B0(n2415), .B1(n816), .Y(
        top_core_EC_ss_in[64]) );
  INVX1 U22077 ( .A(top_core_EC_ss_in[16]), .Y(n3385) );
  OAI22X1 U22078 ( .A0(n2390), .A1(n6288), .B0(n2429), .B1(n817), .Y(
        top_core_EC_ss_in[16]) );
  INVX1 U22079 ( .A(top_core_EC_ss_in[96]), .Y(n2785) );
  OAI22X1 U22080 ( .A0(n2384), .A1(n6208), .B0(n2541), .B1(n818), .Y(
        top_core_EC_ss_in[96]) );
  INVX1 U22081 ( .A(top_core_EC_ss_in[48]), .Y(n3144) );
  OAI22X1 U22082 ( .A0(n2388), .A1(n6256), .B0(n2409), .B1(n819), .Y(
        top_core_EC_ss_in[48]) );
  OAI22X1 U22083 ( .A0(n2385), .A1(n6216), .B0(n2424), .B1(n820), .Y(
        top_core_EC_ss_in[88]) );
  OAI21XL U22084 ( .A0(n2393), .A1(top_core_EC_n946), .B0(n2), .Y(
        top_core_EC_n948) );
  INVX1 U22085 ( .A(n_WR), .Y(n4192) );
  OAI2BB2X1 U22086 ( .B0(n1578), .B1(top_core_io_n5), .A0N(top_core_io_n5), 
        .A1N(top_core_io_NK_0_), .Y(top_core_io_n664) );
  OAI2BB2X1 U22087 ( .B0(top_core_io_n661), .B1(top_core_io_n657), .A0N(
        top_core_io_N81), .A1N(top_core_io_n656), .Y(top_core_io_N90) );
  NOR2X2 U22088 ( .A(n_ADDR[6]), .B(n_WR), .Y(top_core_io_n656) );
  OAI2BB2X1 U22089 ( .B0(top_core_io_n1), .B1(n4260), .A0N(top_core_io_n1), 
        .A1N(n_DIN[0]), .Y(top_core_io_n663) );
  AND3X2 U22090 ( .A(n_ADDR[6]), .B(n4127), .C(n_WR), .Y(top_core_io_n1) );
  OAI21XL U22091 ( .A0(top_core_io_CORE_FULL), .A1(n4144), .B0(
        top_core_io_n655), .Y(top_core_io_n1183) );
  OAI2BB1X1 U22092 ( .A0N(top_core_t_ready), .A1N(n3704), .B0(
        top_core_io_inter_ok), .Y(top_core_io_n655) );
  OAI2BB1X1 U22093 ( .A0N(n_OK), .A1N(n4144), .B0(n3673), .Y(top_core_io_n1182) );
  INVX1 U22094 ( .A(n_START), .Y(n4144) );
  XOR2X1 U22095 ( .A(top_core_clk_slow), .B(top_core_io_div_16_n1), .Y(
        top_core_io_div_16_n3) );
  NOR2BX1 U22096 ( .AN(top_core_io_div_16_c_2_), .B(top_core_io_div_16_n2), 
        .Y(top_core_io_div_16_n1) );
  NAND2BX1 U22097 ( .AN(top_core_io_div_16_n5), .B(top_core_io_div_16_c_1_), 
        .Y(top_core_io_div_16_n2) );
  INVX1 U22098 ( .A(top_core_io_n460), .Y(n4622) );
  AOI22X1 U22099 ( .A0(top_core_Ciphertext[31]), .A1(n3651), .B0(
        top_core_io_Data_reg_19__7_), .B1(n3678), .Y(top_core_io_n460) );
  INVX1 U22100 ( .A(top_core_io_n459), .Y(n4621) );
  AOI22X1 U22101 ( .A0(top_core_Ciphertext[30]), .A1(n3679), .B0(
        top_core_io_Data_reg_19__6_), .B1(n3644), .Y(top_core_io_n459) );
  INVX1 U22102 ( .A(top_core_io_n458), .Y(n4620) );
  AOI22X1 U22103 ( .A0(top_core_Ciphertext[29]), .A1(n3685), .B0(
        top_core_io_Data_reg_19__5_), .B1(n3674), .Y(top_core_io_n458) );
  INVX1 U22104 ( .A(top_core_io_n457), .Y(n4619) );
  AOI22X1 U22105 ( .A0(top_core_Ciphertext[28]), .A1(n3680), .B0(
        top_core_io_Data_reg_19__4_), .B1(n3675), .Y(top_core_io_n457) );
  INVX1 U22106 ( .A(top_core_io_n456), .Y(n4618) );
  AOI22X1 U22107 ( .A0(top_core_Ciphertext[27]), .A1(n3681), .B0(
        top_core_io_Data_reg_19__3_), .B1(n3669), .Y(top_core_io_n456) );
  INVX1 U22108 ( .A(top_core_io_n455), .Y(n4617) );
  AOI22X1 U22109 ( .A0(top_core_Ciphertext[26]), .A1(n3682), .B0(
        top_core_io_Data_reg_19__2_), .B1(n3668), .Y(top_core_io_n455) );
  INVX1 U22110 ( .A(top_core_io_n454), .Y(n4616) );
  AOI22X1 U22111 ( .A0(top_core_Ciphertext[25]), .A1(n3645), .B0(
        top_core_io_Data_reg_19__1_), .B1(n3655), .Y(top_core_io_n454) );
  INVX1 U22112 ( .A(top_core_io_n453), .Y(n4615) );
  AOI22X1 U22113 ( .A0(top_core_Ciphertext[24]), .A1(top_core_c_ready), .B0(
        top_core_io_Data_reg_19__0_), .B1(n3673), .Y(top_core_io_n453) );
  INVX1 U22114 ( .A(top_core_io_n428), .Y(n4590) );
  AOI22X1 U22115 ( .A0(top_core_Ciphertext[63]), .A1(n3646), .B0(
        top_core_io_Data_reg_23__7_), .B1(n3664), .Y(top_core_io_n428) );
  INVX1 U22116 ( .A(top_core_io_n427), .Y(n4589) );
  AOI22X1 U22117 ( .A0(top_core_Ciphertext[62]), .A1(n3646), .B0(
        top_core_io_Data_reg_23__6_), .B1(n3664), .Y(top_core_io_n427) );
  INVX1 U22118 ( .A(top_core_io_n426), .Y(n4588) );
  AOI22X1 U22119 ( .A0(top_core_Ciphertext[61]), .A1(n3646), .B0(
        top_core_io_Data_reg_23__5_), .B1(n3663), .Y(top_core_io_n426) );
  INVX1 U22120 ( .A(top_core_io_n425), .Y(n4587) );
  AOI22X1 U22121 ( .A0(top_core_Ciphertext[60]), .A1(n3646), .B0(
        top_core_io_Data_reg_23__4_), .B1(n3663), .Y(top_core_io_n425) );
  INVX1 U22122 ( .A(top_core_io_n424), .Y(n4586) );
  AOI22X1 U22123 ( .A0(top_core_Ciphertext[59]), .A1(n3647), .B0(
        top_core_io_Data_reg_23__3_), .B1(n3665), .Y(top_core_io_n424) );
  INVX1 U22124 ( .A(top_core_io_n423), .Y(n4585) );
  AOI22X1 U22125 ( .A0(top_core_Ciphertext[58]), .A1(n3647), .B0(
        top_core_io_Data_reg_23__2_), .B1(n3664), .Y(top_core_io_n423) );
  INVX1 U22126 ( .A(top_core_io_n422), .Y(n4584) );
  AOI22X1 U22127 ( .A0(top_core_Ciphertext[57]), .A1(n3647), .B0(
        top_core_io_Data_reg_23__1_), .B1(n3677), .Y(top_core_io_n422) );
  INVX1 U22128 ( .A(top_core_io_n421), .Y(n4583) );
  AOI22X1 U22129 ( .A0(top_core_Ciphertext[56]), .A1(n3647), .B0(
        top_core_io_Data_reg_23__0_), .B1(n3678), .Y(top_core_io_n421) );
  INVX1 U22130 ( .A(top_core_io_n396), .Y(n4558) );
  AOI22X1 U22131 ( .A0(top_core_Ciphertext[95]), .A1(n3649), .B0(
        top_core_io_Data_reg_27__7_), .B1(n3667), .Y(top_core_io_n396) );
  INVX1 U22132 ( .A(top_core_io_n395), .Y(n4557) );
  AOI22X1 U22133 ( .A0(top_core_Ciphertext[94]), .A1(n3649), .B0(
        top_core_io_Data_reg_27__6_), .B1(n3644), .Y(top_core_io_n395) );
  INVX1 U22134 ( .A(top_core_io_n394), .Y(n4556) );
  AOI22X1 U22135 ( .A0(top_core_Ciphertext[93]), .A1(n3649), .B0(
        top_core_io_Data_reg_27__5_), .B1(n3658), .Y(top_core_io_n394) );
  INVX1 U22136 ( .A(top_core_io_n393), .Y(n4555) );
  AOI22X1 U22137 ( .A0(top_core_Ciphertext[92]), .A1(n3649), .B0(
        top_core_io_Data_reg_27__4_), .B1(n3657), .Y(top_core_io_n393) );
  INVX1 U22138 ( .A(top_core_io_n392), .Y(n4554) );
  AOI22X1 U22139 ( .A0(top_core_Ciphertext[91]), .A1(n3649), .B0(
        top_core_io_Data_reg_27__3_), .B1(n3661), .Y(top_core_io_n392) );
  INVX1 U22140 ( .A(top_core_io_n391), .Y(n4553) );
  AOI22X1 U22141 ( .A0(top_core_Ciphertext[90]), .A1(n3649), .B0(
        top_core_io_Data_reg_27__2_), .B1(n3660), .Y(top_core_io_n391) );
  INVX1 U22142 ( .A(top_core_io_n390), .Y(n4552) );
  AOI22X1 U22143 ( .A0(top_core_Ciphertext[89]), .A1(n3649), .B0(
        top_core_io_Data_reg_27__1_), .B1(n3663), .Y(top_core_io_n390) );
  INVX1 U22144 ( .A(top_core_io_n389), .Y(n4551) );
  AOI22X1 U22145 ( .A0(top_core_Ciphertext[88]), .A1(n3649), .B0(
        top_core_io_Data_reg_27__0_), .B1(n3676), .Y(top_core_io_n389) );
  INVX1 U22146 ( .A(top_core_io_n364), .Y(n4526) );
  AOI22X1 U22147 ( .A0(top_core_Ciphertext[127]), .A1(n3651), .B0(
        top_core_io_Data_reg_31__7_), .B1(n3673), .Y(top_core_io_n364) );
  INVX1 U22148 ( .A(top_core_io_n363), .Y(n4525) );
  AOI22X1 U22149 ( .A0(top_core_Ciphertext[126]), .A1(n3651), .B0(
        top_core_io_Data_reg_31__6_), .B1(n3670), .Y(top_core_io_n363) );
  INVX1 U22150 ( .A(top_core_io_n362), .Y(n4524) );
  AOI22X1 U22151 ( .A0(top_core_Ciphertext[125]), .A1(n3651), .B0(
        top_core_io_Data_reg_31__5_), .B1(n3677), .Y(top_core_io_n362) );
  INVX1 U22152 ( .A(top_core_io_n361), .Y(n4523) );
  AOI22X1 U22153 ( .A0(top_core_Ciphertext[124]), .A1(n3651), .B0(
        top_core_io_Data_reg_31__4_), .B1(n3656), .Y(top_core_io_n361) );
  INVX1 U22154 ( .A(top_core_io_n360), .Y(n4522) );
  AOI22X1 U22155 ( .A0(top_core_Ciphertext[123]), .A1(n3651), .B0(
        top_core_io_Data_reg_31__3_), .B1(n3662), .Y(top_core_io_n360) );
  INVX1 U22156 ( .A(top_core_io_n359), .Y(n4521) );
  AOI22X1 U22157 ( .A0(top_core_Ciphertext[122]), .A1(n3651), .B0(
        top_core_io_Data_reg_31__2_), .B1(n3661), .Y(top_core_io_n359) );
  INVX1 U22158 ( .A(top_core_io_n358), .Y(n4520) );
  AOI22X1 U22159 ( .A0(top_core_Ciphertext[121]), .A1(n3651), .B0(
        top_core_io_Data_reg_31__1_), .B1(n3671), .Y(top_core_io_n358) );
  INVX1 U22160 ( .A(top_core_io_n356), .Y(n4519) );
  AOI22X1 U22161 ( .A0(n3651), .A1(top_core_Ciphertext[120]), .B0(
        top_core_io_Data_reg_31__0_), .B1(n3652), .Y(top_core_io_n356) );
  INVX1 U22162 ( .A(top_core_io_NK_1_), .Y(n4261) );
  INVX1 U22163 ( .A(top_core_io_NK_2_), .Y(n4262) );
  INVX1 U22164 ( .A(top_core_io_CipherKey_w_247_), .Y(n4278) );
  INVX1 U22165 ( .A(top_core_io_CipherKey_w_246_), .Y(n4277) );
  INVX1 U22166 ( .A(top_core_io_CipherKey_w_245_), .Y(n4276) );
  INVX1 U22167 ( .A(top_core_io_CipherKey_w_244_), .Y(n4275) );
  INVX1 U22168 ( .A(top_core_io_CipherKey_w_243_), .Y(n4274) );
  INVX1 U22169 ( .A(top_core_io_CipherKey_w_242_), .Y(n4273) );
  INVX1 U22170 ( .A(top_core_io_CipherKey_w_241_), .Y(n4272) );
  INVX1 U22171 ( .A(top_core_io_CipherKey_w_240_), .Y(n4271) );
  INVX1 U22172 ( .A(top_core_io_CipherKey_w_215_), .Y(n4310) );
  INVX1 U22173 ( .A(top_core_io_CipherKey_w_214_), .Y(n4309) );
  INVX1 U22174 ( .A(top_core_io_CipherKey_w_213_), .Y(n4308) );
  INVX1 U22175 ( .A(top_core_io_CipherKey_w_212_), .Y(n4307) );
  INVX1 U22176 ( .A(top_core_io_CipherKey_w_211_), .Y(n4306) );
  INVX1 U22177 ( .A(top_core_io_CipherKey_w_210_), .Y(n4305) );
  INVX1 U22178 ( .A(top_core_io_CipherKey_w_209_), .Y(n4304) );
  INVX1 U22179 ( .A(top_core_io_CipherKey_w_208_), .Y(n4303) );
  INVX1 U22180 ( .A(top_core_io_CipherKey_w_119_), .Y(n4406) );
  INVX1 U22181 ( .A(top_core_io_CipherKey_w_118_), .Y(n4405) );
  INVX1 U22182 ( .A(top_core_io_CipherKey_w_117_), .Y(n4404) );
  INVX1 U22183 ( .A(top_core_io_CipherKey_w_116_), .Y(n4403) );
  INVX1 U22184 ( .A(top_core_io_CipherKey_w_115_), .Y(n4402) );
  INVX1 U22185 ( .A(top_core_io_CipherKey_w_114_), .Y(n4401) );
  INVX1 U22186 ( .A(top_core_io_CipherKey_w_113_), .Y(n4400) );
  INVX1 U22187 ( .A(top_core_io_CipherKey_w_112_), .Y(n4399) );
  INVX1 U22188 ( .A(top_core_io_CipherKey_w_87_), .Y(n4438) );
  INVX1 U22189 ( .A(top_core_io_CipherKey_w_86_), .Y(n4437) );
  INVX1 U22190 ( .A(top_core_io_CipherKey_w_85_), .Y(n4436) );
  INVX1 U22191 ( .A(top_core_io_CipherKey_w_84_), .Y(n4435) );
  INVX1 U22192 ( .A(top_core_io_CipherKey_w_83_), .Y(n4434) );
  INVX1 U22193 ( .A(top_core_io_CipherKey_w_82_), .Y(n4433) );
  INVX1 U22194 ( .A(top_core_io_CipherKey_w_81_), .Y(n4432) );
  INVX1 U22195 ( .A(top_core_io_CipherKey_w_80_), .Y(n4431) );
  INVX1 U22196 ( .A(top_core_io_Plain_text_w_119_), .Y(n4662) );
  INVX1 U22197 ( .A(top_core_io_Plain_text_w_118_), .Y(n4661) );
  INVX1 U22198 ( .A(top_core_io_Plain_text_w_117_), .Y(n4660) );
  INVX1 U22199 ( .A(top_core_io_Plain_text_w_116_), .Y(n4659) );
  INVX1 U22200 ( .A(top_core_io_Plain_text_w_115_), .Y(n4658) );
  INVX1 U22201 ( .A(top_core_io_Plain_text_w_114_), .Y(n4657) );
  INVX1 U22202 ( .A(top_core_io_Plain_text_w_113_), .Y(n4656) );
  INVX1 U22203 ( .A(top_core_io_Plain_text_w_112_), .Y(n4655) );
  INVX1 U22204 ( .A(top_core_io_Plain_text_w_87_), .Y(n4694) );
  INVX1 U22205 ( .A(top_core_io_Plain_text_w_86_), .Y(n4693) );
  INVX1 U22206 ( .A(top_core_io_Plain_text_w_85_), .Y(n4692) );
  INVX1 U22207 ( .A(top_core_io_Plain_text_w_84_), .Y(n4691) );
  INVX1 U22208 ( .A(top_core_io_Plain_text_w_83_), .Y(n4690) );
  INVX1 U22209 ( .A(top_core_io_Plain_text_w_82_), .Y(n4689) );
  INVX1 U22210 ( .A(top_core_io_Plain_text_w_81_), .Y(n4688) );
  INVX1 U22211 ( .A(top_core_io_Plain_text_w_80_), .Y(n4687) );
  INVX1 U22212 ( .A(top_core_io_CipherKey_w_231_), .Y(n4294) );
  INVX1 U22213 ( .A(top_core_io_CipherKey_w_230_), .Y(n4293) );
  INVX1 U22214 ( .A(top_core_io_CipherKey_w_229_), .Y(n4292) );
  INVX1 U22215 ( .A(top_core_io_CipherKey_w_228_), .Y(n4291) );
  INVX1 U22216 ( .A(top_core_io_CipherKey_w_227_), .Y(n4290) );
  INVX1 U22217 ( .A(top_core_io_CipherKey_w_226_), .Y(n4289) );
  INVX1 U22218 ( .A(top_core_io_CipherKey_w_225_), .Y(n4288) );
  INVX1 U22219 ( .A(top_core_io_CipherKey_w_224_), .Y(n4287) );
  INVX1 U22220 ( .A(top_core_io_CipherKey_w_103_), .Y(n4422) );
  INVX1 U22221 ( .A(top_core_io_CipherKey_w_102_), .Y(n4421) );
  INVX1 U22222 ( .A(top_core_io_CipherKey_w_101_), .Y(n4420) );
  INVX1 U22223 ( .A(top_core_io_CipherKey_w_100_), .Y(n4419) );
  INVX1 U22224 ( .A(top_core_io_CipherKey_w_99_), .Y(n4418) );
  INVX1 U22225 ( .A(top_core_io_CipherKey_w_98_), .Y(n4417) );
  INVX1 U22226 ( .A(top_core_io_CipherKey_w_97_), .Y(n4416) );
  INVX1 U22227 ( .A(top_core_io_CipherKey_w_96_), .Y(n4415) );
  INVX1 U22228 ( .A(top_core_io_Plain_text_w_103_), .Y(n4678) );
  INVX1 U22229 ( .A(top_core_io_Plain_text_w_102_), .Y(n4677) );
  INVX1 U22230 ( .A(top_core_io_Plain_text_w_101_), .Y(n4676) );
  INVX1 U22231 ( .A(top_core_io_Plain_text_w_100_), .Y(n4675) );
  INVX1 U22232 ( .A(top_core_io_Plain_text_w_99_), .Y(n4674) );
  INVX1 U22233 ( .A(top_core_io_Plain_text_w_98_), .Y(n4673) );
  INVX1 U22234 ( .A(top_core_io_Plain_text_w_97_), .Y(n4672) );
  INVX1 U22235 ( .A(top_core_io_Plain_text_w_96_), .Y(n4671) );
  INVX1 U22236 ( .A(top_core_io_CipherKey_w_255_), .Y(n4270) );
  INVX1 U22237 ( .A(top_core_io_CipherKey_w_254_), .Y(n4269) );
  INVX1 U22238 ( .A(top_core_io_CipherKey_w_253_), .Y(n4268) );
  INVX1 U22239 ( .A(top_core_io_CipherKey_w_252_), .Y(n4267) );
  INVX1 U22240 ( .A(top_core_io_CipherKey_w_251_), .Y(n4266) );
  INVX1 U22241 ( .A(top_core_io_CipherKey_w_250_), .Y(n4265) );
  INVX1 U22242 ( .A(top_core_io_CipherKey_w_249_), .Y(n4264) );
  INVX1 U22243 ( .A(top_core_io_CipherKey_w_248_), .Y(n4263) );
  INVX1 U22244 ( .A(top_core_io_CipherKey_w_223_), .Y(n4302) );
  INVX1 U22245 ( .A(top_core_io_CipherKey_w_222_), .Y(n4301) );
  INVX1 U22246 ( .A(top_core_io_CipherKey_w_221_), .Y(n4300) );
  INVX1 U22247 ( .A(top_core_io_CipherKey_w_220_), .Y(n4299) );
  INVX1 U22248 ( .A(top_core_io_CipherKey_w_219_), .Y(n4298) );
  INVX1 U22249 ( .A(top_core_io_CipherKey_w_218_), .Y(n4297) );
  INVX1 U22250 ( .A(top_core_io_CipherKey_w_217_), .Y(n4296) );
  INVX1 U22251 ( .A(top_core_io_CipherKey_w_216_), .Y(n4295) );
  INVX1 U22252 ( .A(top_core_io_CipherKey_w_127_), .Y(n4398) );
  INVX1 U22253 ( .A(top_core_io_CipherKey_w_126_), .Y(n4397) );
  INVX1 U22254 ( .A(top_core_io_CipherKey_w_125_), .Y(n4396) );
  INVX1 U22255 ( .A(top_core_io_CipherKey_w_124_), .Y(n4395) );
  INVX1 U22256 ( .A(top_core_io_CipherKey_w_123_), .Y(n4394) );
  INVX1 U22257 ( .A(top_core_io_CipherKey_w_122_), .Y(n4393) );
  INVX1 U22258 ( .A(top_core_io_CipherKey_w_121_), .Y(n4392) );
  INVX1 U22259 ( .A(top_core_io_CipherKey_w_120_), .Y(n4391) );
  INVX1 U22260 ( .A(top_core_io_CipherKey_w_95_), .Y(n4430) );
  INVX1 U22261 ( .A(top_core_io_CipherKey_w_94_), .Y(n4429) );
  INVX1 U22262 ( .A(top_core_io_CipherKey_w_93_), .Y(n4428) );
  INVX1 U22263 ( .A(top_core_io_CipherKey_w_92_), .Y(n4427) );
  INVX1 U22264 ( .A(top_core_io_CipherKey_w_91_), .Y(n4426) );
  INVX1 U22265 ( .A(top_core_io_CipherKey_w_90_), .Y(n4425) );
  INVX1 U22266 ( .A(top_core_io_CipherKey_w_89_), .Y(n4424) );
  INVX1 U22267 ( .A(top_core_io_CipherKey_w_88_), .Y(n4423) );
  INVX1 U22268 ( .A(top_core_io_Plain_text_w_127_), .Y(n4654) );
  INVX1 U22269 ( .A(top_core_io_Plain_text_w_126_), .Y(n4653) );
  INVX1 U22270 ( .A(top_core_io_Plain_text_w_125_), .Y(n4652) );
  INVX1 U22271 ( .A(top_core_io_Plain_text_w_124_), .Y(n4651) );
  INVX1 U22272 ( .A(top_core_io_Plain_text_w_123_), .Y(n4650) );
  INVX1 U22273 ( .A(top_core_io_Plain_text_w_122_), .Y(n4649) );
  INVX1 U22274 ( .A(top_core_io_Plain_text_w_121_), .Y(n4648) );
  INVX1 U22275 ( .A(top_core_io_Plain_text_w_120_), .Y(n4647) );
  INVX1 U22276 ( .A(top_core_io_Plain_text_w_95_), .Y(n4686) );
  INVX1 U22277 ( .A(top_core_io_Plain_text_w_94_), .Y(n4685) );
  INVX1 U22278 ( .A(top_core_io_Plain_text_w_93_), .Y(n4684) );
  INVX1 U22279 ( .A(top_core_io_Plain_text_w_92_), .Y(n4683) );
  INVX1 U22280 ( .A(top_core_io_Plain_text_w_91_), .Y(n4682) );
  INVX1 U22281 ( .A(top_core_io_Plain_text_w_90_), .Y(n4681) );
  INVX1 U22282 ( .A(top_core_io_Plain_text_w_89_), .Y(n4680) );
  INVX1 U22283 ( .A(top_core_io_Plain_text_w_88_), .Y(n4679) );
  INVX1 U22284 ( .A(top_core_io_CipherKey_w_239_), .Y(n4286) );
  INVX1 U22285 ( .A(top_core_io_CipherKey_w_238_), .Y(n4285) );
  INVX1 U22286 ( .A(top_core_io_CipherKey_w_237_), .Y(n4284) );
  INVX1 U22287 ( .A(top_core_io_CipherKey_w_236_), .Y(n4283) );
  INVX1 U22288 ( .A(top_core_io_CipherKey_w_235_), .Y(n4282) );
  INVX1 U22289 ( .A(top_core_io_CipherKey_w_234_), .Y(n4281) );
  INVX1 U22290 ( .A(top_core_io_CipherKey_w_233_), .Y(n4280) );
  INVX1 U22291 ( .A(top_core_io_CipherKey_w_232_), .Y(n4279) );
  INVX1 U22292 ( .A(top_core_io_CipherKey_w_207_), .Y(n4318) );
  INVX1 U22293 ( .A(top_core_io_CipherKey_w_206_), .Y(n4317) );
  INVX1 U22294 ( .A(top_core_io_CipherKey_w_205_), .Y(n4316) );
  INVX1 U22295 ( .A(top_core_io_CipherKey_w_204_), .Y(n4315) );
  INVX1 U22296 ( .A(top_core_io_CipherKey_w_203_), .Y(n4314) );
  INVX1 U22297 ( .A(top_core_io_CipherKey_w_202_), .Y(n4313) );
  INVX1 U22298 ( .A(top_core_io_CipherKey_w_201_), .Y(n4312) );
  INVX1 U22299 ( .A(top_core_io_CipherKey_w_200_), .Y(n4311) );
  INVX1 U22300 ( .A(top_core_io_CipherKey_w_111_), .Y(n4414) );
  INVX1 U22301 ( .A(top_core_io_CipherKey_w_110_), .Y(n4413) );
  INVX1 U22302 ( .A(top_core_io_CipherKey_w_109_), .Y(n4412) );
  INVX1 U22303 ( .A(top_core_io_CipherKey_w_108_), .Y(n4411) );
  INVX1 U22304 ( .A(top_core_io_CipherKey_w_107_), .Y(n4410) );
  INVX1 U22305 ( .A(top_core_io_CipherKey_w_106_), .Y(n4409) );
  INVX1 U22306 ( .A(top_core_io_CipherKey_w_105_), .Y(n4408) );
  INVX1 U22307 ( .A(top_core_io_CipherKey_w_104_), .Y(n4407) );
  INVX1 U22308 ( .A(top_core_io_CipherKey_w_79_), .Y(n4446) );
  INVX1 U22309 ( .A(top_core_io_CipherKey_w_78_), .Y(n4445) );
  INVX1 U22310 ( .A(top_core_io_CipherKey_w_77_), .Y(n4444) );
  INVX1 U22311 ( .A(top_core_io_CipherKey_w_76_), .Y(n4443) );
  INVX1 U22312 ( .A(top_core_io_CipherKey_w_75_), .Y(n4442) );
  INVX1 U22313 ( .A(top_core_io_CipherKey_w_74_), .Y(n4441) );
  INVX1 U22314 ( .A(top_core_io_CipherKey_w_73_), .Y(n4440) );
  INVX1 U22315 ( .A(top_core_io_CipherKey_w_72_), .Y(n4439) );
  INVX1 U22316 ( .A(top_core_io_Plain_text_w_111_), .Y(n4670) );
  INVX1 U22317 ( .A(top_core_io_Plain_text_w_110_), .Y(n4669) );
  INVX1 U22318 ( .A(top_core_io_Plain_text_w_109_), .Y(n4668) );
  INVX1 U22319 ( .A(top_core_io_Plain_text_w_108_), .Y(n4667) );
  INVX1 U22320 ( .A(top_core_io_Plain_text_w_107_), .Y(n4666) );
  INVX1 U22321 ( .A(top_core_io_Plain_text_w_106_), .Y(n4665) );
  INVX1 U22322 ( .A(top_core_io_Plain_text_w_105_), .Y(n4664) );
  INVX1 U22323 ( .A(top_core_io_Plain_text_w_104_), .Y(n4663) );
  INVX1 U22324 ( .A(top_core_io_Plain_text_w_79_), .Y(n4702) );
  INVX1 U22325 ( .A(top_core_io_Plain_text_w_78_), .Y(n4701) );
  INVX1 U22326 ( .A(top_core_io_Plain_text_w_77_), .Y(n4700) );
  INVX1 U22327 ( .A(top_core_io_Plain_text_w_76_), .Y(n4699) );
  INVX1 U22328 ( .A(top_core_io_Plain_text_w_75_), .Y(n4698) );
  INVX1 U22329 ( .A(top_core_io_Plain_text_w_74_), .Y(n4697) );
  INVX1 U22330 ( .A(top_core_io_Plain_text_w_73_), .Y(n4696) );
  INVX1 U22331 ( .A(top_core_io_Plain_text_w_72_), .Y(n4695) );
  INVX1 U22332 ( .A(top_core_io_operation), .Y(n4260) );
  XNOR2X1 U22333 ( .A(top_core_io_div_16_c_1_), .B(top_core_io_div_16_n5), .Y(
        top_core_io_div_16_N7) );
  XNOR2X1 U22334 ( .A(top_core_io_div_16_c_2_), .B(top_core_io_div_16_n2), .Y(
        top_core_io_div_16_N8) );
  INVX1 U22335 ( .A(top_core_io_n484), .Y(n4646) );
  AOI22X1 U22336 ( .A0(top_core_Ciphertext[7]), .A1(n3645), .B0(
        top_core_io_Data_reg_16__7_), .B1(n3672), .Y(top_core_io_n484) );
  INVX1 U22337 ( .A(top_core_io_n483), .Y(n4645) );
  AOI22X1 U22338 ( .A0(top_core_Ciphertext[6]), .A1(n3646), .B0(
        top_core_io_Data_reg_16__6_), .B1(n3672), .Y(top_core_io_n483) );
  INVX1 U22339 ( .A(top_core_io_n482), .Y(n4644) );
  AOI22X1 U22340 ( .A0(top_core_Ciphertext[5]), .A1(n3647), .B0(
        top_core_io_Data_reg_16__5_), .B1(n3671), .Y(top_core_io_n482) );
  INVX1 U22341 ( .A(top_core_io_n481), .Y(n4643) );
  AOI22X1 U22342 ( .A0(top_core_Ciphertext[4]), .A1(n3648), .B0(
        top_core_io_Data_reg_16__4_), .B1(n3671), .Y(top_core_io_n481) );
  INVX1 U22343 ( .A(top_core_io_n480), .Y(n4642) );
  AOI22X1 U22344 ( .A0(top_core_Ciphertext[3]), .A1(n3649), .B0(
        top_core_io_Data_reg_16__3_), .B1(n3670), .Y(top_core_io_n480) );
  INVX1 U22345 ( .A(top_core_io_n479), .Y(n4641) );
  AOI22X1 U22346 ( .A0(top_core_Ciphertext[2]), .A1(n3650), .B0(
        top_core_io_Data_reg_16__2_), .B1(n3670), .Y(top_core_io_n479) );
  INVX1 U22347 ( .A(top_core_io_n478), .Y(n4640) );
  AOI22X1 U22348 ( .A0(top_core_Ciphertext[1]), .A1(n3650), .B0(
        top_core_io_Data_reg_16__1_), .B1(n3669), .Y(top_core_io_n478) );
  INVX1 U22349 ( .A(top_core_io_n477), .Y(n4639) );
  AOI22X1 U22350 ( .A0(top_core_Ciphertext[0]), .A1(n3651), .B0(
        top_core_io_Data_reg_16__0_), .B1(n3669), .Y(top_core_io_n477) );
  INVX1 U22351 ( .A(top_core_io_n476), .Y(n4638) );
  AOI22X1 U22352 ( .A0(top_core_Ciphertext[15]), .A1(n3645), .B0(
        top_core_io_Data_reg_17__7_), .B1(n3668), .Y(top_core_io_n476) );
  INVX1 U22353 ( .A(top_core_io_n475), .Y(n4637) );
  AOI22X1 U22354 ( .A0(top_core_Ciphertext[14]), .A1(n3646), .B0(
        top_core_io_Data_reg_17__6_), .B1(n3668), .Y(top_core_io_n475) );
  INVX1 U22355 ( .A(top_core_io_n474), .Y(n4636) );
  AOI22X1 U22356 ( .A0(top_core_Ciphertext[13]), .A1(n3647), .B0(
        top_core_io_Data_reg_17__5_), .B1(n3667), .Y(top_core_io_n474) );
  INVX1 U22357 ( .A(top_core_io_n473), .Y(n4635) );
  AOI22X1 U22358 ( .A0(top_core_Ciphertext[12]), .A1(n3648), .B0(
        top_core_io_Data_reg_17__4_), .B1(n3667), .Y(top_core_io_n473) );
  INVX1 U22359 ( .A(top_core_io_n472), .Y(n4634) );
  AOI22X1 U22360 ( .A0(top_core_Ciphertext[11]), .A1(n3679), .B0(
        top_core_io_Data_reg_17__3_), .B1(n3668), .Y(top_core_io_n472) );
  INVX1 U22361 ( .A(top_core_io_n471), .Y(n4633) );
  AOI22X1 U22362 ( .A0(top_core_Ciphertext[10]), .A1(n3680), .B0(
        top_core_io_Data_reg_17__2_), .B1(n3663), .Y(top_core_io_n471) );
  INVX1 U22363 ( .A(top_core_io_n470), .Y(n4632) );
  AOI22X1 U22364 ( .A0(top_core_Ciphertext[9]), .A1(n3681), .B0(
        top_core_io_Data_reg_17__1_), .B1(n3666), .Y(top_core_io_n470) );
  INVX1 U22365 ( .A(top_core_io_n469), .Y(n4631) );
  AOI22X1 U22366 ( .A0(top_core_Ciphertext[8]), .A1(n3682), .B0(
        top_core_io_Data_reg_17__0_), .B1(n3677), .Y(top_core_io_n469) );
  INVX1 U22367 ( .A(top_core_io_n468), .Y(n4630) );
  AOI22X1 U22368 ( .A0(top_core_Ciphertext[23]), .A1(n3683), .B0(
        top_core_io_Data_reg_18__7_), .B1(n3672), .Y(top_core_io_n468) );
  INVX1 U22369 ( .A(top_core_io_n467), .Y(n4629) );
  AOI22X1 U22370 ( .A0(top_core_Ciphertext[22]), .A1(n3684), .B0(
        top_core_io_Data_reg_18__6_), .B1(n3671), .Y(top_core_io_n467) );
  INVX1 U22371 ( .A(top_core_io_n466), .Y(n4628) );
  AOI22X1 U22372 ( .A0(top_core_Ciphertext[21]), .A1(n3651), .B0(
        top_core_io_Data_reg_18__5_), .B1(n3653), .Y(top_core_io_n466) );
  INVX1 U22373 ( .A(top_core_io_n465), .Y(n4627) );
  AOI22X1 U22374 ( .A0(top_core_Ciphertext[20]), .A1(n3651), .B0(
        top_core_io_Data_reg_18__4_), .B1(n3653), .Y(top_core_io_n465) );
  INVX1 U22375 ( .A(top_core_io_n464), .Y(n4626) );
  AOI22X1 U22376 ( .A0(top_core_Ciphertext[19]), .A1(n3649), .B0(
        top_core_io_Data_reg_18__3_), .B1(n3655), .Y(top_core_io_n464) );
  INVX1 U22377 ( .A(top_core_io_n463), .Y(n4625) );
  AOI22X1 U22378 ( .A0(top_core_Ciphertext[18]), .A1(n3651), .B0(
        top_core_io_Data_reg_18__2_), .B1(n3665), .Y(top_core_io_n463) );
  INVX1 U22379 ( .A(top_core_io_n462), .Y(n4624) );
  AOI22X1 U22380 ( .A0(top_core_Ciphertext[17]), .A1(n3651), .B0(
        top_core_io_Data_reg_18__1_), .B1(n3654), .Y(top_core_io_n462) );
  INVX1 U22381 ( .A(top_core_io_n461), .Y(n4623) );
  AOI22X1 U22382 ( .A0(top_core_Ciphertext[16]), .A1(n3651), .B0(
        top_core_io_Data_reg_18__0_), .B1(n3686), .Y(top_core_io_n461) );
  INVX1 U22383 ( .A(top_core_io_n452), .Y(n4614) );
  AOI22X1 U22384 ( .A0(top_core_Ciphertext[39]), .A1(n3683), .B0(
        top_core_io_Data_reg_20__7_), .B1(n3669), .Y(top_core_io_n452) );
  INVX1 U22385 ( .A(top_core_io_n451), .Y(n4613) );
  AOI22X1 U22386 ( .A0(top_core_Ciphertext[38]), .A1(n3684), .B0(
        top_core_io_Data_reg_20__6_), .B1(n3672), .Y(top_core_io_n451) );
  INVX1 U22387 ( .A(top_core_io_n450), .Y(n4612) );
  AOI22X1 U22388 ( .A0(top_core_Ciphertext[37]), .A1(n3646), .B0(
        top_core_io_Data_reg_20__5_), .B1(n3666), .Y(top_core_io_n450) );
  INVX1 U22389 ( .A(top_core_io_n449), .Y(n4611) );
  AOI22X1 U22390 ( .A0(top_core_Ciphertext[36]), .A1(n3685), .B0(
        top_core_io_Data_reg_20__4_), .B1(n3666), .Y(top_core_io_n449) );
  INVX1 U22391 ( .A(top_core_io_n448), .Y(n4610) );
  AOI22X1 U22392 ( .A0(top_core_Ciphertext[35]), .A1(n3645), .B0(
        top_core_io_Data_reg_20__3_), .B1(n3675), .Y(top_core_io_n448) );
  INVX1 U22393 ( .A(top_core_io_n447), .Y(n4609) );
  AOI22X1 U22394 ( .A0(top_core_Ciphertext[34]), .A1(n3645), .B0(
        top_core_io_Data_reg_20__2_), .B1(n3676), .Y(top_core_io_n447) );
  INVX1 U22395 ( .A(top_core_io_n446), .Y(n4608) );
  AOI22X1 U22396 ( .A0(top_core_Ciphertext[33]), .A1(n3645), .B0(
        top_core_io_Data_reg_20__1_), .B1(n3659), .Y(top_core_io_n446) );
  INVX1 U22397 ( .A(top_core_io_n445), .Y(n4607) );
  AOI22X1 U22398 ( .A0(top_core_Ciphertext[32]), .A1(n3645), .B0(
        top_core_io_Data_reg_20__0_), .B1(n3658), .Y(top_core_io_n445) );
  INVX1 U22399 ( .A(top_core_io_n444), .Y(n4606) );
  AOI22X1 U22400 ( .A0(top_core_Ciphertext[47]), .A1(n3645), .B0(
        top_core_io_Data_reg_21__7_), .B1(n3664), .Y(top_core_io_n444) );
  INVX1 U22401 ( .A(top_core_io_n443), .Y(n4605) );
  AOI22X1 U22402 ( .A0(top_core_Ciphertext[46]), .A1(n3645), .B0(
        top_core_io_Data_reg_21__6_), .B1(n3663), .Y(top_core_io_n443) );
  INVX1 U22403 ( .A(top_core_io_n442), .Y(n4604) );
  AOI22X1 U22404 ( .A0(top_core_Ciphertext[45]), .A1(n3645), .B0(
        top_core_io_Data_reg_21__5_), .B1(n3667), .Y(top_core_io_n442) );
  INVX1 U22405 ( .A(top_core_io_n441), .Y(n4603) );
  AOI22X1 U22406 ( .A0(top_core_Ciphertext[44]), .A1(n3645), .B0(
        top_core_io_Data_reg_21__4_), .B1(n3656), .Y(top_core_io_n441) );
  INVX1 U22407 ( .A(top_core_io_n440), .Y(n4602) );
  AOI22X1 U22408 ( .A0(top_core_Ciphertext[43]), .A1(n3645), .B0(
        top_core_io_Data_reg_21__3_), .B1(n3671), .Y(top_core_io_n440) );
  INVX1 U22409 ( .A(top_core_io_n439), .Y(n4601) );
  AOI22X1 U22410 ( .A0(top_core_Ciphertext[42]), .A1(n3645), .B0(
        top_core_io_Data_reg_21__2_), .B1(n3670), .Y(top_core_io_n439) );
  INVX1 U22411 ( .A(top_core_io_n438), .Y(n4600) );
  AOI22X1 U22412 ( .A0(top_core_Ciphertext[41]), .A1(n3645), .B0(
        top_core_io_Data_reg_21__1_), .B1(n3657), .Y(top_core_io_n438) );
  INVX1 U22413 ( .A(top_core_io_n437), .Y(n4599) );
  AOI22X1 U22414 ( .A0(top_core_Ciphertext[40]), .A1(n3645), .B0(
        top_core_io_Data_reg_21__0_), .B1(n3662), .Y(top_core_io_n437) );
  INVX1 U22415 ( .A(top_core_io_n436), .Y(n4598) );
  AOI22X1 U22416 ( .A0(top_core_Ciphertext[55]), .A1(n3646), .B0(
        top_core_io_Data_reg_22__7_), .B1(n3674), .Y(top_core_io_n436) );
  INVX1 U22417 ( .A(top_core_io_n435), .Y(n4597) );
  AOI22X1 U22418 ( .A0(top_core_Ciphertext[54]), .A1(n3646), .B0(
        top_core_io_Data_reg_22__6_), .B1(n3660), .Y(top_core_io_n435) );
  INVX1 U22419 ( .A(top_core_io_n434), .Y(n4596) );
  AOI22X1 U22420 ( .A0(top_core_Ciphertext[53]), .A1(n3646), .B0(
        top_core_io_Data_reg_22__5_), .B1(n3656), .Y(top_core_io_n434) );
  INVX1 U22421 ( .A(top_core_io_n433), .Y(n4595) );
  AOI22X1 U22422 ( .A0(top_core_Ciphertext[52]), .A1(n3646), .B0(
        top_core_io_Data_reg_22__4_), .B1(n3674), .Y(top_core_io_n433) );
  INVX1 U22423 ( .A(top_core_io_n432), .Y(n4594) );
  AOI22X1 U22424 ( .A0(top_core_Ciphertext[51]), .A1(n3646), .B0(
        top_core_io_Data_reg_22__3_), .B1(n3659), .Y(top_core_io_n432) );
  INVX1 U22425 ( .A(top_core_io_n431), .Y(n4593) );
  AOI22X1 U22426 ( .A0(top_core_Ciphertext[50]), .A1(n3646), .B0(
        top_core_io_Data_reg_22__2_), .B1(n3658), .Y(top_core_io_n431) );
  INVX1 U22427 ( .A(top_core_io_n430), .Y(n4592) );
  AOI22X1 U22428 ( .A0(top_core_Ciphertext[49]), .A1(n3646), .B0(
        top_core_io_Data_reg_22__1_), .B1(n3665), .Y(top_core_io_n430) );
  INVX1 U22429 ( .A(top_core_io_n429), .Y(n4591) );
  AOI22X1 U22430 ( .A0(top_core_Ciphertext[48]), .A1(n3646), .B0(
        top_core_io_Data_reg_22__0_), .B1(n3665), .Y(top_core_io_n429) );
  INVX1 U22431 ( .A(top_core_io_n420), .Y(n4582) );
  AOI22X1 U22432 ( .A0(top_core_Ciphertext[71]), .A1(n3647), .B0(
        top_core_io_Data_reg_24__7_), .B1(n3674), .Y(top_core_io_n420) );
  INVX1 U22433 ( .A(top_core_io_n419), .Y(n4581) );
  AOI22X1 U22434 ( .A0(top_core_Ciphertext[70]), .A1(n3647), .B0(
        top_core_io_Data_reg_24__6_), .B1(n3675), .Y(top_core_io_n419) );
  INVX1 U22435 ( .A(top_core_io_n418), .Y(n4580) );
  AOI22X1 U22436 ( .A0(top_core_Ciphertext[69]), .A1(n3647), .B0(
        top_core_io_Data_reg_24__5_), .B1(n3654), .Y(top_core_io_n418) );
  INVX1 U22437 ( .A(top_core_io_n417), .Y(n4579) );
  AOI22X1 U22438 ( .A0(top_core_Ciphertext[68]), .A1(n3647), .B0(
        top_core_io_Data_reg_24__4_), .B1(n3654), .Y(top_core_io_n417) );
  INVX1 U22439 ( .A(top_core_io_n416), .Y(n4578) );
  AOI22X1 U22440 ( .A0(top_core_Ciphertext[67]), .A1(n3647), .B0(
        top_core_io_Data_reg_24__3_), .B1(n3667), .Y(top_core_io_n416) );
  INVX1 U22441 ( .A(top_core_io_n415), .Y(n4577) );
  AOI22X1 U22442 ( .A0(top_core_Ciphertext[66]), .A1(n3647), .B0(
        top_core_io_Data_reg_24__2_), .B1(n3655), .Y(top_core_io_n415) );
  INVX1 U22443 ( .A(top_core_io_n414), .Y(n4576) );
  AOI22X1 U22444 ( .A0(top_core_Ciphertext[65]), .A1(n3647), .B0(
        top_core_io_Data_reg_24__1_), .B1(n3659), .Y(top_core_io_n414) );
  INVX1 U22445 ( .A(top_core_io_n413), .Y(n4575) );
  AOI22X1 U22446 ( .A0(top_core_Ciphertext[64]), .A1(n3647), .B0(
        top_core_io_Data_reg_24__0_), .B1(n3662), .Y(top_core_io_n413) );
  INVX1 U22447 ( .A(top_core_io_n412), .Y(n4574) );
  AOI22X1 U22448 ( .A0(top_core_Ciphertext[79]), .A1(n3648), .B0(
        top_core_io_Data_reg_25__7_), .B1(n3662), .Y(top_core_io_n412) );
  INVX1 U22449 ( .A(top_core_io_n411), .Y(n4573) );
  AOI22X1 U22450 ( .A0(top_core_Ciphertext[78]), .A1(n3648), .B0(
        top_core_io_Data_reg_25__6_), .B1(n3662), .Y(top_core_io_n411) );
  INVX1 U22451 ( .A(top_core_io_n410), .Y(n4572) );
  AOI22X1 U22452 ( .A0(top_core_Ciphertext[77]), .A1(n3648), .B0(
        top_core_io_Data_reg_25__5_), .B1(n3661), .Y(top_core_io_n410) );
  INVX1 U22453 ( .A(top_core_io_n409), .Y(n4571) );
  AOI22X1 U22454 ( .A0(top_core_Ciphertext[76]), .A1(n3648), .B0(
        top_core_io_Data_reg_25__4_), .B1(n3661), .Y(top_core_io_n409) );
  INVX1 U22455 ( .A(top_core_io_n408), .Y(n4570) );
  AOI22X1 U22456 ( .A0(top_core_Ciphertext[75]), .A1(n3648), .B0(
        top_core_io_Data_reg_25__3_), .B1(n3660), .Y(top_core_io_n408) );
  INVX1 U22457 ( .A(top_core_io_n407), .Y(n4569) );
  AOI22X1 U22458 ( .A0(top_core_Ciphertext[74]), .A1(n3648), .B0(
        top_core_io_Data_reg_25__2_), .B1(n3660), .Y(top_core_io_n407) );
  INVX1 U22459 ( .A(top_core_io_n406), .Y(n4568) );
  AOI22X1 U22460 ( .A0(top_core_Ciphertext[73]), .A1(n3648), .B0(
        top_core_io_Data_reg_25__1_), .B1(n3670), .Y(top_core_io_n406) );
  INVX1 U22461 ( .A(top_core_io_n405), .Y(n4567) );
  AOI22X1 U22462 ( .A0(top_core_Ciphertext[72]), .A1(n3648), .B0(
        top_core_io_Data_reg_25__0_), .B1(n3669), .Y(top_core_io_n405) );
  INVX1 U22463 ( .A(top_core_io_n404), .Y(n4566) );
  AOI22X1 U22464 ( .A0(top_core_Ciphertext[87]), .A1(n3648), .B0(
        top_core_io_Data_reg_26__7_), .B1(n3652), .Y(top_core_io_n404) );
  INVX1 U22465 ( .A(top_core_io_n403), .Y(n4565) );
  AOI22X1 U22466 ( .A0(top_core_Ciphertext[86]), .A1(n3648), .B0(
        top_core_io_Data_reg_26__6_), .B1(n3672), .Y(top_core_io_n403) );
  INVX1 U22467 ( .A(top_core_io_n402), .Y(n4564) );
  AOI22X1 U22468 ( .A0(top_core_Ciphertext[85]), .A1(n3648), .B0(
        top_core_io_Data_reg_26__5_), .B1(n3666), .Y(top_core_io_n402) );
  INVX1 U22469 ( .A(top_core_io_n401), .Y(n4563) );
  AOI22X1 U22470 ( .A0(top_core_Ciphertext[84]), .A1(n3648), .B0(
        top_core_io_Data_reg_26__4_), .B1(n3673), .Y(top_core_io_n401) );
  INVX1 U22471 ( .A(top_core_io_n400), .Y(n4562) );
  AOI22X1 U22472 ( .A0(top_core_Ciphertext[83]), .A1(n3649), .B0(
        top_core_io_Data_reg_26__3_), .B1(n3661), .Y(top_core_io_n400) );
  INVX1 U22473 ( .A(top_core_io_n399), .Y(n4561) );
  AOI22X1 U22474 ( .A0(top_core_Ciphertext[82]), .A1(n3649), .B0(
        top_core_io_Data_reg_26__2_), .B1(n3665), .Y(top_core_io_n399) );
  INVX1 U22475 ( .A(top_core_io_n398), .Y(n4560) );
  AOI22X1 U22476 ( .A0(top_core_Ciphertext[81]), .A1(n3649), .B0(
        top_core_io_Data_reg_26__1_), .B1(n3652), .Y(top_core_io_n398) );
  INVX1 U22477 ( .A(top_core_io_n397), .Y(n4559) );
  AOI22X1 U22478 ( .A0(top_core_Ciphertext[80]), .A1(n3649), .B0(
        top_core_io_Data_reg_26__0_), .B1(n3686), .Y(top_core_io_n397) );
  INVX1 U22479 ( .A(top_core_io_n388), .Y(n4550) );
  AOI22X1 U22480 ( .A0(top_core_Ciphertext[103]), .A1(n3647), .B0(
        top_core_io_Data_reg_28__7_), .B1(n3659), .Y(top_core_io_n388) );
  INVX1 U22481 ( .A(top_core_io_n387), .Y(n4549) );
  AOI22X1 U22482 ( .A0(top_core_Ciphertext[102]), .A1(n3648), .B0(
        top_core_io_Data_reg_28__6_), .B1(n3659), .Y(top_core_io_n387) );
  INVX1 U22483 ( .A(top_core_io_n386), .Y(n4548) );
  AOI22X1 U22484 ( .A0(top_core_Ciphertext[101]), .A1(n3645), .B0(
        top_core_io_Data_reg_28__5_), .B1(n3658), .Y(top_core_io_n386) );
  INVX1 U22485 ( .A(top_core_io_n385), .Y(n4547) );
  AOI22X1 U22486 ( .A0(top_core_Ciphertext[100]), .A1(n3646), .B0(
        top_core_io_Data_reg_28__4_), .B1(n3658), .Y(top_core_io_n385) );
  INVX1 U22487 ( .A(top_core_io_n384), .Y(n4546) );
  AOI22X1 U22488 ( .A0(top_core_Ciphertext[99]), .A1(n3649), .B0(
        top_core_io_Data_reg_28__3_), .B1(n3657), .Y(top_core_io_n384) );
  INVX1 U22489 ( .A(top_core_io_n383), .Y(n4545) );
  AOI22X1 U22490 ( .A0(top_core_Ciphertext[98]), .A1(n3650), .B0(
        top_core_io_Data_reg_28__2_), .B1(n3657), .Y(top_core_io_n383) );
  INVX1 U22491 ( .A(top_core_io_n382), .Y(n4544) );
  AOI22X1 U22492 ( .A0(top_core_Ciphertext[97]), .A1(n3651), .B0(
        top_core_io_Data_reg_28__1_), .B1(n3664), .Y(top_core_io_n382) );
  INVX1 U22493 ( .A(top_core_io_n381), .Y(n4543) );
  AOI22X1 U22494 ( .A0(top_core_Ciphertext[96]), .A1(n3647), .B0(
        top_core_io_Data_reg_28__0_), .B1(n3668), .Y(top_core_io_n381) );
  INVX1 U22495 ( .A(top_core_io_n380), .Y(n4542) );
  AOI22X1 U22496 ( .A0(top_core_Ciphertext[111]), .A1(n3649), .B0(
        top_core_io_Data_reg_29__7_), .B1(n3676), .Y(top_core_io_n380) );
  INVX1 U22497 ( .A(top_core_io_n379), .Y(n4541) );
  AOI22X1 U22498 ( .A0(top_core_Ciphertext[110]), .A1(n3648), .B0(
        top_core_io_Data_reg_29__6_), .B1(n3673), .Y(top_core_io_n379) );
  INVX1 U22499 ( .A(top_core_io_n378), .Y(n4540) );
  AOI22X1 U22500 ( .A0(top_core_Ciphertext[109]), .A1(n3645), .B0(
        top_core_io_Data_reg_29__5_), .B1(n3657), .Y(top_core_io_n378) );
  INVX1 U22501 ( .A(top_core_io_n377), .Y(n4539) );
  AOI22X1 U22502 ( .A0(top_core_Ciphertext[108]), .A1(n3646), .B0(
        top_core_io_Data_reg_29__4_), .B1(n3660), .Y(top_core_io_n377) );
  INVX1 U22503 ( .A(top_core_io_n376), .Y(n4538) );
  AOI22X1 U22504 ( .A0(top_core_Ciphertext[107]), .A1(n3650), .B0(
        top_core_io_Data_reg_29__3_), .B1(n3656), .Y(top_core_io_n376) );
  INVX1 U22505 ( .A(top_core_io_n375), .Y(n4537) );
  AOI22X1 U22506 ( .A0(top_core_Ciphertext[106]), .A1(n3650), .B0(
        top_core_io_Data_reg_29__2_), .B1(n3656), .Y(top_core_io_n375) );
  INVX1 U22507 ( .A(top_core_io_n374), .Y(n4536) );
  AOI22X1 U22508 ( .A0(top_core_Ciphertext[105]), .A1(n3650), .B0(
        top_core_io_Data_reg_29__1_), .B1(n3655), .Y(top_core_io_n374) );
  INVX1 U22509 ( .A(top_core_io_n373), .Y(n4535) );
  AOI22X1 U22510 ( .A0(top_core_Ciphertext[104]), .A1(n3650), .B0(
        top_core_io_Data_reg_29__0_), .B1(n3655), .Y(top_core_io_n373) );
  INVX1 U22511 ( .A(top_core_io_n372), .Y(n4534) );
  AOI22X1 U22512 ( .A0(top_core_Ciphertext[119]), .A1(n3650), .B0(
        top_core_io_Data_reg_30__7_), .B1(n3674), .Y(top_core_io_n372) );
  INVX1 U22513 ( .A(top_core_io_n371), .Y(n4533) );
  AOI22X1 U22514 ( .A0(top_core_Ciphertext[118]), .A1(n3650), .B0(
        top_core_io_Data_reg_30__6_), .B1(n3678), .Y(top_core_io_n371) );
  INVX1 U22515 ( .A(top_core_io_n370), .Y(n4532) );
  AOI22X1 U22516 ( .A0(top_core_Ciphertext[117]), .A1(n3650), .B0(
        top_core_io_Data_reg_30__5_), .B1(n3654), .Y(top_core_io_n370) );
  INVX1 U22517 ( .A(top_core_io_n369), .Y(n4531) );
  AOI22X1 U22518 ( .A0(top_core_Ciphertext[116]), .A1(n3650), .B0(
        top_core_io_Data_reg_30__4_), .B1(n3654), .Y(top_core_io_n369) );
  INVX1 U22519 ( .A(top_core_io_n368), .Y(n4530) );
  AOI22X1 U22520 ( .A0(top_core_Ciphertext[115]), .A1(n3650), .B0(
        top_core_io_Data_reg_30__3_), .B1(n3653), .Y(top_core_io_n368) );
  INVX1 U22521 ( .A(top_core_io_n367), .Y(n4529) );
  AOI22X1 U22522 ( .A0(top_core_Ciphertext[114]), .A1(n3650), .B0(
        top_core_io_Data_reg_30__2_), .B1(n3653), .Y(top_core_io_n367) );
  INVX1 U22523 ( .A(top_core_io_n366), .Y(n4528) );
  AOI22X1 U22524 ( .A0(top_core_Ciphertext[113]), .A1(n3650), .B0(
        top_core_io_Data_reg_30__1_), .B1(n3652), .Y(top_core_io_n366) );
  INVX1 U22525 ( .A(top_core_io_n365), .Y(n4527) );
  AOI22X1 U22526 ( .A0(top_core_Ciphertext[112]), .A1(n3650), .B0(
        top_core_io_Data_reg_30__0_), .B1(n3652), .Y(top_core_io_n365) );
  NOR2X2 U22527 ( .A(n7023), .B(top_core_KE_Nk0_1_), .Y(top_core_KE_n894) );
  CLKINVX3 U22528 ( .A(top_core_Core_Full), .Y(n6308) );
  NOR2X1 U22529 ( .A(top_core_KE_n2702), .B(top_core_KE_n741), .Y(
        top_core_KE_n2700) );
  AOI221X1 U22530 ( .A0(top_core_KE_n896), .A1(top_core_KE_n2506), .B0(
        top_core_KE_n895), .B1(n7015), .C0(n7011), .Y(top_core_KE_n2702) );
  NOR3X1 U22531 ( .A(top_core_EC_n25), .B(n2431), .C(n4024), .Y(
        top_core_EC_n1014) );
  XOR2X1 U22532 ( .A(top_core_KE_rcon_reg_7_), .B(
        top_core_KE_new_sboxw_192_23_), .Y(top_core_KE_n1974) );
  OAI222XL U22533 ( .A0(n13206), .A1(n13207), .B0(n13208), .B1(n13209), .C0(
        n1340), .C1(n13210), .Y(top_core_KE_new_sboxw_192_23_) );
  AOI211X1 U22534 ( .A0(n13231), .A1(n1152), .B0(n13259), .C0(n13260), .Y(
        n13206) );
  AOI211X1 U22535 ( .A0(n6475), .A1(n13211), .B0(n13212), .C0(n13213), .Y(
        n13210) );
  XOR2X1 U22536 ( .A(top_core_KE_rcon_reg_0_), .B(
        top_core_KE_new_sboxw_192_16_), .Y(top_core_KE_n2002) );
  OAI22X1 U22537 ( .A0(n13491), .A1(n6990), .B0(n1340), .B1(n13492), .Y(
        top_core_KE_new_sboxw_192_16_) );
  AOI222X1 U22538 ( .A0(n13508), .A1(n1185), .B0(n6469), .B1(n13509), .C0(
        n1356), .C1(n13510), .Y(n13491) );
  AOI22X1 U22539 ( .A0(n1356), .A1(n13493), .B0(n13494), .B1(n1185), .Y(n13492) );
  XOR2X1 U22540 ( .A(top_core_KE_rcon_reg_2_), .B(
        top_core_KE_new_sboxw_192_18_), .Y(top_core_KE_n1994) );
  OAI222XL U22541 ( .A0(n13430), .A1(n13207), .B0(n13431), .B1(n13209), .C0(
        n1340), .C1(n13432), .Y(top_core_KE_new_sboxw_192_18_) );
  AOI221X1 U22542 ( .A0(n13403), .A1(n1685), .B0(n1667), .B1(n13448), .C0(
        n13449), .Y(n13431) );
  AOI221X1 U22543 ( .A0(n1667), .A1(n13456), .B0(n13457), .B1(n1668), .C0(
        n13458), .Y(n13430) );
  XOR2X1 U22544 ( .A(top_core_KE_rcon_reg_3_), .B(
        top_core_KE_new_sboxw_192_19_), .Y(top_core_KE_n1990) );
  OAI21XL U22545 ( .A0(n1340), .A1(n13396), .B0(n13397), .Y(
        top_core_KE_new_sboxw_192_19_) );
  AOI211X1 U22546 ( .A0(n13272), .A1(n13416), .B0(n6468), .C0(n13417), .Y(
        n13396) );
  AOI21X1 U22547 ( .A0(n6701), .A1(n13398), .B0(n13399), .Y(n13397) );
  XOR2X1 U22548 ( .A(top_core_KE_rcon_reg_1_), .B(
        top_core_KE_new_sboxw_192_17_), .Y(top_core_KE_n1998) );
  OAI2BB2X1 U22549 ( .B0(n1340), .B1(n13463), .A0N(n1340), .A1N(n13464), .Y(
        top_core_KE_new_sboxw_192_17_) );
  AOI222X1 U22550 ( .A0(n13479), .A1(n1185), .B0(n6475), .B1(n13480), .C0(
        n6469), .C1(n13481), .Y(n13463) );
  OAI221XL U22551 ( .A0(n13465), .A1(n13217), .B0(n1356), .B1(n13466), .C0(
        n13467), .Y(n13464) );
  XOR2X1 U22552 ( .A(top_core_KE_rcon_reg_4_), .B(
        top_core_KE_new_sboxw_192_20_), .Y(top_core_KE_n1986) );
  OAI21XL U22553 ( .A0(n13358), .A1(n6990), .B0(n13359), .Y(
        top_core_KE_new_sboxw_192_20_) );
  AOI222X1 U22554 ( .A0(n1356), .A1(n13377), .B0(n6462), .B1(n13378), .C0(
        n13272), .C1(n13379), .Y(n13358) );
  OAI2BB1X1 U22555 ( .A0N(n13360), .A1N(n13361), .B0(n6990), .Y(n13359) );
  XOR2X1 U22556 ( .A(top_core_KE_rcon_reg_5_), .B(
        top_core_KE_new_sboxw_192_21_), .Y(top_core_KE_n1982) );
  OAI222XL U22557 ( .A0(n13322), .A1(n13209), .B0(n1340), .B1(n13323), .C0(
        n13324), .C1(n13207), .Y(top_core_KE_new_sboxw_192_21_) );
  AOI222X1 U22558 ( .A0(n1667), .A1(n13325), .B0(n13326), .B1(n1671), .C0(
        n6472), .C1(n13327), .Y(n13324) );
  AOI22X1 U22559 ( .A0(n1356), .A1(n13331), .B0(n13332), .B1(n1185), .Y(n13323) );
  XOR2X1 U22560 ( .A(top_core_KE_rcon_reg_6_), .B(
        top_core_KE_new_sboxw_192_22_), .Y(top_core_KE_n1978) );
  OAI22X1 U22561 ( .A0(n1340), .A1(n13269), .B0(n13270), .B1(n6990), .Y(
        top_core_KE_new_sboxw_192_22_) );
  AOI211X1 U22562 ( .A0(n13298), .A1(n1185), .B0(n13299), .C0(n13300), .Y(
        n13269) );
  AOI221X1 U22563 ( .A0(n1356), .A1(n13271), .B0(n13272), .B1(n13273), .C0(
        n13274), .Y(n13270) );
  NOR2X1 U22564 ( .A(n7022), .B(top_core_KE_Nk0_2_), .Y(top_core_KE_n897) );
  OAI21X1 U22565 ( .A0(n7011), .A1(top_core_KE_n2696), .B0(n_RSTB), .Y(
        top_core_KE_n2175) );
  OAI222XL U22566 ( .A0(top_core_EC_n1011), .A1(n4195), .B0(top_core_EC_n1023), 
        .B1(top_core_EC_n1013), .C0(n4028), .C1(n1), .Y(top_core_EC_n1293) );
  AOI211X1 U22567 ( .A0(n4020), .A1(top_core_EC_n1021), .B0(top_core_EC_n1022), 
        .C0(top_core_EC_n1025), .Y(top_core_EC_n1023) );
  NOR3X1 U22568 ( .A(top_core_EC_n25), .B(n3989), .C(n2407), .Y(
        top_core_EC_n1025) );
  AND2X2 U22569 ( .A(top_core_KE_n2692), .B(top_core_KE_n728), .Y(
        top_core_KE_n2181) );
  NAND3X1 U22570 ( .A(n1), .B(top_core_EC_n1024), .C(top_core_Core_Full), .Y(
        top_core_EC_n1013) );
  NOR2X1 U22571 ( .A(n3563), .B(top_core_Core_Full), .Y(top_core_EC_n872) );
  OAI221XL U22572 ( .A0(n3984), .A1(n4028), .B0(n2520), .B1(n3985), .C0(
        top_core_EC_n1016), .Y(top_core_EC_n1015) );
  AOI22X1 U22573 ( .A0(n2393), .A1(top_core_EC_n25), .B0(top_core_EC_n864), 
        .B1(n4022), .Y(top_core_EC_n1016) );
  OAI221XL U22574 ( .A0(n3508), .A1(n4827), .B0(n3516), .B1(
        top_core_EC_ss_n207), .C0(top_core_EC_n858), .Y(top_core_EC_n1160) );
  INVX1 U22575 ( .A(top_core_EC_mix_out_2_), .Y(n4827) );
  AOI22X1 U22576 ( .A0(top_core_Plain_text[122]), .A1(n3526), .B0(
        top_core_EC_round_result_2_), .B1(n3541), .Y(top_core_EC_n858) );
  OAI221XL U22577 ( .A0(n3508), .A1(n4817), .B0(n3516), .B1(
        top_core_EC_ss_n174), .C0(top_core_EC_n855), .Y(top_core_EC_n1157) );
  INVX1 U22578 ( .A(top_core_EC_mix_out_5_), .Y(n4817) );
  AOI22X1 U22579 ( .A0(top_core_Plain_text[125]), .A1(n3526), .B0(
        top_core_EC_round_result_5_), .B1(n3541), .Y(top_core_EC_n855) );
  OAI221XL U22580 ( .A0(n3508), .A1(n4835), .B0(n3516), .B1(
        top_core_EC_ss_n152), .C0(top_core_EC_n853), .Y(top_core_EC_n1155) );
  INVX1 U22581 ( .A(top_core_EC_mix_out_7_), .Y(n4835) );
  AOI22X1 U22582 ( .A0(top_core_Plain_text[127]), .A1(n3526), .B0(
        top_core_EC_round_result_7_), .B1(n3541), .Y(top_core_EC_n853) );
  OAI221XL U22583 ( .A0(n3508), .A1(n4824), .B0(n3516), .B1(
        top_core_EC_ss_n246), .C0(top_core_EC_n850), .Y(top_core_EC_n1152) );
  INVX1 U22584 ( .A(top_core_EC_mix_out_10_), .Y(n4824) );
  AOI22X1 U22585 ( .A0(top_core_Plain_text[114]), .A1(n3526), .B0(
        top_core_EC_round_result_10_), .B1(n3540), .Y(top_core_EC_n850) );
  OAI221XL U22586 ( .A0(n3508), .A1(n4814), .B0(n3517), .B1(
        top_core_EC_ss_n225), .C0(top_core_EC_n847), .Y(top_core_EC_n1149) );
  INVX1 U22587 ( .A(top_core_EC_mix_out_13_), .Y(n4814) );
  AOI22X1 U22588 ( .A0(top_core_Plain_text[117]), .A1(n3527), .B0(
        top_core_EC_round_result_13_), .B1(n3540), .Y(top_core_EC_n847) );
  OAI221XL U22589 ( .A0(n3509), .A1(n4834), .B0(n3517), .B1(
        top_core_EC_ss_n223), .C0(top_core_EC_n845), .Y(top_core_EC_n1147) );
  INVX1 U22590 ( .A(top_core_EC_mix_out_15_), .Y(n4834) );
  AOI22X1 U22591 ( .A0(top_core_Plain_text[119]), .A1(n3527), .B0(
        top_core_EC_round_result_15_), .B1(n3540), .Y(top_core_EC_n845) );
  OAI221XL U22592 ( .A0(n3515), .A1(n4825), .B0(n3517), .B1(
        top_core_EC_ss_n220), .C0(top_core_EC_n842), .Y(top_core_EC_n1144) );
  INVX1 U22593 ( .A(top_core_EC_mix_out_18_), .Y(n4825) );
  AOI22X1 U22594 ( .A0(top_core_Plain_text[106]), .A1(n3527), .B0(
        top_core_EC_round_result_18_), .B1(n3540), .Y(top_core_EC_n842) );
  OAI221XL U22595 ( .A0(n3510), .A1(n4815), .B0(n3517), .B1(
        top_core_EC_ss_n216), .C0(top_core_EC_n839), .Y(top_core_EC_n1141) );
  INVX1 U22596 ( .A(top_core_EC_mix_out_21_), .Y(n4815) );
  AOI22X1 U22597 ( .A0(top_core_Plain_text[109]), .A1(n3527), .B0(
        top_core_EC_round_result_21_), .B1(n3539), .Y(top_core_EC_n839) );
  OAI221XL U22598 ( .A0(n3514), .A1(n4811), .B0(n3517), .B1(
        top_core_EC_ss_n214), .C0(top_core_EC_n837), .Y(top_core_EC_n1139) );
  INVX1 U22599 ( .A(top_core_EC_mix_out_23_), .Y(n4811) );
  AOI22X1 U22600 ( .A0(top_core_Plain_text[111]), .A1(n3527), .B0(
        top_core_EC_round_result_23_), .B1(n3539), .Y(top_core_EC_n837) );
  OAI221XL U22601 ( .A0(n3509), .A1(n4826), .B0(n3520), .B1(
        top_core_EC_ss_n211), .C0(top_core_EC_n834), .Y(top_core_EC_n1136) );
  INVX1 U22602 ( .A(top_core_EC_mix_out_26_), .Y(n4826) );
  AOI22X1 U22603 ( .A0(top_core_Plain_text[98]), .A1(n3528), .B0(
        top_core_EC_round_result_26_), .B1(n3539), .Y(top_core_EC_n834) );
  OAI221XL U22604 ( .A0(n3509), .A1(n4816), .B0(n3523), .B1(
        top_core_EC_ss_n208), .C0(top_core_EC_n831), .Y(top_core_EC_n1133) );
  INVX1 U22605 ( .A(top_core_EC_mix_out_29_), .Y(n4816) );
  AOI22X1 U22606 ( .A0(top_core_Plain_text[101]), .A1(n3528), .B0(
        top_core_EC_round_result_29_), .B1(n3539), .Y(top_core_EC_n831) );
  OAI221XL U22607 ( .A0(n3509), .A1(n4810), .B0(n3518), .B1(
        top_core_EC_ss_n205), .C0(top_core_EC_n829), .Y(top_core_EC_n1131) );
  INVX1 U22608 ( .A(top_core_EC_mix_out_31_), .Y(n4810) );
  AOI22X1 U22609 ( .A0(top_core_Plain_text[103]), .A1(n3528), .B0(
        top_core_EC_round_result_31_), .B1(n3539), .Y(top_core_EC_n829) );
  OAI221XL U22610 ( .A0(n3509), .A1(n4943), .B0(n3516), .B1(
        top_core_EC_ss_n202), .C0(top_core_EC_n826), .Y(top_core_EC_n1128) );
  INVX1 U22611 ( .A(top_core_EC_mix_out_34_), .Y(n4943) );
  AOI22X1 U22612 ( .A0(top_core_Plain_text[90]), .A1(n3528), .B0(
        top_core_EC_round_result_34_), .B1(n3538), .Y(top_core_EC_n826) );
  OAI221XL U22613 ( .A0(n3510), .A1(n4928), .B0(n3518), .B1(
        top_core_EC_ss_n199), .C0(top_core_EC_n823), .Y(top_core_EC_n1125) );
  INVX1 U22614 ( .A(top_core_EC_mix_out_37_), .Y(n4928) );
  AOI22X1 U22615 ( .A0(top_core_Plain_text[93]), .A1(n3526), .B0(
        top_core_EC_round_result_37_), .B1(n3538), .Y(top_core_EC_n823) );
  OAI221XL U22616 ( .A0(n3510), .A1(n4923), .B0(n3518), .B1(
        top_core_EC_ss_n197), .C0(top_core_EC_n821), .Y(top_core_EC_n1123) );
  INVX1 U22617 ( .A(top_core_EC_mix_out_39_), .Y(n4923) );
  AOI22X1 U22618 ( .A0(top_core_Plain_text[95]), .A1(n3529), .B0(
        top_core_EC_round_result_39_), .B1(n3538), .Y(top_core_EC_n821) );
  OAI221XL U22619 ( .A0(n3510), .A1(n4946), .B0(n3518), .B1(
        top_core_EC_ss_n193), .C0(top_core_EC_n818), .Y(top_core_EC_n1120) );
  INVX1 U22620 ( .A(top_core_EC_mix_out_42_), .Y(n4946) );
  AOI22X1 U22621 ( .A0(top_core_Plain_text[82]), .A1(n3532), .B0(
        top_core_EC_round_result_42_), .B1(n3538), .Y(top_core_EC_n818) );
  OAI221XL U22622 ( .A0(n3510), .A1(n4935), .B0(n3518), .B1(
        top_core_EC_ss_n190), .C0(top_core_EC_n815), .Y(top_core_EC_n1117) );
  INVX1 U22623 ( .A(top_core_EC_mix_out_45_), .Y(n4935) );
  AOI22X1 U22624 ( .A0(top_core_Plain_text[85]), .A1(n3526), .B0(
        top_core_EC_round_result_45_), .B1(n3537), .Y(top_core_EC_n815) );
  OAI221XL U22625 ( .A0(n3510), .A1(n4924), .B0(n3518), .B1(
        top_core_EC_ss_n188), .C0(top_core_EC_n813), .Y(top_core_EC_n1115) );
  INVX1 U22626 ( .A(top_core_EC_mix_out_47_), .Y(n4924) );
  AOI22X1 U22627 ( .A0(top_core_Plain_text[87]), .A1(n3533), .B0(
        top_core_EC_round_result_47_), .B1(n3537), .Y(top_core_EC_n813) );
  OAI221XL U22628 ( .A0(n3511), .A1(n4944), .B0(n3519), .B1(
        top_core_EC_ss_n184), .C0(top_core_EC_n810), .Y(top_core_EC_n1112) );
  INVX1 U22629 ( .A(top_core_EC_mix_out_50_), .Y(n4944) );
  AOI22X1 U22630 ( .A0(top_core_Plain_text[74]), .A1(n3529), .B0(
        top_core_EC_round_result_50_), .B1(n3537), .Y(top_core_EC_n810) );
  OAI221XL U22631 ( .A0(n3511), .A1(n4929), .B0(n3519), .B1(
        top_core_EC_ss_n181), .C0(top_core_EC_n807), .Y(top_core_EC_n1109) );
  INVX1 U22632 ( .A(top_core_EC_mix_out_53_), .Y(n4929) );
  AOI22X1 U22633 ( .A0(top_core_Plain_text[77]), .A1(n3529), .B0(
        top_core_EC_round_result_53_), .B1(n3537), .Y(top_core_EC_n807) );
  OAI221XL U22634 ( .A0(n3511), .A1(n4951), .B0(n3519), .B1(
        top_core_EC_ss_n179), .C0(top_core_EC_n805), .Y(top_core_EC_n1107) );
  INVX1 U22635 ( .A(top_core_EC_mix_out_55_), .Y(n4951) );
  AOI22X1 U22636 ( .A0(top_core_Plain_text[79]), .A1(n3529), .B0(
        top_core_EC_round_result_55_), .B1(n3537), .Y(top_core_EC_n805) );
  OAI221XL U22637 ( .A0(n3511), .A1(n4947), .B0(n3519), .B1(
        top_core_EC_ss_n176), .C0(top_core_EC_n802), .Y(top_core_EC_n1104) );
  AOI22X1 U22638 ( .A0(top_core_Plain_text[66]), .A1(n3529), .B0(
        top_core_EC_round_result_58_), .B1(n3536), .Y(top_core_EC_n802) );
  OAI221XL U22639 ( .A0(n3512), .A1(n4936), .B0(n3520), .B1(
        top_core_EC_ss_n172), .C0(top_core_EC_n799), .Y(top_core_EC_n1101) );
  AOI22X1 U22640 ( .A0(top_core_Plain_text[69]), .A1(n3530), .B0(
        top_core_EC_round_result_61_), .B1(n3536), .Y(top_core_EC_n799) );
  OAI221XL U22641 ( .A0(n3512), .A1(n4925), .B0(n3520), .B1(
        top_core_EC_ss_n170), .C0(top_core_EC_n797), .Y(top_core_EC_n1099) );
  AOI22X1 U22642 ( .A0(top_core_Plain_text[71]), .A1(n3530), .B0(
        top_core_EC_round_result_63_), .B1(n3536), .Y(top_core_EC_n797) );
  OAI221XL U22643 ( .A0(n3512), .A1(n4798), .B0(n3520), .B1(
        top_core_EC_ss_n167), .C0(top_core_EC_n794), .Y(top_core_EC_n1096) );
  AOI22X1 U22644 ( .A0(top_core_Plain_text[58]), .A1(n3530), .B0(
        top_core_EC_round_result_66_), .B1(n3536), .Y(top_core_EC_n794) );
  OAI221XL U22645 ( .A0(n3512), .A1(n4787), .B0(n3520), .B1(
        top_core_EC_ss_n164), .C0(top_core_EC_n791), .Y(top_core_EC_n1093) );
  AOI22X1 U22646 ( .A0(top_core_Plain_text[61]), .A1(n3530), .B0(
        top_core_EC_round_result_69_), .B1(n3541), .Y(top_core_EC_n791) );
  OAI221XL U22647 ( .A0(n3512), .A1(n4775), .B0(n3520), .B1(
        top_core_EC_ss_n161), .C0(top_core_EC_n789), .Y(top_core_EC_n1091) );
  AOI22X1 U22648 ( .A0(top_core_Plain_text[63]), .A1(n3530), .B0(
        top_core_EC_round_result_71_), .B1(n3535), .Y(top_core_EC_n789) );
  OAI221XL U22649 ( .A0(n3513), .A1(n4795), .B0(n3521), .B1(
        top_core_EC_ss_n158), .C0(top_core_EC_n786), .Y(top_core_EC_n1088) );
  AOI22X1 U22650 ( .A0(top_core_Plain_text[50]), .A1(n3531), .B0(
        top_core_EC_round_result_74_), .B1(n3540), .Y(top_core_EC_n786) );
  OAI221XL U22651 ( .A0(n3513), .A1(n4780), .B0(n3521), .B1(
        top_core_EC_ss_n155), .C0(top_core_EC_n783), .Y(top_core_EC_n1085) );
  AOI22X1 U22652 ( .A0(top_core_Plain_text[53]), .A1(n3531), .B0(
        top_core_EC_round_result_77_), .B1(n3534), .Y(top_core_EC_n783) );
  OAI221XL U22653 ( .A0(n3513), .A1(n4776), .B0(n3521), .B1(
        top_core_EC_ss_n153), .C0(top_core_EC_n781), .Y(top_core_EC_n1083) );
  AOI22X1 U22654 ( .A0(top_core_Plain_text[55]), .A1(n3531), .B0(
        top_core_EC_round_result_79_), .B1(top_core_EC_n733), .Y(
        top_core_EC_n781) );
  OAI221XL U22655 ( .A0(n3513), .A1(n4799), .B0(n3521), .B1(
        top_core_EC_ss_n149), .C0(top_core_EC_n778), .Y(top_core_EC_n1080) );
  AOI22X1 U22656 ( .A0(top_core_Plain_text[42]), .A1(n3531), .B0(
        top_core_EC_round_result_82_), .B1(top_core_EC_n733), .Y(
        top_core_EC_n778) );
  OAI221XL U22657 ( .A0(n3514), .A1(n4788), .B0(n3522), .B1(
        top_core_EC_ss_n146), .C0(top_core_EC_n775), .Y(top_core_EC_n1077) );
  AOI22X1 U22658 ( .A0(top_core_Plain_text[45]), .A1(n3532), .B0(
        top_core_EC_round_result_85_), .B1(n3541), .Y(top_core_EC_n775) );
  OAI221XL U22659 ( .A0(n3514), .A1(n4777), .B0(n3522), .B1(
        top_core_EC_ss_n144), .C0(top_core_EC_n773), .Y(top_core_EC_n1075) );
  AOI22X1 U22660 ( .A0(top_core_Plain_text[47]), .A1(n3532), .B0(
        top_core_EC_round_result_87_), .B1(n3541), .Y(top_core_EC_n773) );
  OAI221XL U22661 ( .A0(n3514), .A1(n4796), .B0(n3522), .B1(
        top_core_EC_ss_n140), .C0(top_core_EC_n770), .Y(top_core_EC_n1072) );
  AOI22X1 U22662 ( .A0(top_core_Plain_text[34]), .A1(n3532), .B0(
        top_core_EC_round_result_90_), .B1(n3541), .Y(top_core_EC_n770) );
  OAI221XL U22663 ( .A0(n3514), .A1(n4781), .B0(n3522), .B1(
        top_core_EC_ss_n137), .C0(top_core_EC_n767), .Y(top_core_EC_n1069) );
  AOI22X1 U22664 ( .A0(top_core_Plain_text[37]), .A1(n3532), .B0(
        top_core_EC_round_result_93_), .B1(n3535), .Y(top_core_EC_n767) );
  OAI221XL U22665 ( .A0(n3514), .A1(n4802), .B0(n3522), .B1(
        top_core_EC_ss_n135), .C0(top_core_EC_n765), .Y(top_core_EC_n1067) );
  AOI22X1 U22666 ( .A0(top_core_Plain_text[39]), .A1(n3532), .B0(
        top_core_EC_round_result_95_), .B1(n3535), .Y(top_core_EC_n765) );
  OAI221XL U22667 ( .A0(n3515), .A1(n5144), .B0(top_core_EC_n730), .B1(
        top_core_EC_ss_n132), .C0(top_core_EC_n762), .Y(top_core_EC_n1064) );
  AOI22X1 U22668 ( .A0(top_core_Plain_text[26]), .A1(n3533), .B0(
        top_core_EC_round_result_98_), .B1(n3535), .Y(top_core_EC_n762) );
  OAI221XL U22669 ( .A0(n3515), .A1(n5128), .B0(n3521), .B1(
        top_core_EC_ss_n255), .C0(top_core_EC_n759), .Y(top_core_EC_n1061) );
  AOI22X1 U22670 ( .A0(top_core_Plain_text[29]), .A1(n3533), .B0(
        top_core_EC_round_result_101_), .B1(n3535), .Y(top_core_EC_n759) );
  OAI221XL U22671 ( .A0(n3515), .A1(n5150), .B0(n3517), .B1(
        top_core_EC_ss_n253), .C0(top_core_EC_n757), .Y(top_core_EC_n1059) );
  AOI22X1 U22672 ( .A0(top_core_Plain_text[31]), .A1(n3533), .B0(
        top_core_EC_round_result_103_), .B1(n3535), .Y(top_core_EC_n757) );
  OAI221XL U22673 ( .A0(n3515), .A1(n5146), .B0(n3522), .B1(
        top_core_EC_ss_n250), .C0(top_core_EC_n754), .Y(top_core_EC_n1056) );
  AOI22X1 U22674 ( .A0(top_core_Plain_text[18]), .A1(n3533), .B0(
        top_core_EC_round_result_106_), .B1(n3534), .Y(top_core_EC_n754) );
  OAI221XL U22675 ( .A0(n3508), .A1(n5135), .B0(n3523), .B1(
        top_core_EC_ss_n247), .C0(top_core_EC_n751), .Y(top_core_EC_n1053) );
  AOI22X1 U22676 ( .A0(top_core_Plain_text[21]), .A1(n3527), .B0(
        top_core_EC_round_result_109_), .B1(n3539), .Y(top_core_EC_n751) );
  OAI221XL U22677 ( .A0(n3513), .A1(n5123), .B0(n3523), .B1(
        top_core_EC_ss_n244), .C0(top_core_EC_n749), .Y(top_core_EC_n1051) );
  AOI22X1 U22678 ( .A0(top_core_Plain_text[23]), .A1(n3528), .B0(
        top_core_EC_round_result_111_), .B1(n3537), .Y(top_core_EC_n749) );
  OAI221XL U22679 ( .A0(n3510), .A1(n5143), .B0(n3523), .B1(
        top_core_EC_ss_n241), .C0(top_core_EC_n746), .Y(top_core_EC_n1048) );
  AOI22X1 U22680 ( .A0(top_core_Plain_text[10]), .A1(n3531), .B0(
        top_core_EC_round_result_114_), .B1(n3538), .Y(top_core_EC_n746) );
  OAI221XL U22681 ( .A0(n3514), .A1(n5129), .B0(n3523), .B1(
        top_core_EC_ss_n238), .C0(top_core_EC_n743), .Y(top_core_EC_n1045) );
  AOI22X1 U22682 ( .A0(top_core_Plain_text[13]), .A1(n3533), .B0(
        top_core_EC_round_result_117_), .B1(n3534), .Y(top_core_EC_n743) );
  OAI221XL U22683 ( .A0(n3511), .A1(n5125), .B0(n3523), .B1(
        top_core_EC_ss_n236), .C0(top_core_EC_n741), .Y(top_core_EC_n1043) );
  AOI22X1 U22684 ( .A0(top_core_Plain_text[15]), .A1(n3526), .B0(
        top_core_EC_round_result_119_), .B1(n3534), .Y(top_core_EC_n741) );
  OAI221XL U22685 ( .A0(n3513), .A1(n5147), .B0(top_core_EC_n730), .B1(
        top_core_EC_ss_n232), .C0(top_core_EC_n738), .Y(top_core_EC_n1040) );
  AOI22X1 U22686 ( .A0(top_core_Plain_text[2]), .A1(n3529), .B0(
        top_core_EC_round_result_122_), .B1(n3534), .Y(top_core_EC_n738) );
  OAI221XL U22687 ( .A0(n3509), .A1(n5136), .B0(top_core_EC_n730), .B1(
        top_core_EC_ss_n229), .C0(top_core_EC_n735), .Y(top_core_EC_n1037) );
  AOI22X1 U22688 ( .A0(top_core_Plain_text[5]), .A1(n3532), .B0(
        top_core_EC_round_result_125_), .B1(n3534), .Y(top_core_EC_n735) );
  OAI221XL U22689 ( .A0(n3514), .A1(n5124), .B0(n3520), .B1(
        top_core_EC_ss_n227), .C0(top_core_EC_n731), .Y(top_core_EC_n1035) );
  AOI22X1 U22690 ( .A0(top_core_Plain_text[7]), .A1(n3530), .B0(
        top_core_EC_round_result_127_), .B1(n3534), .Y(top_core_EC_n731) );
  OAI221XL U22691 ( .A0(n3508), .A1(n4829), .B0(n3516), .B1(
        top_core_EC_ss_n218), .C0(top_core_EC_n859), .Y(top_core_EC_n1161) );
  INVX1 U22692 ( .A(top_core_EC_mix_out_1_), .Y(n4829) );
  AOI22X1 U22693 ( .A0(top_core_Plain_text[121]), .A1(n3526), .B0(
        top_core_EC_round_result_1_), .B1(n3541), .Y(top_core_EC_n859) );
  OAI221XL U22694 ( .A0(n3508), .A1(n4819), .B0(n3516), .B1(
        top_core_EC_ss_n185), .C0(top_core_EC_n856), .Y(top_core_EC_n1158) );
  INVX1 U22695 ( .A(top_core_EC_mix_out_4_), .Y(n4819) );
  AOI22X1 U22696 ( .A0(top_core_Plain_text[124]), .A1(n3526), .B0(
        top_core_EC_round_result_4_), .B1(n3541), .Y(top_core_EC_n856) );
  OAI221XL U22697 ( .A0(n3508), .A1(n4809), .B0(n3516), .B1(
        top_core_EC_ss_n163), .C0(top_core_EC_n854), .Y(top_core_EC_n1156) );
  INVX1 U22698 ( .A(top_core_EC_mix_out_6_), .Y(n4809) );
  AOI22X1 U22699 ( .A0(top_core_Plain_text[126]), .A1(n3526), .B0(
        top_core_EC_round_result_6_), .B1(n3541), .Y(top_core_EC_n854) );
  OAI221XL U22700 ( .A0(n3508), .A1(n4823), .B0(n3516), .B1(
        top_core_EC_ss_n130), .C0(top_core_EC_n851), .Y(top_core_EC_n1153) );
  INVX1 U22701 ( .A(top_core_EC_mix_out_9_), .Y(n4823) );
  AOI22X1 U22702 ( .A0(top_core_Plain_text[113]), .A1(n3526), .B0(
        top_core_EC_round_result_9_), .B1(n3540), .Y(top_core_EC_n851) );
  OAI221XL U22703 ( .A0(n3511), .A1(n4812), .B0(n3517), .B1(
        top_core_EC_ss_n226), .C0(top_core_EC_n848), .Y(top_core_EC_n1150) );
  INVX1 U22704 ( .A(top_core_EC_mix_out_12_), .Y(n4812) );
  AOI22X1 U22705 ( .A0(top_core_Plain_text[116]), .A1(n3527), .B0(
        top_core_EC_round_result_12_), .B1(n3540), .Y(top_core_EC_n848) );
  OAI221XL U22706 ( .A0(n3512), .A1(n4807), .B0(n3517), .B1(
        top_core_EC_ss_n224), .C0(top_core_EC_n846), .Y(top_core_EC_n1148) );
  INVX1 U22707 ( .A(top_core_EC_mix_out_14_), .Y(n4807) );
  AOI22X1 U22708 ( .A0(top_core_Plain_text[118]), .A1(n3527), .B0(
        top_core_EC_round_result_14_), .B1(n3540), .Y(top_core_EC_n846) );
  OAI221XL U22709 ( .A0(n3511), .A1(n4828), .B0(n3517), .B1(
        top_core_EC_ss_n221), .C0(top_core_EC_n843), .Y(top_core_EC_n1145) );
  INVX1 U22710 ( .A(top_core_EC_mix_out_17_), .Y(n4828) );
  AOI22X1 U22711 ( .A0(top_core_Plain_text[105]), .A1(n3527), .B0(
        top_core_EC_round_result_17_), .B1(n3540), .Y(top_core_EC_n843) );
  OAI221XL U22712 ( .A0(n3508), .A1(n4818), .B0(n3517), .B1(
        top_core_EC_ss_n217), .C0(top_core_EC_n840), .Y(top_core_EC_n1142) );
  INVX1 U22713 ( .A(top_core_EC_mix_out_20_), .Y(n4818) );
  AOI22X1 U22714 ( .A0(top_core_Plain_text[108]), .A1(n3527), .B0(
        top_core_EC_round_result_20_), .B1(n3539), .Y(top_core_EC_n840) );
  OAI221XL U22715 ( .A0(n3513), .A1(n4808), .B0(n3517), .B1(
        top_core_EC_ss_n215), .C0(top_core_EC_n838), .Y(top_core_EC_n1140) );
  INVX1 U22716 ( .A(top_core_EC_mix_out_22_), .Y(n4808) );
  AOI22X1 U22717 ( .A0(top_core_Plain_text[110]), .A1(n3527), .B0(
        top_core_EC_round_result_22_), .B1(n3539), .Y(top_core_EC_n838) );
  OAI221XL U22718 ( .A0(n3509), .A1(n4822), .B0(n3519), .B1(
        top_core_EC_ss_n212), .C0(top_core_EC_n835), .Y(top_core_EC_n1137) );
  INVX1 U22719 ( .A(top_core_EC_mix_out_25_), .Y(n4822) );
  AOI22X1 U22720 ( .A0(top_core_Plain_text[97]), .A1(n3528), .B0(
        top_core_EC_round_result_25_), .B1(n3539), .Y(top_core_EC_n835) );
  OAI221XL U22721 ( .A0(n3509), .A1(n4813), .B0(n3521), .B1(
        top_core_EC_ss_n209), .C0(top_core_EC_n832), .Y(top_core_EC_n1134) );
  INVX1 U22722 ( .A(top_core_EC_mix_out_28_), .Y(n4813) );
  AOI22X1 U22723 ( .A0(top_core_Plain_text[100]), .A1(n3528), .B0(
        top_core_EC_round_result_28_), .B1(n3539), .Y(top_core_EC_n832) );
  OAI221XL U22724 ( .A0(n3509), .A1(n4833), .B0(n3517), .B1(
        top_core_EC_ss_n206), .C0(top_core_EC_n830), .Y(top_core_EC_n1132) );
  INVX1 U22725 ( .A(top_core_EC_mix_out_30_), .Y(n4833) );
  AOI22X1 U22726 ( .A0(top_core_Plain_text[102]), .A1(n3528), .B0(
        top_core_EC_round_result_30_), .B1(n3539), .Y(top_core_EC_n830) );
  OAI221XL U22727 ( .A0(n3509), .A1(n4945), .B0(n3522), .B1(
        top_core_EC_ss_n203), .C0(top_core_EC_n827), .Y(top_core_EC_n1129) );
  INVX1 U22728 ( .A(top_core_EC_mix_out_33_), .Y(n4945) );
  AOI22X1 U22729 ( .A0(top_core_Plain_text[89]), .A1(n3528), .B0(
        top_core_EC_round_result_33_), .B1(n3538), .Y(top_core_EC_n827) );
  OAI221XL U22730 ( .A0(n3510), .A1(n4934), .B0(n3518), .B1(
        top_core_EC_ss_n200), .C0(top_core_EC_n824), .Y(top_core_EC_n1126) );
  INVX1 U22731 ( .A(top_core_EC_mix_out_36_), .Y(n4934) );
  AOI22X1 U22732 ( .A0(top_core_Plain_text[92]), .A1(n3526), .B0(
        top_core_EC_round_result_36_), .B1(n3538), .Y(top_core_EC_n824) );
  OAI221XL U22733 ( .A0(n3510), .A1(n4930), .B0(n3518), .B1(
        top_core_EC_ss_n198), .C0(top_core_EC_n822), .Y(top_core_EC_n1124) );
  INVX1 U22734 ( .A(top_core_EC_mix_out_38_), .Y(n4930) );
  AOI22X1 U22735 ( .A0(top_core_Plain_text[94]), .A1(n3530), .B0(
        top_core_EC_round_result_38_), .B1(n3538), .Y(top_core_EC_n822) );
  OAI221XL U22736 ( .A0(n3510), .A1(n4939), .B0(n3518), .B1(
        top_core_EC_ss_n194), .C0(top_core_EC_n819), .Y(top_core_EC_n1121) );
  INVX1 U22737 ( .A(top_core_EC_mix_out_41_), .Y(n4939) );
  AOI22X1 U22738 ( .A0(top_core_Plain_text[81]), .A1(n3527), .B0(
        top_core_EC_round_result_41_), .B1(n3538), .Y(top_core_EC_n819) );
  OAI221XL U22739 ( .A0(n3510), .A1(n4926), .B0(n3518), .B1(
        top_core_EC_ss_n191), .C0(top_core_EC_n816), .Y(top_core_EC_n1118) );
  INVX1 U22740 ( .A(top_core_EC_mix_out_44_), .Y(n4926) );
  AOI22X1 U22741 ( .A0(top_core_Plain_text[84]), .A1(n3528), .B0(
        top_core_EC_round_result_44_), .B1(n3537), .Y(top_core_EC_n816) );
  OAI221XL U22742 ( .A0(n3510), .A1(n4931), .B0(n3518), .B1(
        top_core_EC_ss_n189), .C0(top_core_EC_n814), .Y(top_core_EC_n1116) );
  INVX1 U22743 ( .A(top_core_EC_mix_out_46_), .Y(n4931) );
  AOI22X1 U22744 ( .A0(top_core_Plain_text[86]), .A1(n3531), .B0(
        top_core_EC_round_result_46_), .B1(n3537), .Y(top_core_EC_n814) );
  OAI221XL U22745 ( .A0(n3511), .A1(n4940), .B0(n3519), .B1(
        top_core_EC_ss_n186), .C0(top_core_EC_n811), .Y(top_core_EC_n1113) );
  INVX1 U22746 ( .A(top_core_EC_mix_out_49_), .Y(n4940) );
  AOI22X1 U22747 ( .A0(top_core_Plain_text[73]), .A1(n3529), .B0(
        top_core_EC_round_result_49_), .B1(n3537), .Y(top_core_EC_n811) );
  OAI221XL U22748 ( .A0(n3511), .A1(n4927), .B0(n3519), .B1(
        top_core_EC_ss_n182), .C0(top_core_EC_n808), .Y(top_core_EC_n1110) );
  INVX1 U22749 ( .A(top_core_EC_mix_out_52_), .Y(n4927) );
  AOI22X1 U22750 ( .A0(top_core_Plain_text[76]), .A1(n3529), .B0(
        top_core_EC_round_result_52_), .B1(n3537), .Y(top_core_EC_n808) );
  OAI221XL U22751 ( .A0(n3511), .A1(n4932), .B0(n3519), .B1(
        top_core_EC_ss_n180), .C0(top_core_EC_n806), .Y(top_core_EC_n1108) );
  INVX1 U22752 ( .A(top_core_EC_mix_out_54_), .Y(n4932) );
  AOI22X1 U22753 ( .A0(top_core_Plain_text[78]), .A1(n3529), .B0(
        top_core_EC_round_result_54_), .B1(n3537), .Y(top_core_EC_n806) );
  OAI221XL U22754 ( .A0(n3511), .A1(n4953), .B0(n3519), .B1(
        top_core_EC_ss_n177), .C0(top_core_EC_n803), .Y(top_core_EC_n1105) );
  INVX1 U22755 ( .A(top_core_EC_mix_out_57_), .Y(n4953) );
  AOI22X1 U22756 ( .A0(top_core_Plain_text[65]), .A1(n3529), .B0(
        top_core_EC_round_result_57_), .B1(n3536), .Y(top_core_EC_n803) );
  OAI221XL U22757 ( .A0(n3512), .A1(n4952), .B0(n3520), .B1(
        top_core_EC_ss_n173), .C0(top_core_EC_n800), .Y(top_core_EC_n1102) );
  AOI22X1 U22758 ( .A0(top_core_Plain_text[68]), .A1(n3530), .B0(
        top_core_EC_round_result_60_), .B1(n3536), .Y(top_core_EC_n800) );
  OAI221XL U22759 ( .A0(n3512), .A1(n4933), .B0(n3520), .B1(
        top_core_EC_ss_n171), .C0(top_core_EC_n798), .Y(top_core_EC_n1100) );
  AOI22X1 U22760 ( .A0(top_core_Plain_text[70]), .A1(n3530), .B0(
        top_core_EC_round_result_62_), .B1(n3536), .Y(top_core_EC_n798) );
  OAI221XL U22761 ( .A0(n3512), .A1(n4804), .B0(n3520), .B1(
        top_core_EC_ss_n168), .C0(top_core_EC_n795), .Y(top_core_EC_n1097) );
  AOI22X1 U22762 ( .A0(top_core_Plain_text[57]), .A1(n3530), .B0(
        top_core_EC_round_result_65_), .B1(n3536), .Y(top_core_EC_n795) );
  OAI221XL U22763 ( .A0(n3512), .A1(n4803), .B0(n3520), .B1(
        top_core_EC_ss_n165), .C0(top_core_EC_n792), .Y(top_core_EC_n1094) );
  AOI22X1 U22764 ( .A0(top_core_Plain_text[60]), .A1(n3530), .B0(
        top_core_EC_round_result_68_), .B1(n3539), .Y(top_core_EC_n792) );
  OAI221XL U22765 ( .A0(n3512), .A1(n4782), .B0(n3520), .B1(
        top_core_EC_ss_n162), .C0(top_core_EC_n790), .Y(top_core_EC_n1092) );
  AOI22X1 U22766 ( .A0(top_core_Plain_text[62]), .A1(n3530), .B0(
        top_core_EC_round_result_70_), .B1(n3537), .Y(top_core_EC_n790) );
  OAI221XL U22767 ( .A0(n3513), .A1(n4797), .B0(n3521), .B1(
        top_core_EC_ss_n159), .C0(top_core_EC_n787), .Y(top_core_EC_n1089) );
  AOI22X1 U22768 ( .A0(top_core_Plain_text[49]), .A1(n3531), .B0(
        top_core_EC_round_result_73_), .B1(n3536), .Y(top_core_EC_n787) );
  OAI221XL U22769 ( .A0(n3513), .A1(n4786), .B0(n3521), .B1(
        top_core_EC_ss_n156), .C0(top_core_EC_n784), .Y(top_core_EC_n1086) );
  AOI22X1 U22770 ( .A0(top_core_Plain_text[52]), .A1(n3531), .B0(
        top_core_EC_round_result_76_), .B1(n3538), .Y(top_core_EC_n784) );
  OAI221XL U22771 ( .A0(n3513), .A1(n4783), .B0(n3521), .B1(
        top_core_EC_ss_n154), .C0(top_core_EC_n782), .Y(top_core_EC_n1084) );
  AOI22X1 U22772 ( .A0(top_core_Plain_text[54]), .A1(n3531), .B0(
        top_core_EC_round_result_78_), .B1(n3541), .Y(top_core_EC_n782) );
  OAI221XL U22773 ( .A0(n3513), .A1(n4792), .B0(n3521), .B1(
        top_core_EC_ss_n150), .C0(top_core_EC_n779), .Y(top_core_EC_n1081) );
  AOI22X1 U22774 ( .A0(top_core_Plain_text[41]), .A1(n3531), .B0(
        top_core_EC_round_result_81_), .B1(n3535), .Y(top_core_EC_n779) );
  OAI221XL U22775 ( .A0(n3514), .A1(n4779), .B0(n3522), .B1(
        top_core_EC_ss_n147), .C0(top_core_EC_n776), .Y(top_core_EC_n1078) );
  AOI22X1 U22776 ( .A0(top_core_Plain_text[44]), .A1(n3532), .B0(
        top_core_EC_round_result_84_), .B1(n3540), .Y(top_core_EC_n776) );
  OAI221XL U22777 ( .A0(n3514), .A1(n4784), .B0(n3522), .B1(
        top_core_EC_ss_n145), .C0(top_core_EC_n774), .Y(top_core_EC_n1076) );
  AOI22X1 U22778 ( .A0(top_core_Plain_text[46]), .A1(n3532), .B0(
        top_core_EC_round_result_86_), .B1(n3534), .Y(top_core_EC_n774) );
  OAI221XL U22779 ( .A0(n3514), .A1(n4791), .B0(n3522), .B1(
        top_core_EC_ss_n142), .C0(top_core_EC_n771), .Y(top_core_EC_n1073) );
  AOI22X1 U22780 ( .A0(top_core_Plain_text[33]), .A1(n3532), .B0(
        top_core_EC_round_result_89_), .B1(n3536), .Y(top_core_EC_n771) );
  OAI221XL U22781 ( .A0(n3514), .A1(n4778), .B0(n3522), .B1(
        top_core_EC_ss_n138), .C0(top_core_EC_n768), .Y(top_core_EC_n1070) );
  AOI22X1 U22782 ( .A0(top_core_Plain_text[36]), .A1(n3532), .B0(
        top_core_EC_round_result_92_), .B1(n3535), .Y(top_core_EC_n768) );
  OAI221XL U22783 ( .A0(n3514), .A1(n4785), .B0(n3522), .B1(
        top_core_EC_ss_n136), .C0(top_core_EC_n766), .Y(top_core_EC_n1068) );
  AOI22X1 U22784 ( .A0(top_core_Plain_text[38]), .A1(n3532), .B0(
        top_core_EC_round_result_94_), .B1(n3535), .Y(top_core_EC_n766) );
  OAI221XL U22785 ( .A0(n3515), .A1(n5140), .B0(n3522), .B1(
        top_core_EC_ss_n133), .C0(top_core_EC_n763), .Y(top_core_EC_n1065) );
  AOI22X1 U22786 ( .A0(top_core_Plain_text[25]), .A1(n3533), .B0(
        top_core_EC_round_result_97_), .B1(n3535), .Y(top_core_EC_n763) );
  OAI221XL U22787 ( .A0(n3515), .A1(n5126), .B0(n3520), .B1(
        top_core_EC_ss_n256), .C0(top_core_EC_n760), .Y(top_core_EC_n1062) );
  AOI22X1 U22788 ( .A0(top_core_Plain_text[28]), .A1(n3533), .B0(
        top_core_EC_round_result_100_), .B1(n3535), .Y(top_core_EC_n760) );
  OAI221XL U22789 ( .A0(n3515), .A1(n5130), .B0(n3523), .B1(
        top_core_EC_ss_n254), .C0(top_core_EC_n758), .Y(top_core_EC_n1060) );
  AOI22X1 U22790 ( .A0(top_core_Plain_text[30]), .A1(n3533), .B0(
        top_core_EC_round_result_102_), .B1(n3535), .Y(top_core_EC_n758) );
  OAI221XL U22791 ( .A0(n3515), .A1(n5152), .B0(n3518), .B1(
        top_core_EC_ss_n251), .C0(top_core_EC_n755), .Y(top_core_EC_n1057) );
  AOI22X1 U22792 ( .A0(top_core_Plain_text[17]), .A1(n3533), .B0(
        top_core_EC_round_result_105_), .B1(n3541), .Y(top_core_EC_n755) );
  OAI221XL U22793 ( .A0(n3512), .A1(n5151), .B0(n3523), .B1(
        top_core_EC_ss_n248), .C0(top_core_EC_n752), .Y(top_core_EC_n1054) );
  AOI22X1 U22794 ( .A0(top_core_Plain_text[20]), .A1(n3530), .B0(
        top_core_EC_round_result_108_), .B1(n3536), .Y(top_core_EC_n752) );
  OAI221XL U22795 ( .A0(n3508), .A1(n5131), .B0(n3523), .B1(
        top_core_EC_ss_n245), .C0(top_core_EC_n750), .Y(top_core_EC_n1052) );
  AOI22X1 U22796 ( .A0(top_core_Plain_text[22]), .A1(n3527), .B0(
        top_core_EC_round_result_110_), .B1(n3535), .Y(top_core_EC_n750) );
  OAI221XL U22797 ( .A0(n3513), .A1(n5145), .B0(n3523), .B1(
        top_core_EC_ss_n242), .C0(top_core_EC_n747), .Y(top_core_EC_n1049) );
  AOI22X1 U22798 ( .A0(top_core_Plain_text[9]), .A1(n3528), .B0(
        top_core_EC_round_result_113_), .B1(n3540), .Y(top_core_EC_n747) );
  OAI221XL U22799 ( .A0(n3509), .A1(n5134), .B0(n3523), .B1(
        top_core_EC_ss_n239), .C0(top_core_EC_n744), .Y(top_core_EC_n1046) );
  AOI22X1 U22800 ( .A0(top_core_Plain_text[12]), .A1(n3531), .B0(
        top_core_EC_round_result_116_), .B1(n3534), .Y(top_core_EC_n744) );
  OAI221XL U22801 ( .A0(n3515), .A1(n5132), .B0(n3523), .B1(
        top_core_EC_ss_n237), .C0(top_core_EC_n742), .Y(top_core_EC_n1044) );
  AOI22X1 U22802 ( .A0(top_core_Plain_text[14]), .A1(n3529), .B0(
        top_core_EC_round_result_118_), .B1(n3534), .Y(top_core_EC_n742) );
  OAI221XL U22803 ( .A0(n3515), .A1(n5139), .B0(n3523), .B1(
        top_core_EC_ss_n233), .C0(top_core_EC_n739), .Y(top_core_EC_n1041) );
  AOI22X1 U22804 ( .A0(top_core_Plain_text[1]), .A1(n3533), .B0(
        top_core_EC_round_result_121_), .B1(n3534), .Y(top_core_EC_n739) );
  OAI221XL U22805 ( .A0(n3510), .A1(n5127), .B0(n3518), .B1(
        top_core_EC_ss_n230), .C0(top_core_EC_n736), .Y(top_core_EC_n1038) );
  AOI22X1 U22806 ( .A0(top_core_Plain_text[4]), .A1(n3530), .B0(
        top_core_EC_round_result_124_), .B1(n3534), .Y(top_core_EC_n736) );
  OAI221XL U22807 ( .A0(n3511), .A1(n5133), .B0(n3516), .B1(
        top_core_EC_ss_n228), .C0(top_core_EC_n734), .Y(top_core_EC_n1036) );
  AOI22X1 U22808 ( .A0(top_core_Plain_text[6]), .A1(n3527), .B0(
        top_core_EC_round_result_126_), .B1(n3534), .Y(top_core_EC_n734) );
  OAI221XL U22809 ( .A0(n3508), .A1(n4840), .B0(n3516), .B1(
        top_core_EC_ss_n257), .C0(top_core_EC_n860), .Y(top_core_EC_n1162) );
  INVX1 U22810 ( .A(top_core_EC_mix_out_0_), .Y(n4840) );
  AOI22X1 U22811 ( .A0(top_core_Plain_text[120]), .A1(n3526), .B0(
        top_core_EC_round_result_0_), .B1(n3541), .Y(top_core_EC_n860) );
  OAI221XL U22812 ( .A0(n3508), .A1(n4831), .B0(n3516), .B1(
        top_core_EC_ss_n141), .C0(top_core_EC_n852), .Y(top_core_EC_n1154) );
  INVX1 U22813 ( .A(top_core_EC_mix_out_8_), .Y(n4831) );
  AOI22X1 U22814 ( .A0(top_core_Plain_text[112]), .A1(n3526), .B0(
        top_core_EC_round_result_8_), .B1(n3540), .Y(top_core_EC_n852) );
  OAI221XL U22815 ( .A0(n3509), .A1(n4839), .B0(n3517), .B1(
        top_core_EC_ss_n222), .C0(top_core_EC_n844), .Y(top_core_EC_n1146) );
  INVX1 U22816 ( .A(top_core_EC_mix_out_16_), .Y(n4839) );
  AOI22X1 U22817 ( .A0(top_core_Plain_text[104]), .A1(n3527), .B0(
        top_core_EC_round_result_16_), .B1(n3540), .Y(top_core_EC_n844) );
  OAI221XL U22818 ( .A0(n3509), .A1(n4830), .B0(n3520), .B1(
        top_core_EC_ss_n213), .C0(top_core_EC_n836), .Y(top_core_EC_n1138) );
  INVX1 U22819 ( .A(top_core_EC_mix_out_24_), .Y(n4830) );
  AOI22X1 U22820 ( .A0(top_core_Plain_text[96]), .A1(n3528), .B0(
        top_core_EC_round_result_24_), .B1(n3539), .Y(top_core_EC_n836) );
  OAI221XL U22821 ( .A0(n3509), .A1(n4954), .B0(n3523), .B1(
        top_core_EC_ss_n204), .C0(top_core_EC_n828), .Y(top_core_EC_n1130) );
  INVX1 U22822 ( .A(top_core_EC_mix_out_32_), .Y(n4954) );
  AOI22X1 U22823 ( .A0(top_core_Plain_text[88]), .A1(n3528), .B0(
        top_core_EC_round_result_32_), .B1(n3538), .Y(top_core_EC_n828) );
  OAI221XL U22824 ( .A0(n3510), .A1(n4948), .B0(n3518), .B1(
        top_core_EC_ss_n195), .C0(top_core_EC_n820), .Y(top_core_EC_n1122) );
  INVX1 U22825 ( .A(top_core_EC_mix_out_40_), .Y(n4948) );
  AOI22X1 U22826 ( .A0(top_core_Plain_text[80]), .A1(n3529), .B0(
        top_core_EC_round_result_40_), .B1(n3538), .Y(top_core_EC_n820) );
  OAI221XL U22827 ( .A0(n3511), .A1(n4949), .B0(n3519), .B1(
        top_core_EC_ss_n187), .C0(top_core_EC_n812), .Y(top_core_EC_n1114) );
  INVX1 U22828 ( .A(top_core_EC_mix_out_48_), .Y(n4949) );
  AOI22X1 U22829 ( .A0(top_core_Plain_text[72]), .A1(n3529), .B0(
        top_core_EC_round_result_48_), .B1(n3537), .Y(top_core_EC_n812) );
  OAI221XL U22830 ( .A0(n3511), .A1(n4956), .B0(n3519), .B1(
        top_core_EC_ss_n178), .C0(top_core_EC_n804), .Y(top_core_EC_n1106) );
  INVX1 U22831 ( .A(top_core_EC_mix_out_56_), .Y(n4956) );
  AOI22X1 U22832 ( .A0(top_core_Plain_text[64]), .A1(n3529), .B0(
        top_core_EC_round_result_56_), .B1(n3536), .Y(top_core_EC_n804) );
  OAI221XL U22833 ( .A0(n3512), .A1(n4806), .B0(n3520), .B1(
        top_core_EC_ss_n169), .C0(top_core_EC_n796), .Y(top_core_EC_n1098) );
  AOI22X1 U22834 ( .A0(top_core_Plain_text[56]), .A1(n3530), .B0(
        top_core_EC_round_result_64_), .B1(n3536), .Y(top_core_EC_n796) );
  OAI221XL U22835 ( .A0(n3513), .A1(n4805), .B0(n3521), .B1(
        top_core_EC_ss_n160), .C0(top_core_EC_n788), .Y(top_core_EC_n1090) );
  AOI22X1 U22836 ( .A0(top_core_Plain_text[48]), .A1(n3531), .B0(
        top_core_EC_round_result_72_), .B1(n3535), .Y(top_core_EC_n788) );
  OAI221XL U22837 ( .A0(n3513), .A1(n4800), .B0(n3521), .B1(
        top_core_EC_ss_n151), .C0(top_core_EC_n780), .Y(top_core_EC_n1082) );
  AOI22X1 U22838 ( .A0(top_core_Plain_text[40]), .A1(n3531), .B0(
        top_core_EC_round_result_80_), .B1(n3539), .Y(top_core_EC_n780) );
  OAI221XL U22839 ( .A0(n3514), .A1(n4801), .B0(n3522), .B1(
        top_core_EC_ss_n143), .C0(top_core_EC_n772), .Y(top_core_EC_n1074) );
  AOI22X1 U22840 ( .A0(top_core_Plain_text[32]), .A1(n3532), .B0(
        top_core_EC_round_result_88_), .B1(n3537), .Y(top_core_EC_n772) );
  OAI221XL U22841 ( .A0(n3515), .A1(n5149), .B0(n3516), .B1(
        top_core_EC_ss_n134), .C0(top_core_EC_n764), .Y(top_core_EC_n1066) );
  AOI22X1 U22842 ( .A0(top_core_Plain_text[24]), .A1(n3533), .B0(
        top_core_EC_round_result_96_), .B1(n3535), .Y(top_core_EC_n764) );
  OAI221XL U22843 ( .A0(n3515), .A1(n5154), .B0(n3519), .B1(
        top_core_EC_ss_n252), .C0(top_core_EC_n756), .Y(top_core_EC_n1058) );
  AOI22X1 U22844 ( .A0(top_core_Plain_text[16]), .A1(n3533), .B0(
        top_core_EC_round_result_104_), .B1(n3534), .Y(top_core_EC_n756) );
  OAI221XL U22845 ( .A0(n3510), .A1(n5153), .B0(n3523), .B1(
        top_core_EC_ss_n243), .C0(top_core_EC_n748), .Y(top_core_EC_n1050) );
  AOI22X1 U22846 ( .A0(top_core_Plain_text[8]), .A1(n3532), .B0(
        top_core_EC_round_result_112_), .B1(n3539), .Y(top_core_EC_n748) );
  OAI221XL U22847 ( .A0(n3512), .A1(n5148), .B0(n3519), .B1(
        top_core_EC_ss_n234), .C0(top_core_EC_n740), .Y(top_core_EC_n1042) );
  AOI22X1 U22848 ( .A0(top_core_Plain_text[0]), .A1(n3528), .B0(
        top_core_EC_round_result_120_), .B1(n3534), .Y(top_core_EC_n740) );
  OAI221XL U22849 ( .A0(n3508), .A1(n4838), .B0(n3516), .B1(
        top_core_EC_ss_n196), .C0(top_core_EC_n857), .Y(top_core_EC_n1159) );
  INVX1 U22850 ( .A(top_core_EC_mix_out_3_), .Y(n4838) );
  AOI22X1 U22851 ( .A0(top_core_Plain_text[123]), .A1(n3526), .B0(
        top_core_EC_round_result_3_), .B1(n3541), .Y(top_core_EC_n857) );
  OAI221XL U22852 ( .A0(n3508), .A1(n4820), .B0(n3516), .B1(
        top_core_EC_ss_n235), .C0(top_core_EC_n849), .Y(top_core_EC_n1151) );
  INVX1 U22853 ( .A(top_core_EC_mix_out_11_), .Y(n4820) );
  AOI22X1 U22854 ( .A0(top_core_Plain_text[115]), .A1(n3526), .B0(
        top_core_EC_round_result_11_), .B1(n3540), .Y(top_core_EC_n849) );
  OAI221XL U22855 ( .A0(n3515), .A1(n4837), .B0(n3517), .B1(
        top_core_EC_ss_n219), .C0(top_core_EC_n841), .Y(top_core_EC_n1143) );
  INVX1 U22856 ( .A(top_core_EC_mix_out_19_), .Y(n4837) );
  AOI22X1 U22857 ( .A0(top_core_Plain_text[107]), .A1(n3527), .B0(
        top_core_EC_round_result_19_), .B1(n3540), .Y(top_core_EC_n841) );
  OAI221XL U22858 ( .A0(n3509), .A1(n4821), .B0(n3518), .B1(
        top_core_EC_ss_n210), .C0(top_core_EC_n833), .Y(top_core_EC_n1135) );
  INVX1 U22859 ( .A(top_core_EC_mix_out_27_), .Y(n4821) );
  AOI22X1 U22860 ( .A0(top_core_Plain_text[99]), .A1(n3528), .B0(
        top_core_EC_round_result_27_), .B1(n3539), .Y(top_core_EC_n833) );
  OAI221XL U22861 ( .A0(n3509), .A1(n4941), .B0(n3516), .B1(
        top_core_EC_ss_n201), .C0(top_core_EC_n825), .Y(top_core_EC_n1127) );
  INVX1 U22862 ( .A(top_core_EC_mix_out_35_), .Y(n4941) );
  AOI22X1 U22863 ( .A0(top_core_Plain_text[91]), .A1(n3528), .B0(
        top_core_EC_round_result_35_), .B1(n3538), .Y(top_core_EC_n825) );
  OAI221XL U22864 ( .A0(n3510), .A1(n4937), .B0(n3518), .B1(
        top_core_EC_ss_n192), .C0(top_core_EC_n817), .Y(top_core_EC_n1119) );
  INVX1 U22865 ( .A(top_core_EC_mix_out_43_), .Y(n4937) );
  AOI22X1 U22866 ( .A0(top_core_Plain_text[83]), .A1(n3532), .B0(
        top_core_EC_round_result_43_), .B1(n3538), .Y(top_core_EC_n817) );
  OAI221XL U22867 ( .A0(n3511), .A1(n4938), .B0(n3519), .B1(
        top_core_EC_ss_n183), .C0(top_core_EC_n809), .Y(top_core_EC_n1111) );
  INVX1 U22868 ( .A(top_core_EC_mix_out_51_), .Y(n4938) );
  AOI22X1 U22869 ( .A0(top_core_Plain_text[75]), .A1(n3529), .B0(
        top_core_EC_round_result_51_), .B1(n3537), .Y(top_core_EC_n809) );
  OAI221XL U22870 ( .A0(n3511), .A1(n4942), .B0(n3519), .B1(
        top_core_EC_ss_n175), .C0(top_core_EC_n801), .Y(top_core_EC_n1103) );
  AOI22X1 U22871 ( .A0(top_core_Plain_text[67]), .A1(n3529), .B0(
        top_core_EC_round_result_59_), .B1(n3536), .Y(top_core_EC_n801) );
  OAI221XL U22872 ( .A0(n3512), .A1(n4793), .B0(n3520), .B1(
        top_core_EC_ss_n166), .C0(top_core_EC_n793), .Y(top_core_EC_n1095) );
  AOI22X1 U22873 ( .A0(top_core_Plain_text[59]), .A1(n3530), .B0(
        top_core_EC_round_result_67_), .B1(n3536), .Y(top_core_EC_n793) );
  OAI221XL U22874 ( .A0(n3513), .A1(n4794), .B0(n3521), .B1(
        top_core_EC_ss_n157), .C0(top_core_EC_n785), .Y(top_core_EC_n1087) );
  AOI22X1 U22875 ( .A0(top_core_Plain_text[51]), .A1(n3531), .B0(
        top_core_EC_round_result_75_), .B1(n3540), .Y(top_core_EC_n785) );
  OAI221XL U22876 ( .A0(n3513), .A1(n4789), .B0(n3521), .B1(
        top_core_EC_ss_n148), .C0(top_core_EC_n777), .Y(top_core_EC_n1079) );
  AOI22X1 U22877 ( .A0(top_core_Plain_text[43]), .A1(n3531), .B0(
        top_core_EC_round_result_83_), .B1(n3536), .Y(top_core_EC_n777) );
  OAI221XL U22878 ( .A0(n3514), .A1(n4790), .B0(n3522), .B1(
        top_core_EC_ss_n139), .C0(top_core_EC_n769), .Y(top_core_EC_n1071) );
  AOI22X1 U22879 ( .A0(top_core_Plain_text[35]), .A1(n3532), .B0(
        top_core_EC_round_result_91_), .B1(n3538), .Y(top_core_EC_n769) );
  OAI221XL U22880 ( .A0(n3515), .A1(n5138), .B0(n3521), .B1(
        top_core_EC_ss_n131), .C0(top_core_EC_n761), .Y(top_core_EC_n1063) );
  AOI22X1 U22881 ( .A0(top_core_Plain_text[27]), .A1(n3533), .B0(
        top_core_EC_round_result_99_), .B1(n3535), .Y(top_core_EC_n761) );
  OAI221XL U22882 ( .A0(n3515), .A1(n5141), .B0(n3517), .B1(
        top_core_EC_ss_n249), .C0(top_core_EC_n753), .Y(top_core_EC_n1055) );
  AOI22X1 U22883 ( .A0(top_core_Plain_text[19]), .A1(n3533), .B0(
        top_core_EC_round_result_107_), .B1(n3537), .Y(top_core_EC_n753) );
  OAI221XL U22884 ( .A0(n3514), .A1(n5142), .B0(n3523), .B1(
        top_core_EC_ss_n240), .C0(top_core_EC_n745), .Y(top_core_EC_n1047) );
  AOI22X1 U22885 ( .A0(top_core_Plain_text[11]), .A1(n3533), .B0(
        top_core_EC_round_result_115_), .B1(n3538), .Y(top_core_EC_n745) );
  OAI221XL U22886 ( .A0(n3512), .A1(n5137), .B0(n3522), .B1(
        top_core_EC_ss_n231), .C0(top_core_EC_n737), .Y(top_core_EC_n1039) );
  AOI22X1 U22887 ( .A0(top_core_Plain_text[3]), .A1(n3531), .B0(
        top_core_EC_round_result_123_), .B1(n3534), .Y(top_core_EC_n737) );
  OAI221XL U22888 ( .A0(n4212), .A1(n3567), .B0(n6260), .B1(n3569), .C0(
        top_core_EC_n964), .Y(top_core_EC_n1246) );
  INVX1 U22889 ( .A(top_core_Plain_text[84]), .Y(n4212) );
  AOI22X1 U22890 ( .A0(n3574), .A1(top_core_EC_mix_out_44_), .B0(
        top_core_EC_add_out_r_44_), .B1(n3580), .Y(top_core_EC_n964) );
  OAI221XL U22891 ( .A0(n4213), .A1(n3567), .B0(n6259), .B1(n3569), .C0(
        top_core_EC_n963), .Y(top_core_EC_n1245) );
  INVX1 U22892 ( .A(top_core_Plain_text[85]), .Y(n4213) );
  AOI22X1 U22893 ( .A0(n3575), .A1(top_core_EC_mix_out_45_), .B0(
        top_core_EC_add_out_r_45_), .B1(n3580), .Y(top_core_EC_n963) );
  OAI221XL U22894 ( .A0(n4214), .A1(n3567), .B0(n6258), .B1(n3569), .C0(
        top_core_EC_n962), .Y(top_core_EC_n1244) );
  INVX1 U22895 ( .A(top_core_Plain_text[86]), .Y(n4214) );
  AOI22X1 U22896 ( .A0(n3576), .A1(top_core_EC_mix_out_46_), .B0(
        top_core_EC_add_out_r_46_), .B1(n3580), .Y(top_core_EC_n962) );
  OAI221XL U22897 ( .A0(n4215), .A1(n3567), .B0(n6257), .B1(n3569), .C0(
        top_core_EC_n961), .Y(top_core_EC_n1243) );
  INVX1 U22898 ( .A(top_core_Plain_text[87]), .Y(n4215) );
  AOI22X1 U22899 ( .A0(n3574), .A1(top_core_EC_mix_out_47_), .B0(
        top_core_EC_add_out_r_47_), .B1(n3580), .Y(top_core_EC_n961) );
  OAI221XL U22900 ( .A0(n4200), .A1(top_core_EC_n947), .B0(n6256), .B1(n3569), 
        .C0(top_core_EC_n960), .Y(top_core_EC_n1242) );
  INVX1 U22901 ( .A(top_core_Plain_text[72]), .Y(n4200) );
  AOI22X1 U22902 ( .A0(n3576), .A1(top_core_EC_mix_out_48_), .B0(
        top_core_EC_add_out_r_48_), .B1(top_core_EC_n951), .Y(top_core_EC_n960) );
  OAI221XL U22903 ( .A0(n4201), .A1(top_core_EC_n947), .B0(n6255), .B1(n3569), 
        .C0(top_core_EC_n959), .Y(top_core_EC_n1241) );
  INVX1 U22904 ( .A(top_core_Plain_text[73]), .Y(n4201) );
  AOI22X1 U22905 ( .A0(n3576), .A1(top_core_EC_mix_out_49_), .B0(
        top_core_EC_add_out_r_49_), .B1(top_core_EC_n951), .Y(top_core_EC_n959) );
  OAI221XL U22906 ( .A0(n4202), .A1(top_core_EC_n947), .B0(n6254), .B1(n3569), 
        .C0(top_core_EC_n958), .Y(top_core_EC_n1240) );
  INVX1 U22907 ( .A(top_core_Plain_text[74]), .Y(n4202) );
  AOI22X1 U22908 ( .A0(n3576), .A1(top_core_EC_mix_out_50_), .B0(
        top_core_EC_add_out_r_50_), .B1(top_core_EC_n951), .Y(top_core_EC_n958) );
  OAI221XL U22909 ( .A0(n4203), .A1(top_core_EC_n947), .B0(n6253), .B1(n3569), 
        .C0(top_core_EC_n957), .Y(top_core_EC_n1239) );
  INVX1 U22910 ( .A(top_core_Plain_text[75]), .Y(n4203) );
  AOI22X1 U22911 ( .A0(n3576), .A1(top_core_EC_mix_out_51_), .B0(
        top_core_EC_add_out_r_51_), .B1(top_core_EC_n951), .Y(top_core_EC_n957) );
  OAI221XL U22912 ( .A0(n4204), .A1(n3565), .B0(n6252), .B1(n3569), .C0(
        top_core_EC_n956), .Y(top_core_EC_n1238) );
  INVX1 U22913 ( .A(top_core_Plain_text[76]), .Y(n4204) );
  AOI22X1 U22914 ( .A0(n3576), .A1(top_core_EC_mix_out_52_), .B0(
        top_core_EC_add_out_r_52_), .B1(top_core_EC_n951), .Y(top_core_EC_n956) );
  OAI221XL U22915 ( .A0(n4205), .A1(n3566), .B0(n6251), .B1(n3569), .C0(
        top_core_EC_n955), .Y(top_core_EC_n1237) );
  INVX1 U22916 ( .A(top_core_Plain_text[77]), .Y(n4205) );
  AOI22X1 U22917 ( .A0(n3576), .A1(top_core_EC_mix_out_53_), .B0(
        top_core_EC_add_out_r_53_), .B1(top_core_EC_n951), .Y(top_core_EC_n955) );
  OAI221XL U22918 ( .A0(n4206), .A1(n3567), .B0(n6250), .B1(n3569), .C0(
        top_core_EC_n954), .Y(top_core_EC_n1236) );
  INVX1 U22919 ( .A(top_core_Plain_text[78]), .Y(n4206) );
  AOI22X1 U22920 ( .A0(n3576), .A1(top_core_EC_mix_out_54_), .B0(
        top_core_EC_add_out_r_54_), .B1(top_core_EC_n951), .Y(top_core_EC_n954) );
  OAI221XL U22921 ( .A0(n4207), .A1(n3564), .B0(n6249), .B1(n3569), .C0(
        top_core_EC_n953), .Y(top_core_EC_n1235) );
  INVX1 U22922 ( .A(top_core_Plain_text[79]), .Y(n4207) );
  AOI22X1 U22923 ( .A0(n3576), .A1(top_core_EC_mix_out_55_), .B0(
        top_core_EC_add_out_r_55_), .B1(top_core_EC_n951), .Y(top_core_EC_n953) );
  OAI221XL U22924 ( .A0(n4198), .A1(n3565), .B0(n6248), .B1(n3569), .C0(
        top_core_EC_n952), .Y(top_core_EC_n1234) );
  INVX1 U22925 ( .A(top_core_Plain_text[64]), .Y(n4198) );
  AOI22X1 U22926 ( .A0(n3576), .A1(top_core_EC_mix_out_56_), .B0(
        top_core_EC_add_out_r_56_), .B1(top_core_EC_n951), .Y(top_core_EC_n952) );
  OAI221XL U22927 ( .A0(n4251), .A1(n3564), .B0(n6301), .B1(n3572), .C0(
        top_core_EC_n1005), .Y(top_core_EC_n1287) );
  INVX1 U22928 ( .A(top_core_Plain_text[123]), .Y(n4251) );
  AOI22X1 U22929 ( .A0(top_core_EC_n950), .A1(top_core_EC_mix_out_3_), .B0(
        top_core_EC_add_out_r_3_), .B1(n3578), .Y(top_core_EC_n1005) );
  OAI221XL U22930 ( .A0(n4252), .A1(n3564), .B0(n6300), .B1(n3572), .C0(
        top_core_EC_n1004), .Y(top_core_EC_n1286) );
  INVX1 U22931 ( .A(top_core_Plain_text[124]), .Y(n4252) );
  AOI22X1 U22932 ( .A0(top_core_EC_n950), .A1(top_core_EC_mix_out_4_), .B0(
        top_core_EC_add_out_r_4_), .B1(n3579), .Y(top_core_EC_n1004) );
  OAI221XL U22933 ( .A0(n4253), .A1(n3564), .B0(n6299), .B1(n3572), .C0(
        top_core_EC_n1003), .Y(top_core_EC_n1285) );
  INVX1 U22934 ( .A(top_core_Plain_text[125]), .Y(n4253) );
  AOI22X1 U22935 ( .A0(top_core_EC_n950), .A1(top_core_EC_mix_out_5_), .B0(
        top_core_EC_add_out_r_5_), .B1(n3580), .Y(top_core_EC_n1003) );
  OAI221XL U22936 ( .A0(n4254), .A1(n3564), .B0(n6298), .B1(n3572), .C0(
        top_core_EC_n1002), .Y(top_core_EC_n1284) );
  INVX1 U22937 ( .A(top_core_Plain_text[126]), .Y(n4254) );
  AOI22X1 U22938 ( .A0(top_core_EC_n950), .A1(top_core_EC_mix_out_6_), .B0(
        top_core_EC_add_out_r_6_), .B1(n3578), .Y(top_core_EC_n1002) );
  OAI221XL U22939 ( .A0(n4255), .A1(n3564), .B0(n6297), .B1(n3572), .C0(
        top_core_EC_n1001), .Y(top_core_EC_n1283) );
  INVX1 U22940 ( .A(top_core_Plain_text[127]), .Y(n4255) );
  AOI22X1 U22941 ( .A0(top_core_EC_n950), .A1(top_core_EC_mix_out_7_), .B0(
        top_core_EC_add_out_r_7_), .B1(n3579), .Y(top_core_EC_n1001) );
  OAI221XL U22942 ( .A0(n4240), .A1(n3564), .B0(n6296), .B1(n3572), .C0(
        top_core_EC_n1000), .Y(top_core_EC_n1282) );
  INVX1 U22943 ( .A(top_core_Plain_text[112]), .Y(n4240) );
  AOI22X1 U22944 ( .A0(top_core_EC_n950), .A1(top_core_EC_mix_out_8_), .B0(
        top_core_EC_add_out_r_8_), .B1(n3580), .Y(top_core_EC_n1000) );
  OAI221XL U22945 ( .A0(n4241), .A1(n3564), .B0(n6295), .B1(n3572), .C0(
        top_core_EC_n999), .Y(top_core_EC_n1281) );
  INVX1 U22946 ( .A(top_core_Plain_text[113]), .Y(n4241) );
  AOI22X1 U22947 ( .A0(top_core_EC_n950), .A1(top_core_EC_mix_out_9_), .B0(
        top_core_EC_add_out_r_9_), .B1(n3578), .Y(top_core_EC_n999) );
  OAI221XL U22948 ( .A0(n4242), .A1(n3564), .B0(n6294), .B1(n3572), .C0(
        top_core_EC_n998), .Y(top_core_EC_n1280) );
  INVX1 U22949 ( .A(top_core_Plain_text[114]), .Y(n4242) );
  AOI22X1 U22950 ( .A0(top_core_EC_n950), .A1(top_core_EC_mix_out_10_), .B0(
        top_core_EC_add_out_r_10_), .B1(n3579), .Y(top_core_EC_n998) );
  OAI221XL U22951 ( .A0(n4243), .A1(n3564), .B0(n6293), .B1(n3572), .C0(
        top_core_EC_n997), .Y(top_core_EC_n1279) );
  INVX1 U22952 ( .A(top_core_Plain_text[115]), .Y(n4243) );
  AOI22X1 U22953 ( .A0(top_core_EC_n950), .A1(top_core_EC_mix_out_11_), .B0(
        top_core_EC_add_out_r_11_), .B1(n3580), .Y(top_core_EC_n997) );
  OAI221XL U22954 ( .A0(n4244), .A1(n3565), .B0(n6292), .B1(n3572), .C0(
        top_core_EC_n996), .Y(top_core_EC_n1278) );
  INVX1 U22955 ( .A(top_core_Plain_text[116]), .Y(n4244) );
  AOI22X1 U22956 ( .A0(n3574), .A1(top_core_EC_mix_out_12_), .B0(
        top_core_EC_add_out_r_12_), .B1(n3578), .Y(top_core_EC_n996) );
  OAI221XL U22957 ( .A0(n4245), .A1(n3565), .B0(n6291), .B1(n3572), .C0(
        top_core_EC_n995), .Y(top_core_EC_n1277) );
  INVX1 U22958 ( .A(top_core_Plain_text[117]), .Y(n4245) );
  AOI22X1 U22959 ( .A0(n3574), .A1(top_core_EC_mix_out_13_), .B0(
        top_core_EC_add_out_r_13_), .B1(n3578), .Y(top_core_EC_n995) );
  OAI221XL U22960 ( .A0(n4246), .A1(n3565), .B0(n6290), .B1(n3572), .C0(
        top_core_EC_n994), .Y(top_core_EC_n1276) );
  INVX1 U22961 ( .A(top_core_Plain_text[118]), .Y(n4246) );
  AOI22X1 U22962 ( .A0(n3574), .A1(top_core_EC_mix_out_14_), .B0(
        top_core_EC_add_out_r_14_), .B1(n3578), .Y(top_core_EC_n994) );
  OAI221XL U22963 ( .A0(n4247), .A1(n3565), .B0(n6289), .B1(n3572), .C0(
        top_core_EC_n993), .Y(top_core_EC_n1275) );
  INVX1 U22964 ( .A(top_core_Plain_text[119]), .Y(n4247) );
  AOI22X1 U22965 ( .A0(n3574), .A1(top_core_EC_mix_out_15_), .B0(
        top_core_EC_add_out_r_15_), .B1(n3578), .Y(top_core_EC_n993) );
  OAI221XL U22966 ( .A0(n4232), .A1(n3565), .B0(n6288), .B1(n3572), .C0(
        top_core_EC_n992), .Y(top_core_EC_n1274) );
  INVX1 U22967 ( .A(top_core_Plain_text[104]), .Y(n4232) );
  AOI22X1 U22968 ( .A0(n3574), .A1(top_core_EC_mix_out_16_), .B0(
        top_core_EC_add_out_r_16_), .B1(n3578), .Y(top_core_EC_n992) );
  OAI221XL U22969 ( .A0(n4233), .A1(n3565), .B0(n6287), .B1(n3571), .C0(
        top_core_EC_n991), .Y(top_core_EC_n1273) );
  INVX1 U22970 ( .A(top_core_Plain_text[105]), .Y(n4233) );
  AOI22X1 U22971 ( .A0(n3574), .A1(top_core_EC_mix_out_17_), .B0(
        top_core_EC_add_out_r_17_), .B1(n3578), .Y(top_core_EC_n991) );
  OAI221XL U22972 ( .A0(n4234), .A1(n3565), .B0(n6286), .B1(n3571), .C0(
        top_core_EC_n990), .Y(top_core_EC_n1272) );
  INVX1 U22973 ( .A(top_core_Plain_text[106]), .Y(n4234) );
  AOI22X1 U22974 ( .A0(n3574), .A1(top_core_EC_mix_out_18_), .B0(
        top_core_EC_add_out_r_18_), .B1(n3578), .Y(top_core_EC_n990) );
  OAI221XL U22975 ( .A0(n4235), .A1(n3565), .B0(n6285), .B1(n3571), .C0(
        top_core_EC_n989), .Y(top_core_EC_n1271) );
  INVX1 U22976 ( .A(top_core_Plain_text[107]), .Y(n4235) );
  AOI22X1 U22977 ( .A0(n3574), .A1(top_core_EC_mix_out_19_), .B0(
        top_core_EC_add_out_r_19_), .B1(n3578), .Y(top_core_EC_n989) );
  OAI221XL U22978 ( .A0(n4236), .A1(n3565), .B0(n6284), .B1(n3571), .C0(
        top_core_EC_n988), .Y(top_core_EC_n1270) );
  INVX1 U22979 ( .A(top_core_Plain_text[108]), .Y(n4236) );
  AOI22X1 U22980 ( .A0(n3574), .A1(top_core_EC_mix_out_20_), .B0(
        top_core_EC_add_out_r_20_), .B1(n3578), .Y(top_core_EC_n988) );
  OAI221XL U22981 ( .A0(n4237), .A1(n3565), .B0(n6283), .B1(n3571), .C0(
        top_core_EC_n987), .Y(top_core_EC_n1269) );
  INVX1 U22982 ( .A(top_core_Plain_text[109]), .Y(n4237) );
  AOI22X1 U22983 ( .A0(n3574), .A1(top_core_EC_mix_out_21_), .B0(
        top_core_EC_add_out_r_21_), .B1(n3578), .Y(top_core_EC_n987) );
  OAI221XL U22984 ( .A0(n4238), .A1(n3565), .B0(n6282), .B1(n3571), .C0(
        top_core_EC_n986), .Y(top_core_EC_n1268) );
  INVX1 U22985 ( .A(top_core_Plain_text[110]), .Y(n4238) );
  AOI22X1 U22986 ( .A0(n3574), .A1(top_core_EC_mix_out_22_), .B0(
        top_core_EC_add_out_r_22_), .B1(n3578), .Y(top_core_EC_n986) );
  OAI221XL U22987 ( .A0(n4239), .A1(n3565), .B0(n6281), .B1(n3571), .C0(
        top_core_EC_n985), .Y(top_core_EC_n1267) );
  INVX1 U22988 ( .A(top_core_Plain_text[111]), .Y(n4239) );
  AOI22X1 U22989 ( .A0(n3574), .A1(top_core_EC_mix_out_23_), .B0(
        top_core_EC_add_out_r_23_), .B1(n3578), .Y(top_core_EC_n985) );
  OAI221XL U22990 ( .A0(n4224), .A1(n3566), .B0(n6280), .B1(n3571), .C0(
        top_core_EC_n984), .Y(top_core_EC_n1266) );
  INVX1 U22991 ( .A(top_core_Plain_text[96]), .Y(n4224) );
  AOI22X1 U22992 ( .A0(n3575), .A1(top_core_EC_mix_out_24_), .B0(
        top_core_EC_add_out_r_24_), .B1(n3579), .Y(top_core_EC_n984) );
  OAI221XL U22993 ( .A0(n4225), .A1(n3566), .B0(n6279), .B1(n3571), .C0(
        top_core_EC_n983), .Y(top_core_EC_n1265) );
  INVX1 U22994 ( .A(top_core_Plain_text[97]), .Y(n4225) );
  AOI22X1 U22995 ( .A0(n3575), .A1(top_core_EC_mix_out_25_), .B0(
        top_core_EC_add_out_r_25_), .B1(n3579), .Y(top_core_EC_n983) );
  OAI221XL U22996 ( .A0(n4226), .A1(n3566), .B0(n6278), .B1(n3571), .C0(
        top_core_EC_n982), .Y(top_core_EC_n1264) );
  INVX1 U22997 ( .A(top_core_Plain_text[98]), .Y(n4226) );
  AOI22X1 U22998 ( .A0(n3575), .A1(top_core_EC_mix_out_26_), .B0(
        top_core_EC_add_out_r_26_), .B1(n3579), .Y(top_core_EC_n982) );
  OAI221XL U22999 ( .A0(n4227), .A1(n3566), .B0(n6277), .B1(n3571), .C0(
        top_core_EC_n981), .Y(top_core_EC_n1263) );
  INVX1 U23000 ( .A(top_core_Plain_text[99]), .Y(n4227) );
  AOI22X1 U23001 ( .A0(n3575), .A1(top_core_EC_mix_out_27_), .B0(
        top_core_EC_add_out_r_27_), .B1(n3579), .Y(top_core_EC_n981) );
  OAI221XL U23002 ( .A0(n4228), .A1(n3566), .B0(n6276), .B1(n3571), .C0(
        top_core_EC_n980), .Y(top_core_EC_n1262) );
  INVX1 U23003 ( .A(top_core_Plain_text[100]), .Y(n4228) );
  AOI22X1 U23004 ( .A0(n3575), .A1(top_core_EC_mix_out_28_), .B0(
        top_core_EC_add_out_r_28_), .B1(n3579), .Y(top_core_EC_n980) );
  OAI221XL U23005 ( .A0(n4229), .A1(n3566), .B0(n6275), .B1(n3571), .C0(
        top_core_EC_n979), .Y(top_core_EC_n1261) );
  INVX1 U23006 ( .A(top_core_Plain_text[101]), .Y(n4229) );
  AOI22X1 U23007 ( .A0(n3575), .A1(top_core_EC_mix_out_29_), .B0(
        top_core_EC_add_out_r_29_), .B1(n3579), .Y(top_core_EC_n979) );
  OAI221XL U23008 ( .A0(n4230), .A1(n3566), .B0(n6274), .B1(n3570), .C0(
        top_core_EC_n978), .Y(top_core_EC_n1260) );
  INVX1 U23009 ( .A(top_core_Plain_text[102]), .Y(n4230) );
  AOI22X1 U23010 ( .A0(n3575), .A1(top_core_EC_mix_out_30_), .B0(
        top_core_EC_add_out_r_30_), .B1(n3579), .Y(top_core_EC_n978) );
  OAI221XL U23011 ( .A0(n4231), .A1(n3566), .B0(n6273), .B1(n3570), .C0(
        top_core_EC_n977), .Y(top_core_EC_n1259) );
  INVX1 U23012 ( .A(top_core_Plain_text[103]), .Y(n4231) );
  AOI22X1 U23013 ( .A0(n3575), .A1(top_core_EC_mix_out_31_), .B0(
        top_core_EC_add_out_r_31_), .B1(n3579), .Y(top_core_EC_n977) );
  OAI221XL U23014 ( .A0(n4216), .A1(n3566), .B0(n6272), .B1(n3570), .C0(
        top_core_EC_n976), .Y(top_core_EC_n1258) );
  INVX1 U23015 ( .A(top_core_Plain_text[88]), .Y(n4216) );
  AOI22X1 U23016 ( .A0(n3575), .A1(top_core_EC_mix_out_32_), .B0(
        top_core_EC_add_out_r_32_), .B1(n3579), .Y(top_core_EC_n976) );
  OAI221XL U23017 ( .A0(n4217), .A1(n3566), .B0(n6271), .B1(n3570), .C0(
        top_core_EC_n975), .Y(top_core_EC_n1257) );
  INVX1 U23018 ( .A(top_core_Plain_text[89]), .Y(n4217) );
  AOI22X1 U23019 ( .A0(n3575), .A1(top_core_EC_mix_out_33_), .B0(
        top_core_EC_add_out_r_33_), .B1(n3579), .Y(top_core_EC_n975) );
  OAI221XL U23020 ( .A0(n4218), .A1(n3566), .B0(n6270), .B1(n3570), .C0(
        top_core_EC_n974), .Y(top_core_EC_n1256) );
  INVX1 U23021 ( .A(top_core_Plain_text[90]), .Y(n4218) );
  AOI22X1 U23022 ( .A0(n3575), .A1(top_core_EC_mix_out_34_), .B0(
        top_core_EC_add_out_r_34_), .B1(n3579), .Y(top_core_EC_n974) );
  OAI221XL U23023 ( .A0(n4219), .A1(n3566), .B0(n6269), .B1(n3570), .C0(
        top_core_EC_n973), .Y(top_core_EC_n1255) );
  INVX1 U23024 ( .A(top_core_Plain_text[91]), .Y(n4219) );
  AOI22X1 U23025 ( .A0(n3575), .A1(top_core_EC_mix_out_35_), .B0(
        top_core_EC_add_out_r_35_), .B1(n3579), .Y(top_core_EC_n973) );
  OAI221XL U23026 ( .A0(n4220), .A1(n3567), .B0(n6268), .B1(n3570), .C0(
        top_core_EC_n972), .Y(top_core_EC_n1254) );
  INVX1 U23027 ( .A(top_core_Plain_text[92]), .Y(n4220) );
  AOI22X1 U23028 ( .A0(n3575), .A1(top_core_EC_mix_out_36_), .B0(
        top_core_EC_add_out_r_36_), .B1(n3580), .Y(top_core_EC_n972) );
  OAI221XL U23029 ( .A0(n4221), .A1(n3567), .B0(n6267), .B1(n3570), .C0(
        top_core_EC_n971), .Y(top_core_EC_n1253) );
  INVX1 U23030 ( .A(top_core_Plain_text[93]), .Y(n4221) );
  AOI22X1 U23031 ( .A0(n3576), .A1(top_core_EC_mix_out_37_), .B0(
        top_core_EC_add_out_r_37_), .B1(n3580), .Y(top_core_EC_n971) );
  OAI221XL U23032 ( .A0(n4222), .A1(n3567), .B0(n6266), .B1(n3570), .C0(
        top_core_EC_n970), .Y(top_core_EC_n1252) );
  INVX1 U23033 ( .A(top_core_Plain_text[94]), .Y(n4222) );
  AOI22X1 U23034 ( .A0(n3574), .A1(top_core_EC_mix_out_38_), .B0(
        top_core_EC_add_out_r_38_), .B1(n3580), .Y(top_core_EC_n970) );
  OAI221XL U23035 ( .A0(n4223), .A1(n3567), .B0(n6265), .B1(n3570), .C0(
        top_core_EC_n969), .Y(top_core_EC_n1251) );
  INVX1 U23036 ( .A(top_core_Plain_text[95]), .Y(n4223) );
  AOI22X1 U23037 ( .A0(n3575), .A1(top_core_EC_mix_out_39_), .B0(
        top_core_EC_add_out_r_39_), .B1(n3580), .Y(top_core_EC_n969) );
  OAI221XL U23038 ( .A0(n4208), .A1(n3567), .B0(n6264), .B1(n3570), .C0(
        top_core_EC_n968), .Y(top_core_EC_n1250) );
  INVX1 U23039 ( .A(top_core_Plain_text[80]), .Y(n4208) );
  AOI22X1 U23040 ( .A0(n3576), .A1(top_core_EC_mix_out_40_), .B0(
        top_core_EC_add_out_r_40_), .B1(n3580), .Y(top_core_EC_n968) );
  OAI221XL U23041 ( .A0(n4209), .A1(n3567), .B0(n6263), .B1(n3570), .C0(
        top_core_EC_n967), .Y(top_core_EC_n1249) );
  INVX1 U23042 ( .A(top_core_Plain_text[81]), .Y(n4209) );
  AOI22X1 U23043 ( .A0(n3574), .A1(top_core_EC_mix_out_41_), .B0(
        top_core_EC_add_out_r_41_), .B1(n3580), .Y(top_core_EC_n967) );
  OAI221XL U23044 ( .A0(n4210), .A1(n3567), .B0(n6262), .B1(n3570), .C0(
        top_core_EC_n966), .Y(top_core_EC_n1248) );
  INVX1 U23045 ( .A(top_core_Plain_text[82]), .Y(n4210) );
  AOI22X1 U23046 ( .A0(n3575), .A1(top_core_EC_mix_out_42_), .B0(
        top_core_EC_add_out_r_42_), .B1(n3580), .Y(top_core_EC_n966) );
  OAI221XL U23047 ( .A0(n4211), .A1(n3567), .B0(n6261), .B1(n3570), .C0(
        top_core_EC_n965), .Y(top_core_EC_n1247) );
  INVX1 U23048 ( .A(top_core_Plain_text[83]), .Y(n4211) );
  AOI22X1 U23049 ( .A0(n3576), .A1(top_core_EC_mix_out_43_), .B0(
        top_core_EC_add_out_r_43_), .B1(n3580), .Y(top_core_EC_n965) );
  OAI221XL U23050 ( .A0(n4199), .A1(n3566), .B0(n6247), .B1(n3571), .C0(
        top_core_EC_n949), .Y(top_core_EC_n1233) );
  INVX1 U23051 ( .A(top_core_Plain_text[65]), .Y(n4199) );
  AOI22X1 U23052 ( .A0(n3576), .A1(top_core_EC_mix_out_57_), .B0(
        top_core_EC_add_out_r_57_), .B1(top_core_EC_n951), .Y(top_core_EC_n949) );
  OAI221XL U23053 ( .A0(n4947), .A1(n3544), .B0(n3549), .B1(n192), .C0(
        top_core_EC_n942), .Y(top_core_EC_n1232) );
  AOI22X1 U23054 ( .A0(n3554), .A1(top_core_Plain_text[66]), .B0(
        top_core_EC_round_result_r_58_), .B1(n3561), .Y(top_core_EC_n942) );
  OAI221XL U23055 ( .A0(n4942), .A1(n3544), .B0(n3549), .B1(n193), .C0(
        top_core_EC_n941), .Y(top_core_EC_n1231) );
  AOI22X1 U23056 ( .A0(n3554), .A1(top_core_Plain_text[67]), .B0(
        top_core_EC_round_result_r_59_), .B1(n3563), .Y(top_core_EC_n941) );
  OAI221XL U23057 ( .A0(n4952), .A1(n3544), .B0(n3549), .B1(n128), .C0(
        top_core_EC_n940), .Y(top_core_EC_n1230) );
  AOI22X1 U23058 ( .A0(n3554), .A1(top_core_Plain_text[68]), .B0(
        top_core_EC_round_result_r_60_), .B1(n3562), .Y(top_core_EC_n940) );
  OAI221XL U23059 ( .A0(n4936), .A1(n3544), .B0(n3549), .B1(n194), .C0(
        top_core_EC_n939), .Y(top_core_EC_n1229) );
  AOI22X1 U23060 ( .A0(n3554), .A1(top_core_Plain_text[69]), .B0(
        top_core_EC_round_result_r_61_), .B1(n3560), .Y(top_core_EC_n939) );
  OAI221XL U23061 ( .A0(n4933), .A1(n3544), .B0(n3549), .B1(n195), .C0(
        top_core_EC_n938), .Y(top_core_EC_n1228) );
  AOI22X1 U23062 ( .A0(n3554), .A1(top_core_Plain_text[70]), .B0(
        top_core_EC_round_result_r_62_), .B1(n3559), .Y(top_core_EC_n938) );
  OAI221XL U23063 ( .A0(n4925), .A1(n3544), .B0(n3549), .B1(n196), .C0(
        top_core_EC_n937), .Y(top_core_EC_n1227) );
  AOI22X1 U23064 ( .A0(n3554), .A1(top_core_Plain_text[71]), .B0(
        top_core_EC_round_result_r_63_), .B1(n3561), .Y(top_core_EC_n937) );
  OAI221XL U23065 ( .A0(n4806), .A1(n3544), .B0(n3549), .B1(n197), .C0(
        top_core_EC_n936), .Y(top_core_EC_n1226) );
  AOI22X1 U23066 ( .A0(n3554), .A1(top_core_Plain_text[56]), .B0(
        top_core_EC_round_result_r_64_), .B1(n3563), .Y(top_core_EC_n936) );
  OAI221XL U23067 ( .A0(n4804), .A1(n3544), .B0(n3549), .B1(n198), .C0(
        top_core_EC_n935), .Y(top_core_EC_n1225) );
  AOI22X1 U23068 ( .A0(n3554), .A1(top_core_Plain_text[57]), .B0(
        top_core_EC_round_result_r_65_), .B1(n3562), .Y(top_core_EC_n935) );
  OAI221XL U23069 ( .A0(n4798), .A1(n3544), .B0(n3549), .B1(n199), .C0(
        top_core_EC_n934), .Y(top_core_EC_n1224) );
  AOI22X1 U23070 ( .A0(n3554), .A1(top_core_Plain_text[58]), .B0(
        top_core_EC_round_result_r_66_), .B1(n3560), .Y(top_core_EC_n934) );
  OAI221XL U23071 ( .A0(n4793), .A1(n3544), .B0(n3549), .B1(n200), .C0(
        top_core_EC_n933), .Y(top_core_EC_n1223) );
  AOI22X1 U23072 ( .A0(n3554), .A1(top_core_Plain_text[59]), .B0(
        top_core_EC_round_result_r_67_), .B1(n3559), .Y(top_core_EC_n933) );
  OAI221XL U23073 ( .A0(n4803), .A1(n3544), .B0(n3549), .B1(n152), .C0(
        top_core_EC_n932), .Y(top_core_EC_n1222) );
  AOI22X1 U23074 ( .A0(n3554), .A1(top_core_Plain_text[60]), .B0(
        top_core_EC_round_result_r_68_), .B1(n3563), .Y(top_core_EC_n932) );
  OAI221XL U23075 ( .A0(n4787), .A1(n3544), .B0(n3549), .B1(n127), .C0(
        top_core_EC_n931), .Y(top_core_EC_n1221) );
  AOI22X1 U23076 ( .A0(n3554), .A1(top_core_Plain_text[61]), .B0(
        top_core_EC_round_result_r_69_), .B1(n3563), .Y(top_core_EC_n931) );
  OAI221XL U23077 ( .A0(n4782), .A1(n3545), .B0(n3549), .B1(n126), .C0(
        top_core_EC_n930), .Y(top_core_EC_n1220) );
  AOI22X1 U23078 ( .A0(n3555), .A1(top_core_Plain_text[62]), .B0(
        top_core_EC_round_result_r_70_), .B1(n3563), .Y(top_core_EC_n930) );
  OAI221XL U23079 ( .A0(n4775), .A1(n3545), .B0(n3552), .B1(n153), .C0(
        top_core_EC_n929), .Y(top_core_EC_n1219) );
  AOI22X1 U23080 ( .A0(n3555), .A1(top_core_Plain_text[63]), .B0(
        top_core_EC_round_result_r_71_), .B1(n3563), .Y(top_core_EC_n929) );
  OAI221XL U23081 ( .A0(n4805), .A1(n3545), .B0(n3550), .B1(n201), .C0(
        top_core_EC_n928), .Y(top_core_EC_n1218) );
  AOI22X1 U23082 ( .A0(n3555), .A1(top_core_Plain_text[48]), .B0(
        top_core_EC_round_result_r_72_), .B1(n3563), .Y(top_core_EC_n928) );
  OAI221XL U23083 ( .A0(n4797), .A1(n3545), .B0(n3551), .B1(n154), .C0(
        top_core_EC_n927), .Y(top_core_EC_n1217) );
  AOI22X1 U23084 ( .A0(n3555), .A1(top_core_Plain_text[49]), .B0(
        top_core_EC_round_result_r_73_), .B1(n3563), .Y(top_core_EC_n927) );
  OAI221XL U23085 ( .A0(n4795), .A1(n3545), .B0(n3549), .B1(n202), .C0(
        top_core_EC_n926), .Y(top_core_EC_n1216) );
  AOI22X1 U23086 ( .A0(n3555), .A1(top_core_Plain_text[50]), .B0(
        top_core_EC_round_result_r_74_), .B1(n3563), .Y(top_core_EC_n926) );
  OAI221XL U23087 ( .A0(n4794), .A1(n3545), .B0(n3552), .B1(n203), .C0(
        top_core_EC_n925), .Y(top_core_EC_n1215) );
  AOI22X1 U23088 ( .A0(n3555), .A1(top_core_Plain_text[51]), .B0(
        top_core_EC_round_result_r_75_), .B1(n3563), .Y(top_core_EC_n925) );
  OAI221XL U23089 ( .A0(n4786), .A1(n3545), .B0(n3550), .B1(n155), .C0(
        top_core_EC_n924), .Y(top_core_EC_n1214) );
  AOI22X1 U23090 ( .A0(n3555), .A1(top_core_Plain_text[52]), .B0(
        top_core_EC_round_result_r_76_), .B1(n3563), .Y(top_core_EC_n924) );
  OAI221XL U23091 ( .A0(n4780), .A1(n3545), .B0(n3551), .B1(n204), .C0(
        top_core_EC_n923), .Y(top_core_EC_n1213) );
  AOI22X1 U23092 ( .A0(n3555), .A1(top_core_Plain_text[53]), .B0(
        top_core_EC_round_result_r_77_), .B1(n3563), .Y(top_core_EC_n923) );
  OAI221XL U23093 ( .A0(n4783), .A1(n3545), .B0(n3549), .B1(n205), .C0(
        top_core_EC_n922), .Y(top_core_EC_n1212) );
  AOI22X1 U23094 ( .A0(n3555), .A1(top_core_Plain_text[54]), .B0(
        top_core_EC_round_result_r_78_), .B1(n3563), .Y(top_core_EC_n922) );
  OAI221XL U23095 ( .A0(n4776), .A1(n3545), .B0(n3552), .B1(n206), .C0(
        top_core_EC_n921), .Y(top_core_EC_n1211) );
  AOI22X1 U23096 ( .A0(n3555), .A1(top_core_Plain_text[55]), .B0(
        top_core_EC_round_result_r_79_), .B1(n3563), .Y(top_core_EC_n921) );
  OAI221XL U23097 ( .A0(n4800), .A1(n3545), .B0(n3550), .B1(n207), .C0(
        top_core_EC_n920), .Y(top_core_EC_n1210) );
  AOI22X1 U23098 ( .A0(n3555), .A1(top_core_Plain_text[40]), .B0(
        top_core_EC_round_result_r_80_), .B1(n3562), .Y(top_core_EC_n920) );
  OAI221XL U23099 ( .A0(n4792), .A1(n3545), .B0(n3551), .B1(n208), .C0(
        top_core_EC_n919), .Y(top_core_EC_n1209) );
  AOI22X1 U23100 ( .A0(n3555), .A1(top_core_Plain_text[41]), .B0(
        top_core_EC_round_result_r_81_), .B1(n3562), .Y(top_core_EC_n919) );
  OAI221XL U23101 ( .A0(n4799), .A1(n3546), .B0(n3550), .B1(n209), .C0(
        top_core_EC_n918), .Y(top_core_EC_n1208) );
  AOI22X1 U23102 ( .A0(n3556), .A1(top_core_Plain_text[42]), .B0(
        top_core_EC_round_result_r_82_), .B1(n3562), .Y(top_core_EC_n918) );
  OAI221XL U23103 ( .A0(n4789), .A1(n3546), .B0(n3550), .B1(n210), .C0(
        top_core_EC_n917), .Y(top_core_EC_n1207) );
  AOI22X1 U23104 ( .A0(n3556), .A1(top_core_Plain_text[43]), .B0(
        top_core_EC_round_result_r_83_), .B1(n3562), .Y(top_core_EC_n917) );
  OAI221XL U23105 ( .A0(n4779), .A1(n3546), .B0(n3550), .B1(n156), .C0(
        top_core_EC_n916), .Y(top_core_EC_n1206) );
  AOI22X1 U23106 ( .A0(n3556), .A1(top_core_Plain_text[44]), .B0(
        top_core_EC_round_result_r_84_), .B1(n3562), .Y(top_core_EC_n916) );
  OAI221XL U23107 ( .A0(n4788), .A1(n3546), .B0(n3550), .B1(n125), .C0(
        top_core_EC_n915), .Y(top_core_EC_n1205) );
  AOI22X1 U23108 ( .A0(n3556), .A1(top_core_Plain_text[45]), .B0(
        top_core_EC_round_result_r_85_), .B1(n3562), .Y(top_core_EC_n915) );
  OAI221XL U23109 ( .A0(n4784), .A1(n3546), .B0(n3550), .B1(n124), .C0(
        top_core_EC_n914), .Y(top_core_EC_n1204) );
  AOI22X1 U23110 ( .A0(n3556), .A1(top_core_Plain_text[46]), .B0(
        top_core_EC_round_result_r_86_), .B1(n3562), .Y(top_core_EC_n914) );
  OAI221XL U23111 ( .A0(n4777), .A1(n3546), .B0(n3550), .B1(n123), .C0(
        top_core_EC_n913), .Y(top_core_EC_n1203) );
  AOI22X1 U23112 ( .A0(n3556), .A1(top_core_Plain_text[47]), .B0(
        top_core_EC_round_result_r_87_), .B1(n3562), .Y(top_core_EC_n913) );
  OAI221XL U23113 ( .A0(n4801), .A1(n3546), .B0(n3550), .B1(n211), .C0(
        top_core_EC_n912), .Y(top_core_EC_n1202) );
  AOI22X1 U23114 ( .A0(n3556), .A1(top_core_Plain_text[32]), .B0(
        top_core_EC_round_result_r_88_), .B1(n3562), .Y(top_core_EC_n912) );
  OAI221XL U23115 ( .A0(n4791), .A1(n3546), .B0(n3550), .B1(n157), .C0(
        top_core_EC_n911), .Y(top_core_EC_n1201) );
  AOI22X1 U23116 ( .A0(n3556), .A1(top_core_Plain_text[33]), .B0(
        top_core_EC_round_result_r_89_), .B1(n3562), .Y(top_core_EC_n911) );
  OAI221XL U23117 ( .A0(n4796), .A1(n3546), .B0(n3550), .B1(n212), .C0(
        top_core_EC_n910), .Y(top_core_EC_n1200) );
  AOI22X1 U23118 ( .A0(n3556), .A1(top_core_Plain_text[34]), .B0(
        top_core_EC_round_result_r_90_), .B1(n3562), .Y(top_core_EC_n910) );
  OAI221XL U23119 ( .A0(n4790), .A1(n3546), .B0(n3550), .B1(n213), .C0(
        top_core_EC_n909), .Y(top_core_EC_n1199) );
  AOI22X1 U23120 ( .A0(n3556), .A1(top_core_Plain_text[35]), .B0(
        top_core_EC_round_result_r_91_), .B1(n3562), .Y(top_core_EC_n909) );
  OAI221XL U23121 ( .A0(n4778), .A1(n3546), .B0(n3550), .B1(n122), .C0(
        top_core_EC_n908), .Y(top_core_EC_n1198) );
  AOI22X1 U23122 ( .A0(n3556), .A1(top_core_Plain_text[36]), .B0(
        top_core_EC_round_result_r_92_), .B1(n3561), .Y(top_core_EC_n908) );
  OAI221XL U23123 ( .A0(n4781), .A1(n3546), .B0(n3550), .B1(n214), .C0(
        top_core_EC_n907), .Y(top_core_EC_n1197) );
  AOI22X1 U23124 ( .A0(n3556), .A1(top_core_Plain_text[37]), .B0(
        top_core_EC_round_result_r_93_), .B1(n3561), .Y(top_core_EC_n907) );
  OAI221XL U23125 ( .A0(n4785), .A1(n3546), .B0(n3551), .B1(n215), .C0(
        top_core_EC_n906), .Y(top_core_EC_n1196) );
  AOI22X1 U23126 ( .A0(n3557), .A1(top_core_Plain_text[38]), .B0(
        top_core_EC_round_result_r_94_), .B1(n3561), .Y(top_core_EC_n906) );
  OAI221XL U23127 ( .A0(n4802), .A1(n3547), .B0(n3551), .B1(n216), .C0(
        top_core_EC_n905), .Y(top_core_EC_n1195) );
  AOI22X1 U23128 ( .A0(n3554), .A1(top_core_Plain_text[39]), .B0(
        top_core_EC_round_result_r_95_), .B1(n3561), .Y(top_core_EC_n905) );
  OAI221XL U23129 ( .A0(n5149), .A1(n3544), .B0(n3551), .B1(n217), .C0(
        top_core_EC_n904), .Y(top_core_EC_n1194) );
  AOI22X1 U23130 ( .A0(n3555), .A1(top_core_Plain_text[24]), .B0(
        top_core_EC_round_result_r_96_), .B1(n3561), .Y(top_core_EC_n904) );
  OAI221XL U23131 ( .A0(n5140), .A1(n3545), .B0(n3551), .B1(n218), .C0(
        top_core_EC_n903), .Y(top_core_EC_n1193) );
  AOI22X1 U23132 ( .A0(n3556), .A1(top_core_Plain_text[25]), .B0(
        top_core_EC_round_result_r_97_), .B1(n3561), .Y(top_core_EC_n903) );
  OAI221XL U23133 ( .A0(n5144), .A1(n3546), .B0(n3551), .B1(n219), .C0(
        top_core_EC_n902), .Y(top_core_EC_n1192) );
  AOI22X1 U23134 ( .A0(n3557), .A1(top_core_Plain_text[26]), .B0(
        top_core_EC_round_result_r_98_), .B1(n3561), .Y(top_core_EC_n902) );
  OAI221XL U23135 ( .A0(n5138), .A1(n3547), .B0(n3551), .B1(n220), .C0(
        top_core_EC_n901), .Y(top_core_EC_n1191) );
  AOI22X1 U23136 ( .A0(n3554), .A1(top_core_Plain_text[27]), .B0(
        top_core_EC_round_result_r_99_), .B1(n3561), .Y(top_core_EC_n901) );
  OAI221XL U23137 ( .A0(n5126), .A1(n3544), .B0(n3551), .B1(n158), .C0(
        top_core_EC_n900), .Y(top_core_EC_n1190) );
  AOI22X1 U23138 ( .A0(n3555), .A1(top_core_Plain_text[28]), .B0(
        top_core_EC_round_result_r_100_), .B1(n3561), .Y(top_core_EC_n900) );
  OAI221XL U23139 ( .A0(n5128), .A1(n3545), .B0(n3551), .B1(n134), .C0(
        top_core_EC_n899), .Y(top_core_EC_n1189) );
  AOI22X1 U23140 ( .A0(n3556), .A1(top_core_Plain_text[29]), .B0(
        top_core_EC_round_result_r_101_), .B1(n3561), .Y(top_core_EC_n899) );
  OAI221XL U23141 ( .A0(n5130), .A1(n3546), .B0(n3551), .B1(n133), .C0(
        top_core_EC_n898), .Y(top_core_EC_n1188) );
  AOI22X1 U23142 ( .A0(n3557), .A1(top_core_Plain_text[30]), .B0(
        top_core_EC_round_result_r_102_), .B1(n3561), .Y(top_core_EC_n898) );
  OAI221XL U23143 ( .A0(n5150), .A1(n3547), .B0(n3551), .B1(n159), .C0(
        top_core_EC_n897), .Y(top_core_EC_n1187) );
  AOI22X1 U23144 ( .A0(n3554), .A1(top_core_Plain_text[31]), .B0(
        top_core_EC_round_result_r_103_), .B1(n3561), .Y(top_core_EC_n897) );
  OAI221XL U23145 ( .A0(n5154), .A1(n3544), .B0(n3551), .B1(n221), .C0(
        top_core_EC_n896), .Y(top_core_EC_n1186) );
  AOI22X1 U23146 ( .A0(n3555), .A1(top_core_Plain_text[16]), .B0(
        top_core_EC_round_result_r_104_), .B1(n3560), .Y(top_core_EC_n896) );
  OAI221XL U23147 ( .A0(n5152), .A1(n3545), .B0(n3551), .B1(n160), .C0(
        top_core_EC_n895), .Y(top_core_EC_n1185) );
  AOI22X1 U23148 ( .A0(n3556), .A1(top_core_Plain_text[17]), .B0(
        top_core_EC_round_result_r_105_), .B1(n3560), .Y(top_core_EC_n895) );
  OAI221XL U23149 ( .A0(n5146), .A1(n3547), .B0(top_core_EC_n870), .B1(n222), 
        .C0(top_core_EC_n894), .Y(top_core_EC_n1184) );
  AOI22X1 U23150 ( .A0(n3557), .A1(top_core_Plain_text[18]), .B0(
        top_core_EC_round_result_r_106_), .B1(n3560), .Y(top_core_EC_n894) );
  OAI221XL U23151 ( .A0(n5141), .A1(n3547), .B0(top_core_EC_n870), .B1(n223), 
        .C0(top_core_EC_n893), .Y(top_core_EC_n1183) );
  AOI22X1 U23152 ( .A0(n3557), .A1(top_core_Plain_text[19]), .B0(
        top_core_EC_round_result_r_107_), .B1(n3560), .Y(top_core_EC_n893) );
  OAI221XL U23153 ( .A0(n5151), .A1(n3547), .B0(top_core_EC_n870), .B1(n161), 
        .C0(top_core_EC_n892), .Y(top_core_EC_n1182) );
  AOI22X1 U23154 ( .A0(n3557), .A1(top_core_Plain_text[20]), .B0(
        top_core_EC_round_result_r_108_), .B1(n3560), .Y(top_core_EC_n892) );
  OAI221XL U23155 ( .A0(n5135), .A1(n3547), .B0(n3552), .B1(n224), .C0(
        top_core_EC_n891), .Y(top_core_EC_n1181) );
  AOI22X1 U23156 ( .A0(n3557), .A1(top_core_Plain_text[21]), .B0(
        top_core_EC_round_result_r_109_), .B1(n3560), .Y(top_core_EC_n891) );
  OAI221XL U23157 ( .A0(n5131), .A1(n3547), .B0(n3552), .B1(n225), .C0(
        top_core_EC_n890), .Y(top_core_EC_n1180) );
  AOI22X1 U23158 ( .A0(n3557), .A1(top_core_Plain_text[22]), .B0(
        top_core_EC_round_result_r_110_), .B1(n3560), .Y(top_core_EC_n890) );
  OAI221XL U23159 ( .A0(n5123), .A1(n3547), .B0(n3552), .B1(n226), .C0(
        top_core_EC_n889), .Y(top_core_EC_n1179) );
  AOI22X1 U23160 ( .A0(n3557), .A1(top_core_Plain_text[23]), .B0(
        top_core_EC_round_result_r_111_), .B1(n3560), .Y(top_core_EC_n889) );
  OAI221XL U23161 ( .A0(n5153), .A1(n3547), .B0(n3550), .B1(n227), .C0(
        top_core_EC_n888), .Y(top_core_EC_n1178) );
  AOI22X1 U23162 ( .A0(n3557), .A1(top_core_Plain_text[8]), .B0(
        top_core_EC_round_result_r_112_), .B1(n3560), .Y(top_core_EC_n888) );
  OAI221XL U23163 ( .A0(n5145), .A1(n3547), .B0(n3551), .B1(n228), .C0(
        top_core_EC_n887), .Y(top_core_EC_n1177) );
  AOI22X1 U23164 ( .A0(n3557), .A1(top_core_Plain_text[9]), .B0(
        top_core_EC_round_result_r_113_), .B1(n3560), .Y(top_core_EC_n887) );
  OAI221XL U23165 ( .A0(n5143), .A1(n3547), .B0(n3549), .B1(n229), .C0(
        top_core_EC_n886), .Y(top_core_EC_n1176) );
  AOI22X1 U23166 ( .A0(n3557), .A1(top_core_Plain_text[10]), .B0(
        top_core_EC_round_result_r_114_), .B1(n3560), .Y(top_core_EC_n886) );
  OAI221XL U23167 ( .A0(n5142), .A1(n3547), .B0(n3551), .B1(n230), .C0(
        top_core_EC_n885), .Y(top_core_EC_n1175) );
  AOI22X1 U23168 ( .A0(n3557), .A1(top_core_Plain_text[11]), .B0(
        top_core_EC_round_result_r_115_), .B1(n3560), .Y(top_core_EC_n885) );
  OAI221XL U23169 ( .A0(n5134), .A1(n3547), .B0(n3552), .B1(n162), .C0(
        top_core_EC_n884), .Y(top_core_EC_n1174) );
  AOI22X1 U23170 ( .A0(n3557), .A1(top_core_Plain_text[12]), .B0(
        top_core_EC_round_result_r_116_), .B1(n3559), .Y(top_core_EC_n884) );
  OAI221XL U23171 ( .A0(n5129), .A1(n3547), .B0(n3550), .B1(n132), .C0(
        top_core_EC_n883), .Y(top_core_EC_n1173) );
  AOI22X1 U23172 ( .A0(n3557), .A1(top_core_Plain_text[13]), .B0(
        top_core_EC_round_result_r_117_), .B1(n3559), .Y(top_core_EC_n883) );
  OAI221XL U23173 ( .A0(n5132), .A1(top_core_EC_n869), .B0(n3552), .B1(n131), 
        .C0(top_core_EC_n882), .Y(top_core_EC_n1172) );
  AOI22X1 U23174 ( .A0(top_core_EC_n872), .A1(top_core_Plain_text[14]), .B0(
        top_core_EC_round_result_r_118_), .B1(n3559), .Y(top_core_EC_n882) );
  OAI221XL U23175 ( .A0(n5125), .A1(top_core_EC_n869), .B0(n3552), .B1(n130), 
        .C0(top_core_EC_n881), .Y(top_core_EC_n1171) );
  AOI22X1 U23176 ( .A0(top_core_EC_n872), .A1(top_core_Plain_text[15]), .B0(
        top_core_EC_round_result_r_119_), .B1(n3559), .Y(top_core_EC_n881) );
  OAI221XL U23177 ( .A0(n5148), .A1(top_core_EC_n869), .B0(n3552), .B1(n231), 
        .C0(top_core_EC_n880), .Y(top_core_EC_n1170) );
  AOI22X1 U23178 ( .A0(n3557), .A1(top_core_Plain_text[0]), .B0(
        top_core_EC_round_result_r_120_), .B1(n3559), .Y(top_core_EC_n880) );
  OAI221XL U23179 ( .A0(n5139), .A1(n3547), .B0(n3552), .B1(n163), .C0(
        top_core_EC_n879), .Y(top_core_EC_n1169) );
  AOI22X1 U23180 ( .A0(n3554), .A1(top_core_Plain_text[1]), .B0(
        top_core_EC_round_result_r_121_), .B1(n3559), .Y(top_core_EC_n879) );
  OAI221XL U23181 ( .A0(n5147), .A1(n3544), .B0(n3552), .B1(n232), .C0(
        top_core_EC_n878), .Y(top_core_EC_n1168) );
  AOI22X1 U23182 ( .A0(n3555), .A1(top_core_Plain_text[2]), .B0(
        top_core_EC_round_result_r_122_), .B1(n3559), .Y(top_core_EC_n878) );
  OAI221XL U23183 ( .A0(n5137), .A1(n3545), .B0(n3552), .B1(n233), .C0(
        top_core_EC_n877), .Y(top_core_EC_n1167) );
  AOI22X1 U23184 ( .A0(n3556), .A1(top_core_Plain_text[3]), .B0(
        top_core_EC_round_result_r_123_), .B1(n3559), .Y(top_core_EC_n877) );
  OAI221XL U23185 ( .A0(n5127), .A1(n3546), .B0(n3552), .B1(n129), .C0(
        top_core_EC_n876), .Y(top_core_EC_n1166) );
  AOI22X1 U23186 ( .A0(n3556), .A1(top_core_Plain_text[4]), .B0(
        top_core_EC_round_result_r_124_), .B1(n3559), .Y(top_core_EC_n876) );
  OAI221XL U23187 ( .A0(n5136), .A1(n3545), .B0(n3552), .B1(n234), .C0(
        top_core_EC_n875), .Y(top_core_EC_n1165) );
  AOI22X1 U23188 ( .A0(n3557), .A1(top_core_Plain_text[5]), .B0(
        top_core_EC_round_result_r_125_), .B1(n3559), .Y(top_core_EC_n875) );
  OAI221XL U23189 ( .A0(n5133), .A1(n3547), .B0(n3552), .B1(n235), .C0(
        top_core_EC_n874), .Y(top_core_EC_n1164) );
  AOI22X1 U23190 ( .A0(n3554), .A1(top_core_Plain_text[6]), .B0(
        top_core_EC_round_result_r_126_), .B1(n3559), .Y(top_core_EC_n874) );
  OAI221XL U23191 ( .A0(n5124), .A1(n3544), .B0(n3552), .B1(n236), .C0(
        top_core_EC_n871), .Y(top_core_EC_n1163) );
  AOI22X1 U23192 ( .A0(n3555), .A1(top_core_Plain_text[7]), .B0(
        top_core_EC_round_result_r_127_), .B1(n3559), .Y(top_core_EC_n871) );
  OAI221XL U23193 ( .A0(n1500), .A1(top_core_KE_n2709), .B0(n7002), .B1(n151), 
        .C0(top_core_KE_n2710), .Y(top_core_KE_n4924) );
  XNOR2X1 U23194 ( .A(top_core_KE_rcon_reg_2_), .B(top_core_KE_rcon_reg_7_), 
        .Y(top_core_KE_n2709) );
  OAI221XL U23195 ( .A0(n4248), .A1(n3564), .B0(n6304), .B1(top_core_EC_n948), 
        .C0(top_core_EC_n1008), .Y(top_core_EC_n1290) );
  INVX1 U23196 ( .A(top_core_Plain_text[120]), .Y(n4248) );
  AOI22X1 U23197 ( .A0(top_core_EC_n950), .A1(top_core_EC_mix_out_0_), .B0(
        top_core_EC_add_out_r_0_), .B1(n3578), .Y(top_core_EC_n1008) );
  OAI221XL U23198 ( .A0(n4249), .A1(n3564), .B0(n6303), .B1(n3571), .C0(
        top_core_EC_n1007), .Y(top_core_EC_n1289) );
  INVX1 U23199 ( .A(top_core_Plain_text[121]), .Y(n4249) );
  AOI22X1 U23200 ( .A0(n3576), .A1(top_core_EC_mix_out_1_), .B0(
        top_core_EC_add_out_r_1_), .B1(n3579), .Y(top_core_EC_n1007) );
  OAI221XL U23201 ( .A0(n4250), .A1(n3564), .B0(n6302), .B1(n3572), .C0(
        top_core_EC_n1006), .Y(top_core_EC_n1288) );
  INVX1 U23202 ( .A(top_core_Plain_text[122]), .Y(n4250) );
  AOI22X1 U23203 ( .A0(n3576), .A1(top_core_EC_mix_out_2_), .B0(
        top_core_EC_add_out_r_2_), .B1(n3580), .Y(top_core_EC_n1006) );
  NAND3X1 U23204 ( .A(top_core_KE_n728), .B(n1226), .C(top_core_KE_n875), .Y(
        top_core_KE_n874) );
  NAND3X1 U23205 ( .A(top_core_KE_n728), .B(n7007), .C(top_core_KE_n878), .Y(
        top_core_KE_n877) );
  NAND3X1 U23206 ( .A(top_core_KE_n728), .B(n1226), .C(top_core_KE_n887), .Y(
        top_core_KE_n886) );
  OAI221XL U23207 ( .A0(n6768), .A1(n2241), .B0(n2249), .B1(top_core_KE_n650), 
        .C0(top_core_KE_n1954), .Y(top_core_KE_n4719) );
  INVX1 U23208 ( .A(top_core_KE_n1802), .Y(n6768) );
  AOI222X1 U23209 ( .A0(n2259), .A1(n1717), .B0(n2268), .B1(
        top_core_KE_CipherKey0_200_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_136_), .Y(top_core_KE_n1954) );
  OAI221XL U23210 ( .A0(n6428), .A1(n2243), .B0(n2248), .B1(top_core_KE_n658), 
        .C0(top_core_KE_n1970), .Y(top_core_KE_n4727) );
  INVX1 U23211 ( .A(top_core_KE_n1869), .Y(n6428) );
  AOI222X1 U23212 ( .A0(n2258), .A1(n1746), .B0(n2267), .B1(
        top_core_KE_CipherKey0_192_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_128_), .Y(top_core_KE_n1970) );
  OAI221XL U23213 ( .A0(n6765), .A1(n2241), .B0(n2249), .B1(top_core_KE_n649), 
        .C0(top_core_KE_n1952), .Y(top_core_KE_n4718) );
  INVX1 U23214 ( .A(top_core_KE_n1794), .Y(n6765) );
  AOI222X1 U23215 ( .A0(n2259), .A1(n1710), .B0(n2268), .B1(
        top_core_KE_CipherKey0_201_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_137_), .Y(top_core_KE_n1952) );
  OAI221XL U23216 ( .A0(n6425), .A1(n2241), .B0(n2248), .B1(top_core_KE_n657), 
        .C0(top_core_KE_n1968), .Y(top_core_KE_n4726) );
  INVX1 U23217 ( .A(top_core_KE_n1858), .Y(n6425) );
  AOI222X1 U23218 ( .A0(n2258), .A1(n1739), .B0(n2267), .B1(
        top_core_KE_CipherKey0_193_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_129_), .Y(top_core_KE_n1968) );
  OAI221XL U23219 ( .A0(n6761), .A1(n2241), .B0(n2249), .B1(top_core_KE_n648), 
        .C0(top_core_KE_n1950), .Y(top_core_KE_n4717) );
  INVX1 U23220 ( .A(top_core_KE_n1786), .Y(n6761) );
  AOI222X1 U23221 ( .A0(n2259), .A1(n1703), .B0(n2268), .B1(
        top_core_KE_CipherKey0_202_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_138_), .Y(top_core_KE_n1950) );
  OAI221XL U23222 ( .A0(n6418), .A1(n2239), .B0(n2248), .B1(top_core_KE_n656), 
        .C0(top_core_KE_n1966), .Y(top_core_KE_n4725) );
  INVX1 U23223 ( .A(top_core_KE_n1850), .Y(n6418) );
  AOI222X1 U23224 ( .A0(n2258), .A1(n1732), .B0(n2267), .B1(
        top_core_KE_CipherKey0_194_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_130_), .Y(top_core_KE_n1966) );
  OAI221XL U23225 ( .A0(n6758), .A1(n2241), .B0(n2249), .B1(top_core_KE_n647), 
        .C0(top_core_KE_n1948), .Y(top_core_KE_n4716) );
  INVX1 U23226 ( .A(top_core_KE_n1778), .Y(n6758) );
  AOI222X1 U23227 ( .A0(n2259), .A1(n1347), .B0(n2268), .B1(
        top_core_KE_CipherKey0_203_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_139_), .Y(top_core_KE_n1948) );
  OAI221XL U23228 ( .A0(n6421), .A1(n2237), .B0(n2248), .B1(top_core_KE_n655), 
        .C0(top_core_KE_n1964), .Y(top_core_KE_n4724) );
  INVX1 U23229 ( .A(top_core_KE_n1842), .Y(n6421) );
  AOI222X1 U23230 ( .A0(n2258), .A1(n1349), .B0(n2267), .B1(
        top_core_KE_CipherKey0_195_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_131_), .Y(top_core_KE_n1964) );
  OAI221XL U23231 ( .A0(n6755), .A1(n2241), .B0(n2249), .B1(top_core_KE_n646), 
        .C0(top_core_KE_n1946), .Y(top_core_KE_n4715) );
  INVX1 U23232 ( .A(top_core_KE_n1770), .Y(n6755) );
  AOI222X1 U23233 ( .A0(n2259), .A1(n1351), .B0(n2268), .B1(
        top_core_KE_CipherKey0_204_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_140_), .Y(top_core_KE_n1946) );
  OAI221XL U23234 ( .A0(n6414), .A1(n2242), .B0(n2248), .B1(top_core_KE_n654), 
        .C0(top_core_KE_n1962), .Y(top_core_KE_n4723) );
  INVX1 U23235 ( .A(top_core_KE_n1834), .Y(n6414) );
  AOI222X1 U23236 ( .A0(n2258), .A1(n1353), .B0(n2267), .B1(
        top_core_KE_CipherKey0_196_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_132_), .Y(top_core_KE_n1962) );
  OAI221XL U23237 ( .A0(n6752), .A1(n2241), .B0(n2249), .B1(top_core_KE_n645), 
        .C0(top_core_KE_n1944), .Y(top_core_KE_n4714) );
  INVX1 U23238 ( .A(top_core_KE_n1762), .Y(n6752) );
  AOI222X1 U23239 ( .A0(n2259), .A1(n1696), .B0(n2268), .B1(
        top_core_KE_CipherKey0_205_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_141_), .Y(top_core_KE_n1944) );
  OAI221XL U23240 ( .A0(n6411), .A1(n2243), .B0(n2248), .B1(top_core_KE_n653), 
        .C0(top_core_KE_n1960), .Y(top_core_KE_n4722) );
  INVX1 U23241 ( .A(top_core_KE_n1826), .Y(n6411) );
  AOI222X1 U23242 ( .A0(n2258), .A1(n1725), .B0(n2267), .B1(
        top_core_KE_CipherKey0_197_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_133_), .Y(top_core_KE_n1960) );
  OAI221XL U23243 ( .A0(n6687), .A1(n2241), .B0(n2249), .B1(top_core_KE_n642), 
        .C0(top_core_KE_n1938), .Y(top_core_KE_n4711) );
  INVX1 U23244 ( .A(top_core_KE_n1738), .Y(n6687) );
  AOI222X1 U23245 ( .A0(n2259), .A1(n1688), .B0(n2268), .B1(
        top_core_KE_CipherKey0_208_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_144_), .Y(top_core_KE_n1938) );
  OAI221XL U23246 ( .A0(n6680), .A1(n2241), .B0(n2249), .B1(top_core_KE_n641), 
        .C0(top_core_KE_n1936), .Y(top_core_KE_n4710) );
  INVX1 U23247 ( .A(top_core_KE_n1730), .Y(n6680) );
  AOI222X1 U23248 ( .A0(n2259), .A1(n1681), .B0(n2268), .B1(
        top_core_KE_CipherKey0_209_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_145_), .Y(top_core_KE_n1936) );
  OAI221XL U23249 ( .A0(n6665), .A1(n2241), .B0(n2249), .B1(top_core_KE_n640), 
        .C0(top_core_KE_n1934), .Y(top_core_KE_n4709) );
  INVX1 U23250 ( .A(top_core_KE_n1722), .Y(n6665) );
  AOI222X1 U23251 ( .A0(n2259), .A1(n1674), .B0(n2268), .B1(
        top_core_KE_CipherKey0_210_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_146_), .Y(top_core_KE_n1934) );
  OAI221XL U23252 ( .A0(n6632), .A1(n2242), .B0(n2250), .B1(top_core_KE_n639), 
        .C0(top_core_KE_n1932), .Y(top_core_KE_n4708) );
  INVX1 U23253 ( .A(top_core_KE_n1714), .Y(n6632) );
  AOI222X1 U23254 ( .A0(n2260), .A1(n1363), .B0(n2269), .B1(
        top_core_KE_CipherKey0_211_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_147_), .Y(top_core_KE_n1932) );
  OAI221XL U23255 ( .A0(n6537), .A1(n2242), .B0(n2250), .B1(top_core_KE_n638), 
        .C0(top_core_KE_n1930), .Y(top_core_KE_n4707) );
  INVX1 U23256 ( .A(top_core_KE_n1706), .Y(n6537) );
  AOI222X1 U23257 ( .A0(n2260), .A1(n1367), .B0(n2269), .B1(
        top_core_KE_CipherKey0_212_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_148_), .Y(top_core_KE_n1930) );
  OAI221XL U23258 ( .A0(n6447), .A1(n2242), .B0(n2250), .B1(top_core_KE_n637), 
        .C0(top_core_KE_n1928), .Y(top_core_KE_n4706) );
  INVX1 U23259 ( .A(top_core_KE_n1698), .Y(n6447) );
  AOI222X1 U23260 ( .A0(n2260), .A1(n1667), .B0(n2269), .B1(
        top_core_KE_CipherKey0_213_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_149_), .Y(top_core_KE_n1928) );
  OAI221XL U23261 ( .A0(n6399), .A1(n2242), .B0(n2250), .B1(top_core_KE_n636), 
        .C0(top_core_KE_n1926), .Y(top_core_KE_n4705) );
  INVX1 U23262 ( .A(top_core_KE_n1690), .Y(n6399) );
  AOI222X1 U23263 ( .A0(n2260), .A1(n1356), .B0(n2269), .B1(
        top_core_KE_CipherKey0_214_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_150_), .Y(top_core_KE_n1926) );
  OAI221XL U23264 ( .A0(n6391), .A1(n2241), .B0(n2249), .B1(top_core_KE_n644), 
        .C0(top_core_KE_n1942), .Y(top_core_KE_n4713) );
  INVX1 U23265 ( .A(top_core_KE_n1754), .Y(n6391) );
  AOI222X1 U23266 ( .A0(n2259), .A1(n1355), .B0(n2268), .B1(
        top_core_KE_CipherKey0_206_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_142_), .Y(top_core_KE_n1942) );
  OAI221XL U23267 ( .A0(n6382), .A1(n2238), .B0(n2248), .B1(top_core_KE_n652), 
        .C0(top_core_KE_n1958), .Y(top_core_KE_n4721) );
  INVX1 U23268 ( .A(top_core_KE_n1818), .Y(n6382) );
  AOI222X1 U23269 ( .A0(n2258), .A1(n1342), .B0(n2267), .B1(
        top_core_KE_CipherKey0_198_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_134_), .Y(top_core_KE_n1958) );
  OAI221XL U23270 ( .A0(n6335), .A1(n2242), .B0(n2250), .B1(top_core_KE_n635), 
        .C0(top_core_KE_n1924), .Y(top_core_KE_n4704) );
  INVX1 U23271 ( .A(top_core_KE_n1682), .Y(n6335) );
  AOI222X1 U23272 ( .A0(n2260), .A1(n1340), .B0(n2269), .B1(
        top_core_KE_CipherKey0_215_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_151_), .Y(top_core_KE_n1924) );
  OAI221XL U23273 ( .A0(n6326), .A1(n2241), .B0(n2249), .B1(top_core_KE_n643), 
        .C0(top_core_KE_n1940), .Y(top_core_KE_n4712) );
  INVX1 U23274 ( .A(top_core_KE_n1746), .Y(n6326) );
  AOI222X1 U23275 ( .A0(n2259), .A1(n1337), .B0(n2268), .B1(
        top_core_KE_CipherKey0_207_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_143_), .Y(top_core_KE_n1940) );
  OAI221XL U23276 ( .A0(n6322), .A1(n2241), .B0(n2249), .B1(top_core_KE_n651), 
        .C0(top_core_KE_n1956), .Y(top_core_KE_n4720) );
  INVX1 U23277 ( .A(top_core_KE_n1810), .Y(n6322) );
  AOI222X1 U23278 ( .A0(n2259), .A1(n1336), .B0(n2268), .B1(
        top_core_KE_CipherKey0_199_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_135_), .Y(top_core_KE_n1956) );
  OAI221XL U23279 ( .A0(top_core_KE_n1805), .A1(n2347), .B0(n2290), .B1(n6997), 
        .C0(top_core_KE_n2662), .Y(top_core_KE_n4912) );
  AOI222X1 U23280 ( .A0(n2343), .A1(top_core_KE_n1809), .B0(n2324), .B1(
        top_core_KE_CipherKey0_7_), .C0(n2333), .C1(top_core_KE_n1807), .Y(
        top_core_KE_n2662) );
  OAI221XL U23281 ( .A0(top_core_KE_n1741), .A1(n2348), .B0(n2290), .B1(n6993), 
        .C0(top_core_KE_n2630), .Y(top_core_KE_n4904) );
  AOI222X1 U23282 ( .A0(n2343), .A1(top_core_KE_n1745), .B0(n2324), .B1(
        top_core_KE_CipherKey0_15_), .C0(n2333), .C1(top_core_KE_n1743), .Y(
        top_core_KE_n2630) );
  OAI221XL U23283 ( .A0(top_core_KE_n1677), .A1(n2348), .B0(n2289), .B1(n6992), 
        .C0(top_core_KE_n2598), .Y(top_core_KE_n4896) );
  AOI222X1 U23284 ( .A0(n2342), .A1(top_core_KE_n1681), .B0(n2323), .B1(
        top_core_KE_CipherKey0_23_), .C0(n2332), .C1(top_core_KE_n1679), .Y(
        top_core_KE_n2598) );
  OAI221XL U23285 ( .A0(n6688), .A1(n2243), .B0(n2251), .B1(n6689), .C0(
        top_core_KE_n1892), .Y(top_core_KE_n4680) );
  INVX1 U23286 ( .A(top_core_KE_n1482), .Y(n6688) );
  AOI222X1 U23287 ( .A0(top_core_KE_n1875), .A1(top_core_KE_prev_key1_reg_112_), .B0(n2271), .B1(top_core_KE_CipherKey0_240_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_176_), .Y(top_core_KE_n1892) );
  OAI221XL U23288 ( .A0(n6681), .A1(n2243), .B0(n2251), .B1(n6682), .C0(
        top_core_KE_n1891), .Y(top_core_KE_n4679) );
  INVX1 U23289 ( .A(top_core_KE_n1474), .Y(n6681) );
  AOI222X1 U23290 ( .A0(top_core_KE_n1875), .A1(top_core_KE_prev_key1_reg_113_), .B0(n2271), .B1(top_core_KE_CipherKey0_241_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_177_), .Y(top_core_KE_n1891) );
  OAI221XL U23291 ( .A0(n6666), .A1(n2243), .B0(n2251), .B1(n6667), .C0(
        top_core_KE_n1890), .Y(top_core_KE_n4678) );
  INVX1 U23292 ( .A(top_core_KE_n1466), .Y(n6666) );
  AOI222X1 U23293 ( .A0(top_core_KE_n1875), .A1(top_core_KE_prev_key1_reg_114_), .B0(n2271), .B1(top_core_KE_CipherKey0_242_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_178_), .Y(top_core_KE_n1890) );
  OAI221XL U23294 ( .A0(n6638), .A1(n2243), .B0(n2251), .B1(n6639), .C0(
        top_core_KE_n1889), .Y(top_core_KE_n4677) );
  INVX1 U23295 ( .A(top_core_KE_n1458), .Y(n6638) );
  AOI222X1 U23296 ( .A0(top_core_KE_n1875), .A1(top_core_KE_prev_key1_reg_115_), .B0(n2271), .B1(top_core_KE_CipherKey0_243_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_179_), .Y(top_core_KE_n1889) );
  OAI221XL U23297 ( .A0(n6559), .A1(n2243), .B0(n2251), .B1(n6560), .C0(
        top_core_KE_n1888), .Y(top_core_KE_n4676) );
  INVX1 U23298 ( .A(top_core_KE_n1450), .Y(n6559) );
  AOI222X1 U23299 ( .A0(top_core_KE_n1875), .A1(top_core_KE_prev_key1_reg_116_), .B0(n2271), .B1(top_core_KE_CipherKey0_244_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_180_), .Y(top_core_KE_n1888) );
  OAI221XL U23300 ( .A0(n6479), .A1(n2243), .B0(n2251), .B1(n6480), .C0(
        top_core_KE_n1887), .Y(top_core_KE_n4675) );
  INVX1 U23301 ( .A(top_core_KE_n1442), .Y(n6479) );
  AOI222X1 U23302 ( .A0(top_core_KE_n1875), .A1(top_core_KE_prev_key1_reg_117_), .B0(n2271), .B1(top_core_KE_CipherKey0_245_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_181_), .Y(top_core_KE_n1887) );
  OAI221XL U23303 ( .A0(n6401), .A1(n2243), .B0(n2251), .B1(n6402), .C0(
        top_core_KE_n1886), .Y(top_core_KE_n4674) );
  INVX1 U23304 ( .A(top_core_KE_n1434), .Y(n6401) );
  AOI222X1 U23305 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_118_), .B0(n2271), .B1(top_core_KE_CipherKey0_246_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_182_), .Y(top_core_KE_n1886) );
  OAI221XL U23306 ( .A0(n6393), .A1(n2243), .B0(n2251), .B1(n6394), .C0(
        top_core_KE_n1885), .Y(top_core_KE_n4673) );
  INVX1 U23307 ( .A(top_core_KE_n1426), .Y(n6393) );
  AOI222X1 U23308 ( .A0(top_core_KE_n1875), .A1(top_core_KE_prev_key1_reg_119_), .B0(n2271), .B1(top_core_KE_CipherKey0_247_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_183_), .Y(top_core_KE_n1885) );
  OAI221XL U23309 ( .A0(top_core_KE_n1613), .A1(n2349), .B0(n2288), .B1(n6358), 
        .C0(top_core_KE_n2558), .Y(top_core_KE_n4888) );
  AOI222X1 U23310 ( .A0(n2342), .A1(top_core_KE_n1617), .B0(n2323), .B1(
        top_core_KE_CipherKey0_31_), .C0(n2332), .C1(top_core_KE_n1615), .Y(
        top_core_KE_n2558) );
  OAI221XL U23311 ( .A0(top_core_KE_n1653), .A1(n2349), .B0(n2289), .B1(n1171), 
        .C0(top_core_KE_n2583), .Y(top_core_KE_n4893) );
  AOI222X1 U23312 ( .A0(n2342), .A1(top_core_KE_n1657), .B0(n2323), .B1(
        top_core_KE_CipherKey0_26_), .C0(n2332), .C1(top_core_KE_n1655), .Y(
        top_core_KE_n2583) );
  OAI221XL U23313 ( .A0(n6343), .A1(n2241), .B0(top_core_KE_n1873), .B1(n6341), 
        .C0(top_core_KE_n1874), .Y(top_core_KE_n4665) );
  INVX1 U23314 ( .A(top_core_KE_n1362), .Y(n6343) );
  AOI222X1 U23315 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_127_), .B0(n2266), .B1(top_core_KE_CipherKey0_255_), .C0(top_core_KE_n1877), .C1(
        top_core_KE_CipherKey0_191_), .Y(top_core_KE_n1874) );
  OAI221XL U23316 ( .A0(n6769), .A1(n2236), .B0(n2247), .B1(n6982), .C0(
        top_core_KE_n1900), .Y(top_core_KE_n4688) );
  INVX1 U23317 ( .A(top_core_KE_n1546), .Y(n6769) );
  AOI222X1 U23318 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_104_), .B0(n2270), .B1(top_core_KE_CipherKey0_232_), .C0(top_core_KE_n1877), .C1(
        top_core_KE_CipherKey0_168_), .Y(top_core_KE_n1900) );
  OAI221XL U23319 ( .A0(n6429), .A1(n2240), .B0(n2251), .B1(n6977), .C0(
        top_core_KE_n1907), .Y(top_core_KE_n4695) );
  INVX1 U23320 ( .A(top_core_KE_n1610), .Y(n6429) );
  AOI222X1 U23321 ( .A0(n2255), .A1(top_core_KE_prev_key1_reg_96_), .B0(n2270), 
        .B1(top_core_KE_CipherKey0_224_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_160_), .Y(top_core_KE_n1907) );
  OAI221XL U23322 ( .A0(n6766), .A1(n2237), .B0(n2244), .B1(n6972), .C0(
        top_core_KE_n1899), .Y(top_core_KE_n4687) );
  INVX1 U23323 ( .A(top_core_KE_n1538), .Y(n6766) );
  AOI222X1 U23324 ( .A0(n2258), .A1(top_core_KE_prev_key1_reg_105_), .B0(n2270), .B1(top_core_KE_CipherKey0_233_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_169_), .Y(top_core_KE_n1899) );
  OAI221XL U23325 ( .A0(n6426), .A1(n2242), .B0(n2246), .B1(n6967), .C0(
        top_core_KE_n1906), .Y(top_core_KE_n4694) );
  INVX1 U23326 ( .A(top_core_KE_n1602), .Y(n6426) );
  AOI222X1 U23327 ( .A0(n2259), .A1(top_core_KE_prev_key1_reg_97_), .B0(n2270), 
        .B1(top_core_KE_CipherKey0_225_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_161_), .Y(top_core_KE_n1906) );
  OAI221XL U23328 ( .A0(n6762), .A1(n2243), .B0(n2245), .B1(n6961), .C0(
        top_core_KE_n1898), .Y(top_core_KE_n4686) );
  INVX1 U23329 ( .A(top_core_KE_n1530), .Y(n6762) );
  AOI222X1 U23330 ( .A0(top_core_KE_n1875), .A1(top_core_KE_prev_key1_reg_106_), .B0(n2270), .B1(top_core_KE_CipherKey0_234_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_170_), .Y(top_core_KE_n1898) );
  OAI221XL U23331 ( .A0(n6417), .A1(n2236), .B0(n2244), .B1(n6955), .C0(
        top_core_KE_n2698), .Y(top_core_KE_n4920) );
  INVX1 U23332 ( .A(top_core_KE_n1594), .Y(n6417) );
  AOI222X1 U23333 ( .A0(n2254), .A1(top_core_KE_prev_key1_reg_98_), .B0(n2264), 
        .B1(top_core_KE_CipherKey0_226_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_162_), .Y(top_core_KE_n2698) );
  OAI221XL U23334 ( .A0(n6759), .A1(n2238), .B0(n2250), .B1(n6945), .C0(
        top_core_KE_n1897), .Y(top_core_KE_n4685) );
  INVX1 U23335 ( .A(top_core_KE_n1522), .Y(n6759) );
  AOI222X1 U23336 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_107_), .B0(n2270), .B1(top_core_KE_CipherKey0_235_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_171_), .Y(top_core_KE_n1897) );
  OAI221XL U23337 ( .A0(n6422), .A1(n2236), .B0(n2248), .B1(n6930), .C0(
        top_core_KE_n1905), .Y(top_core_KE_n4693) );
  INVX1 U23338 ( .A(top_core_KE_n1586), .Y(n6422) );
  AOI222X1 U23339 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_99_), .B0(n2270), 
        .B1(top_core_KE_CipherKey0_227_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_163_), .Y(top_core_KE_n1905) );
  OAI221XL U23340 ( .A0(n6756), .A1(n2243), .B0(n2251), .B1(n6900), .C0(
        top_core_KE_n1896), .Y(top_core_KE_n4684) );
  INVX1 U23341 ( .A(top_core_KE_n1514), .Y(n6756) );
  AOI222X1 U23342 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_108_), .B0(n2271), .B1(top_core_KE_CipherKey0_236_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_172_), .Y(top_core_KE_n1896) );
  OAI221XL U23343 ( .A0(n6415), .A1(n2240), .B0(n2249), .B1(n6854), .C0(
        top_core_KE_n1904), .Y(top_core_KE_n4692) );
  INVX1 U23344 ( .A(top_core_KE_n1578), .Y(n6415) );
  AOI222X1 U23345 ( .A0(n2260), .A1(top_core_KE_prev_key1_reg_100_), .B0(n2270), .B1(top_core_KE_CipherKey0_228_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_164_), .Y(top_core_KE_n1904) );
  OAI221XL U23346 ( .A0(n6753), .A1(n2243), .B0(n2251), .B1(n6820), .C0(
        top_core_KE_n1895), .Y(top_core_KE_n4683) );
  INVX1 U23347 ( .A(top_core_KE_n1506), .Y(n6753) );
  AOI222X1 U23348 ( .A0(top_core_KE_n1875), .A1(top_core_KE_prev_key1_reg_109_), .B0(n2271), .B1(top_core_KE_CipherKey0_237_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_173_), .Y(top_core_KE_n1895) );
  OAI221XL U23349 ( .A0(n6412), .A1(n2241), .B0(n2247), .B1(n6781), .C0(
        top_core_KE_n1903), .Y(top_core_KE_n4691) );
  INVX1 U23350 ( .A(top_core_KE_n1570), .Y(n6412) );
  AOI222X1 U23351 ( .A0(n2254), .A1(top_core_KE_prev_key1_reg_101_), .B0(n2270), .B1(top_core_KE_CipherKey0_229_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_165_), .Y(top_core_KE_n1903) );
  OAI221XL U23352 ( .A0(n6716), .A1(n2243), .B0(n2251), .B1(n6717), .C0(
        top_core_KE_n1894), .Y(top_core_KE_n4682) );
  INVX1 U23353 ( .A(top_core_KE_n1498), .Y(n6716) );
  AOI222X1 U23354 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_110_), .B0(n2271), .B1(top_core_KE_CipherKey0_238_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_174_), .Y(top_core_KE_n1894) );
  OAI221XL U23355 ( .A0(n6383), .A1(n2239), .B0(n2251), .B1(n6384), .C0(
        top_core_KE_n1902), .Y(top_core_KE_n4690) );
  INVX1 U23356 ( .A(top_core_KE_n1562), .Y(n6383) );
  AOI222X1 U23357 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_102_), .B0(n2270), .B1(top_core_KE_CipherKey0_230_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_166_), .Y(top_core_KE_n1902) );
  OAI221XL U23358 ( .A0(n6376), .A1(n2237), .B0(n2244), .B1(n6377), .C0(
        top_core_KE_n1901), .Y(top_core_KE_n4689) );
  INVX1 U23359 ( .A(top_core_KE_n1554), .Y(n6376) );
  AOI222X1 U23360 ( .A0(n2255), .A1(top_core_KE_prev_key1_reg_103_), .B0(n2270), .B1(top_core_KE_CipherKey0_231_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_167_), .Y(top_core_KE_n1901) );
  OAI221XL U23361 ( .A0(n6327), .A1(n2243), .B0(n2251), .B1(n6328), .C0(
        top_core_KE_n1893), .Y(top_core_KE_n4681) );
  INVX1 U23362 ( .A(top_core_KE_n1490), .Y(n6327) );
  AOI222X1 U23363 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_111_), .B0(n2271), .B1(top_core_KE_CipherKey0_239_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_175_), .Y(top_core_KE_n1893) );
  OAI221XL U23364 ( .A0(top_core_KE_n1972), .A1(n2243), .B0(n2248), .B1(n6337), 
        .C0(top_core_KE_n1973), .Y(top_core_KE_n4728) );
  AOI222X1 U23365 ( .A0(n2258), .A1(top_core_KE_prev_key1_reg_63_), .B0(n2267), 
        .B1(top_core_KE_CipherKey0_191_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_127_), .Y(top_core_KE_n1973) );
  XNOR2X1 U23366 ( .A(top_core_KE_n1974), .B(top_core_KE_n1975), .Y(
        top_core_KE_n1972) );
  OAI221XL U23367 ( .A0(n6464), .A1(n2239), .B0(top_core_KE_n1873), .B1(n6695), 
        .C0(top_core_KE_n1884), .Y(top_core_KE_n4672) );
  INVX1 U23368 ( .A(top_core_KE_n1418), .Y(n6464) );
  AOI222X1 U23369 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_120_), .B0(
        top_core_KE_n1876), .B1(top_core_KE_CipherKey0_248_), .C0(
        top_core_KE_n1877), .C1(top_core_KE_CipherKey0_184_), .Y(
        top_core_KE_n1884) );
  OAI221XL U23370 ( .A0(n6459), .A1(n2237), .B0(top_core_KE_n1873), .B1(n6674), 
        .C0(top_core_KE_n1882), .Y(top_core_KE_n4670) );
  INVX1 U23371 ( .A(top_core_KE_n1402), .Y(n6459) );
  AOI222X1 U23372 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_122_), .B0(n2267), .B1(top_core_KE_CipherKey0_250_), .C0(top_core_KE_n1877), .C1(
        top_core_KE_CipherKey0_186_), .Y(top_core_KE_n1882) );
  OAI221XL U23373 ( .A0(n6456), .A1(n2242), .B0(top_core_KE_n1873), .B1(n6655), 
        .C0(top_core_KE_n1881), .Y(top_core_KE_n4669) );
  INVX1 U23374 ( .A(top_core_KE_n1394), .Y(n6456) );
  AOI222X1 U23375 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_123_), .B0(n2268), .B1(top_core_KE_CipherKey0_251_), .C0(top_core_KE_n1877), .C1(
        top_core_KE_CipherKey0_187_), .Y(top_core_KE_n1881) );
  OAI221XL U23376 ( .A0(n6453), .A1(n2238), .B0(n2244), .B1(n6607), .C0(
        top_core_KE_n1880), .Y(top_core_KE_n4668) );
  INVX1 U23377 ( .A(top_core_KE_n1386), .Y(n6453) );
  AOI222X1 U23378 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_124_), .B0(n2271), .B1(top_core_KE_CipherKey0_252_), .C0(top_core_KE_n1877), .C1(
        top_core_KE_CipherKey0_188_), .Y(top_core_KE_n1880) );
  OAI221XL U23379 ( .A0(n6450), .A1(n2238), .B0(n2249), .B1(n6524), .C0(
        top_core_KE_n1879), .Y(top_core_KE_n4667) );
  INVX1 U23380 ( .A(top_core_KE_n1378), .Y(n6450) );
  AOI222X1 U23381 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_125_), .B0(n2265), .B1(top_core_KE_CipherKey0_253_), .C0(top_core_KE_n1877), .C1(
        top_core_KE_CipherKey0_189_), .Y(top_core_KE_n1879) );
  OAI221XL U23382 ( .A0(n6436), .A1(n2236), .B0(n2250), .B1(n6435), .C0(
        top_core_KE_n1878), .Y(top_core_KE_n4666) );
  INVX1 U23383 ( .A(top_core_KE_n1370), .Y(n6436) );
  AOI222X1 U23384 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_126_), .B0(n2270), .B1(top_core_KE_CipherKey0_254_), .C0(top_core_KE_n1877), .C1(
        top_core_KE_CipherKey0_190_), .Y(top_core_KE_n1878) );
  OAI221XL U23385 ( .A0(n6316), .A1(n2240), .B0(n2248), .B1(n6314), .C0(
        top_core_KE_n1883), .Y(top_core_KE_n4671) );
  INVX1 U23386 ( .A(top_core_KE_n1410), .Y(n6316) );
  AOI222X1 U23387 ( .A0(n2261), .A1(top_core_KE_prev_key1_reg_121_), .B0(n2269), .B1(top_core_KE_CipherKey0_249_), .C0(top_core_KE_n1877), .C1(
        top_core_KE_CipherKey0_185_), .Y(top_core_KE_n1883) );
  OAI221XL U23388 ( .A0(top_core_KE_n2073), .A1(n2238), .B0(top_core_KE_n1873), 
        .B1(n6975), .C0(top_core_KE_n2074), .Y(top_core_KE_n4759) );
  AOI222X1 U23389 ( .A0(n2254), .A1(top_core_KE_prev_key1_reg_32_), .B0(
        top_core_KE_n1876), .B1(top_core_KE_CipherKey0_160_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_96_), .Y(top_core_KE_n2074) );
  XNOR2X1 U23390 ( .A(top_core_KE_new_sboxw_192_24_), .B(top_core_KE_n2075), 
        .Y(top_core_KE_n2073) );
  OAI221XL U23391 ( .A0(top_core_KE_n2070), .A1(n2238), .B0(top_core_KE_n1873), 
        .B1(n6965), .C0(top_core_KE_n2071), .Y(top_core_KE_n4758) );
  AOI222X1 U23392 ( .A0(n2259), .A1(top_core_KE_prev_key1_reg_33_), .B0(
        top_core_KE_n1876), .B1(top_core_KE_CipherKey0_161_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_97_), .Y(top_core_KE_n2071) );
  XNOR2X1 U23393 ( .A(top_core_KE_new_sboxw_192_25_), .B(top_core_KE_n2072), 
        .Y(top_core_KE_n2070) );
  OAI221XL U23394 ( .A0(top_core_KE_n2043), .A1(n2239), .B0(n2246), .B1(n6959), 
        .C0(top_core_KE_n2044), .Y(top_core_KE_n4749) );
  AOI222X1 U23395 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_42_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_170_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_106_), .Y(top_core_KE_n2044) );
  XNOR2X1 U23396 ( .A(top_core_KE_new_sboxw_192_2_), .B(top_core_KE_n2045), 
        .Y(top_core_KE_n2043) );
  OAI221XL U23397 ( .A0(top_core_KE_n2067), .A1(n2238), .B0(top_core_KE_n1873), 
        .B1(n6953), .C0(top_core_KE_n2068), .Y(top_core_KE_n4757) );
  AOI222X1 U23398 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_34_), .B0(
        top_core_KE_n1876), .B1(top_core_KE_CipherKey0_162_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_98_), .Y(top_core_KE_n2068) );
  XNOR2X1 U23399 ( .A(top_core_KE_new_sboxw_192_26_), .B(top_core_KE_n2069), 
        .Y(top_core_KE_n2067) );
  OAI221XL U23400 ( .A0(top_core_KE_n2040), .A1(n2239), .B0(n2246), .B1(n6938), 
        .C0(top_core_KE_n2041), .Y(top_core_KE_n4748) );
  AOI222X1 U23401 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_43_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_171_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_107_), .Y(top_core_KE_n2041) );
  XNOR2X1 U23402 ( .A(top_core_KE_new_sboxw_192_3_), .B(top_core_KE_n2042), 
        .Y(top_core_KE_n2040) );
  OAI221XL U23403 ( .A0(top_core_KE_n2037), .A1(n2239), .B0(n2246), .B1(n6877), 
        .C0(top_core_KE_n2038), .Y(top_core_KE_n4747) );
  AOI222X1 U23404 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_44_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_172_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_108_), .Y(top_core_KE_n2038) );
  XNOR2X1 U23405 ( .A(top_core_KE_new_sboxw_192_4_), .B(top_core_KE_n2039), 
        .Y(top_core_KE_n2037) );
  OAI221XL U23406 ( .A0(top_core_KE_n2034), .A1(n2239), .B0(n2246), .B1(n6810), 
        .C0(top_core_KE_n2035), .Y(top_core_KE_n4746) );
  AOI222X1 U23407 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_45_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_173_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_109_), .Y(top_core_KE_n2035) );
  XNOR2X1 U23408 ( .A(top_core_KE_new_sboxw_192_5_), .B(top_core_KE_n2036), 
        .Y(top_core_KE_n2034) );
  OAI221XL U23409 ( .A0(top_core_KE_n2000), .A1(n2240), .B0(n2247), .B1(n6692), 
        .C0(top_core_KE_n2001), .Y(top_core_KE_n4735) );
  AOI222X1 U23410 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_56_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_184_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_120_), .Y(top_core_KE_n2001) );
  XNOR2X1 U23411 ( .A(top_core_KE_n2002), .B(top_core_KE_n2003), .Y(
        top_core_KE_n2000) );
  OAI221XL U23412 ( .A0(top_core_KE_n2025), .A1(n2240), .B0(n2247), .B1(n6685), 
        .C0(top_core_KE_n2026), .Y(top_core_KE_n4743) );
  AOI222X1 U23413 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_48_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_176_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_112_), .Y(top_core_KE_n2026) );
  XNOR2X1 U23414 ( .A(top_core_KE_new_sboxw_192_8_), .B(top_core_KE_n2027), 
        .Y(top_core_KE_n2025) );
  OAI221XL U23415 ( .A0(top_core_KE_n2022), .A1(n2240), .B0(n2247), .B1(n6678), 
        .C0(top_core_KE_n2023), .Y(top_core_KE_n4742) );
  AOI222X1 U23416 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_49_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_177_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_113_), .Y(top_core_KE_n2023) );
  XNOR2X1 U23417 ( .A(top_core_KE_new_sboxw_192_9_), .B(top_core_KE_n2024), 
        .Y(top_core_KE_n2022) );
  OAI221XL U23418 ( .A0(top_core_KE_n1992), .A1(n2240), .B0(n2247), .B1(n6671), 
        .C0(top_core_KE_n1993), .Y(top_core_KE_n4733) );
  AOI222X1 U23419 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_58_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_186_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_122_), .Y(top_core_KE_n1993) );
  XNOR2X1 U23420 ( .A(top_core_KE_n1994), .B(top_core_KE_n1995), .Y(
        top_core_KE_n1992) );
  OAI221XL U23421 ( .A0(top_core_KE_n2019), .A1(n2240), .B0(n2247), .B1(n6663), 
        .C0(top_core_KE_n2020), .Y(top_core_KE_n4741) );
  AOI222X1 U23422 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_50_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_178_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_114_), .Y(top_core_KE_n2020) );
  XNOR2X1 U23423 ( .A(top_core_KE_new_sboxw_192_10_), .B(top_core_KE_n2021), 
        .Y(top_core_KE_n2019) );
  OAI221XL U23424 ( .A0(top_core_KE_n1988), .A1(n2236), .B0(n2248), .B1(n6647), 
        .C0(top_core_KE_n1989), .Y(top_core_KE_n4732) );
  AOI222X1 U23425 ( .A0(n2258), .A1(top_core_KE_prev_key1_reg_59_), .B0(n2267), 
        .B1(top_core_KE_CipherKey0_187_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_123_), .Y(top_core_KE_n1989) );
  XNOR2X1 U23426 ( .A(top_core_KE_n1990), .B(top_core_KE_n1991), .Y(
        top_core_KE_n1988) );
  OAI221XL U23427 ( .A0(top_core_KE_n2016), .A1(n2240), .B0(n2247), .B1(n6630), 
        .C0(top_core_KE_n2017), .Y(top_core_KE_n4740) );
  AOI222X1 U23428 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_51_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_179_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_115_), .Y(top_core_KE_n2017) );
  XNOR2X1 U23429 ( .A(top_core_KE_new_sboxw_192_11_), .B(top_core_KE_n2018), 
        .Y(top_core_KE_n2016) );
  OAI221XL U23430 ( .A0(top_core_KE_n1984), .A1(n2240), .B0(n2248), .B1(n6583), 
        .C0(top_core_KE_n1985), .Y(top_core_KE_n4731) );
  AOI222X1 U23431 ( .A0(n2258), .A1(top_core_KE_prev_key1_reg_60_), .B0(n2267), 
        .B1(top_core_KE_CipherKey0_188_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_124_), .Y(top_core_KE_n1985) );
  XNOR2X1 U23432 ( .A(top_core_KE_n1986), .B(top_core_KE_n1987), .Y(
        top_core_KE_n1984) );
  OAI221XL U23433 ( .A0(top_core_KE_n2013), .A1(n2240), .B0(n2247), .B1(n6535), 
        .C0(top_core_KE_n2014), .Y(top_core_KE_n4739) );
  AOI222X1 U23434 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_52_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_180_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_116_), .Y(top_core_KE_n2014) );
  XNOR2X1 U23435 ( .A(top_core_KE_new_sboxw_192_12_), .B(top_core_KE_n2015), 
        .Y(top_core_KE_n2013) );
  OAI221XL U23436 ( .A0(top_core_KE_n1980), .A1(n2241), .B0(n2248), .B1(n6513), 
        .C0(top_core_KE_n1981), .Y(top_core_KE_n4730) );
  AOI222X1 U23437 ( .A0(n2258), .A1(top_core_KE_prev_key1_reg_61_), .B0(n2267), 
        .B1(top_core_KE_CipherKey0_189_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_125_), .Y(top_core_KE_n1981) );
  XNOR2X1 U23438 ( .A(top_core_KE_n1982), .B(top_core_KE_n1983), .Y(
        top_core_KE_n1980) );
  OAI221XL U23439 ( .A0(top_core_KE_n2010), .A1(n2240), .B0(n2247), .B1(n6444), 
        .C0(top_core_KE_n2011), .Y(top_core_KE_n4738) );
  AOI222X1 U23440 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_53_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_181_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_117_), .Y(top_core_KE_n2011) );
  XNOR2X1 U23441 ( .A(top_core_KE_new_sboxw_192_13_), .B(top_core_KE_n2012), 
        .Y(top_core_KE_n2010) );
  OAI221XL U23442 ( .A0(top_core_KE_n1976), .A1(n2239), .B0(n2248), .B1(n6405), 
        .C0(top_core_KE_n1977), .Y(top_core_KE_n4729) );
  AOI222X1 U23443 ( .A0(n2258), .A1(top_core_KE_prev_key1_reg_62_), .B0(n2267), 
        .B1(top_core_KE_CipherKey0_190_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_126_), .Y(top_core_KE_n1977) );
  XNOR2X1 U23444 ( .A(top_core_KE_n1978), .B(top_core_KE_n1979), .Y(
        top_core_KE_n1976) );
  OAI221XL U23445 ( .A0(top_core_KE_n2007), .A1(n2240), .B0(n2247), .B1(n6396), 
        .C0(top_core_KE_n2008), .Y(top_core_KE_n4737) );
  AOI222X1 U23446 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_54_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_182_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_118_), .Y(top_core_KE_n2008) );
  XNOR2X1 U23447 ( .A(top_core_KE_new_sboxw_192_14_), .B(top_core_KE_n2009), 
        .Y(top_core_KE_n2007) );
  OAI221XL U23448 ( .A0(top_core_KE_n2031), .A1(n2239), .B0(n2246), .B1(n6388), 
        .C0(top_core_KE_n2032), .Y(top_core_KE_n4745) );
  AOI222X1 U23449 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_46_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_174_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_110_), .Y(top_core_KE_n2032) );
  XNOR2X1 U23450 ( .A(top_core_KE_new_sboxw_192_6_), .B(top_core_KE_n2033), 
        .Y(top_core_KE_n2031) );
  OAI221XL U23451 ( .A0(top_core_KE_n2004), .A1(n2240), .B0(n2247), .B1(n6332), 
        .C0(top_core_KE_n2005), .Y(top_core_KE_n4736) );
  AOI222X1 U23452 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_55_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_183_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_119_), .Y(top_core_KE_n2005) );
  XNOR2X1 U23453 ( .A(top_core_KE_new_sboxw_192_15_), .B(top_core_KE_n2006), 
        .Y(top_core_KE_n2004) );
  OAI221XL U23454 ( .A0(top_core_KE_n2028), .A1(n2240), .B0(n2247), .B1(n6323), 
        .C0(top_core_KE_n2029), .Y(top_core_KE_n4744) );
  AOI222X1 U23455 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_47_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_175_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_111_), .Y(top_core_KE_n2029) );
  XNOR2X1 U23456 ( .A(top_core_KE_new_sboxw_192_7_), .B(top_core_KE_n2030), 
        .Y(top_core_KE_n2028) );
  OAI221XL U23457 ( .A0(top_core_KE_n1996), .A1(n2240), .B0(n2247), .B1(n6310), 
        .C0(top_core_KE_n1997), .Y(top_core_KE_n4734) );
  AOI222X1 U23458 ( .A0(n2257), .A1(top_core_KE_prev_key1_reg_57_), .B0(n2266), 
        .B1(top_core_KE_CipherKey0_185_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_121_), .Y(top_core_KE_n1997) );
  XNOR2X1 U23459 ( .A(top_core_KE_n1998), .B(top_core_KE_n1999), .Y(
        top_core_KE_n1996) );
  OAI221XL U23460 ( .A0(top_core_KE_n2049), .A1(n2239), .B0(n2246), .B1(n6980), 
        .C0(top_core_KE_n2050), .Y(top_core_KE_n4751) );
  AOI222X1 U23461 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_40_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_168_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_104_), .Y(top_core_KE_n2050) );
  XNOR2X1 U23462 ( .A(top_core_KE_new_sboxw_192_0_), .B(top_core_KE_n2051), 
        .Y(top_core_KE_n2049) );
  OAI221XL U23463 ( .A0(top_core_KE_n2046), .A1(n2239), .B0(n2246), .B1(n6970), 
        .C0(top_core_KE_n2047), .Y(top_core_KE_n4750) );
  AOI222X1 U23464 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_41_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_169_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_105_), .Y(top_core_KE_n2047) );
  XNOR2X1 U23465 ( .A(top_core_KE_new_sboxw_192_1_), .B(top_core_KE_n2048), 
        .Y(top_core_KE_n2046) );
  OAI221XL U23466 ( .A0(top_core_KE_n2064), .A1(n2239), .B0(n2246), .B1(n6923), 
        .C0(top_core_KE_n2065), .Y(top_core_KE_n4756) );
  AOI222X1 U23467 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_35_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_163_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_99_), .Y(top_core_KE_n2065) );
  XNOR2X1 U23468 ( .A(top_core_KE_new_sboxw_192_27_), .B(top_core_KE_n2066), 
        .Y(top_core_KE_n2064) );
  OAI221XL U23469 ( .A0(top_core_KE_n2061), .A1(n2239), .B0(n2246), .B1(n6831), 
        .C0(top_core_KE_n2062), .Y(top_core_KE_n4755) );
  AOI222X1 U23470 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_36_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_164_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_100_), .Y(top_core_KE_n2062) );
  XNOR2X1 U23471 ( .A(top_core_KE_new_sboxw_192_28_), .B(top_core_KE_n2063), 
        .Y(top_core_KE_n2061) );
  OAI221XL U23472 ( .A0(top_core_KE_n2058), .A1(n2239), .B0(n2246), .B1(n6747), 
        .C0(top_core_KE_n2059), .Y(top_core_KE_n4754) );
  AOI222X1 U23473 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_37_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_165_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_101_), .Y(top_core_KE_n2059) );
  XNOR2X1 U23474 ( .A(top_core_KE_new_sboxw_192_29_), .B(top_core_KE_n2060), 
        .Y(top_core_KE_n2058) );
  OAI221XL U23475 ( .A0(top_core_KE_n2055), .A1(n2239), .B0(n2246), .B1(n6380), 
        .C0(top_core_KE_n2056), .Y(top_core_KE_n4753) );
  AOI222X1 U23476 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_38_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_166_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_102_), .Y(top_core_KE_n2056) );
  XNOR2X1 U23477 ( .A(top_core_KE_new_sboxw_192_30_), .B(top_core_KE_n2057), 
        .Y(top_core_KE_n2055) );
  OAI221XL U23478 ( .A0(top_core_KE_n2052), .A1(n2239), .B0(n2246), .B1(n6319), 
        .C0(top_core_KE_n2053), .Y(top_core_KE_n4752) );
  AOI222X1 U23479 ( .A0(n2256), .A1(top_core_KE_prev_key1_reg_39_), .B0(n2265), 
        .B1(top_core_KE_CipherKey0_167_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_103_), .Y(top_core_KE_n2053) );
  XNOR2X1 U23480 ( .A(top_core_KE_new_sboxw_192_31_), .B(top_core_KE_n2054), 
        .Y(top_core_KE_n2052) );
  OAI221XL U23481 ( .A0(top_core_KE_n1757), .A1(n2348), .B0(n2290), .B1(n1796), 
        .C0(top_core_KE_n2638), .Y(top_core_KE_n4906) );
  AOI222X1 U23482 ( .A0(n2343), .A1(top_core_KE_n1761), .B0(n2324), .B1(
        top_core_KE_CipherKey0_13_), .C0(n2333), .C1(top_core_KE_n1759), .Y(
        top_core_KE_n2638) );
  OAI221XL U23483 ( .A0(top_core_KE_n1821), .A1(n2347), .B0(n2290), .B1(n1817), 
        .C0(top_core_KE_n2670), .Y(top_core_KE_n4914) );
  AOI222X1 U23484 ( .A0(n2343), .A1(top_core_KE_n1825), .B0(n2324), .B1(
        top_core_KE_CipherKey0_5_), .C0(n2333), .C1(top_core_KE_n1823), .Y(
        top_core_KE_n2670) );
  OAI221XL U23485 ( .A0(top_core_KE_n1693), .A1(n2348), .B0(n2289), .B1(n1775), 
        .C0(top_core_KE_n2606), .Y(top_core_KE_n4898) );
  AOI222X1 U23486 ( .A0(n2342), .A1(top_core_KE_n1697), .B0(n2323), .B1(
        top_core_KE_CipherKey0_21_), .C0(n2332), .C1(top_core_KE_n1695), .Y(
        top_core_KE_n2606) );
  OAI221XL U23487 ( .A0(top_core_KE_n2148), .A1(n2236), .B0(n2244), .B1(n6996), 
        .C0(top_core_KE_n2149), .Y(top_core_KE_n4784) );
  AOI222X1 U23488 ( .A0(n2254), .A1(n1335), .B0(n2264), .B1(
        top_core_KE_CipherKey0_135_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_71_), .Y(top_core_KE_n2149) );
  XNOR2X1 U23489 ( .A(top_core_KE_n2150), .B(n6423), .Y(top_core_KE_n2148) );
  INVX1 U23490 ( .A(top_core_KE_new_sboxw_192_31_), .Y(n6423) );
  OAI221XL U23491 ( .A0(top_core_KE_n2145), .A1(n2236), .B0(n2244), .B1(n6984), 
        .C0(top_core_KE_n2146), .Y(top_core_KE_n4783) );
  AOI222X1 U23492 ( .A0(n2254), .A1(n1810), .B0(n2264), .B1(
        top_core_KE_CipherKey0_136_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_72_), .Y(top_core_KE_n2146) );
  XNOR2X1 U23493 ( .A(top_core_KE_n2147), .B(n6767), .Y(top_core_KE_n2145) );
  INVX1 U23494 ( .A(top_core_KE_new_sboxw_192_0_), .Y(n6767) );
  OAI221XL U23495 ( .A0(top_core_KE_n2142), .A1(n2236), .B0(n2244), .B1(n6974), 
        .C0(top_core_KE_n2143), .Y(top_core_KE_n4782) );
  AOI222X1 U23496 ( .A0(n2254), .A1(n1803), .B0(n2264), .B1(
        top_core_KE_CipherKey0_137_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_73_), .Y(top_core_KE_n2143) );
  XNOR2X1 U23497 ( .A(top_core_KE_n2144), .B(n6764), .Y(top_core_KE_n2142) );
  INVX1 U23498 ( .A(top_core_KE_new_sboxw_192_1_), .Y(n6764) );
  OAI221XL U23499 ( .A0(top_core_KE_n2160), .A1(n2236), .B0(n2244), .B1(n6932), 
        .C0(top_core_KE_n2161), .Y(top_core_KE_n4788) );
  AOI222X1 U23500 ( .A0(n2254), .A1(n1348), .B0(n2264), .B1(
        top_core_KE_CipherKey0_131_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_67_), .Y(top_core_KE_n2161) );
  XNOR2X1 U23501 ( .A(top_core_KE_n2162), .B(n6420), .Y(top_core_KE_n2160) );
  INVX1 U23502 ( .A(top_core_KE_new_sboxw_192_27_), .Y(n6420) );
  OAI221XL U23503 ( .A0(top_core_KE_n2157), .A1(n2236), .B0(n2244), .B1(n6856), 
        .C0(top_core_KE_n2158), .Y(top_core_KE_n4787) );
  AOI222X1 U23504 ( .A0(n2254), .A1(n1352), .B0(n2264), .B1(
        top_core_KE_CipherKey0_132_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_68_), .Y(top_core_KE_n2158) );
  XNOR2X1 U23505 ( .A(top_core_KE_n2159), .B(n6413), .Y(top_core_KE_n2157) );
  INVX1 U23506 ( .A(top_core_KE_new_sboxw_192_28_), .Y(n6413) );
  OAI221XL U23507 ( .A0(top_core_KE_n2154), .A1(n2236), .B0(n2244), .B1(n6784), 
        .C0(top_core_KE_n2155), .Y(top_core_KE_n4786) );
  AOI222X1 U23508 ( .A0(n2254), .A1(n1822), .B0(n2264), .B1(
        top_core_KE_CipherKey0_133_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_69_), .Y(top_core_KE_n2155) );
  XNOR2X1 U23509 ( .A(top_core_KE_n2156), .B(n6410), .Y(top_core_KE_n2154) );
  INVX1 U23510 ( .A(top_core_KE_new_sboxw_192_29_), .Y(n6410) );
  OAI221XL U23511 ( .A0(top_core_KE_n2151), .A1(n2236), .B0(n2244), .B1(n6387), 
        .C0(top_core_KE_n2152), .Y(top_core_KE_n4785) );
  AOI222X1 U23512 ( .A0(n2254), .A1(n1343), .B0(n2264), .B1(
        top_core_KE_CipherKey0_134_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_70_), .Y(top_core_KE_n2152) );
  XNOR2X1 U23513 ( .A(top_core_KE_n2153), .B(n6409), .Y(top_core_KE_n2151) );
  INVX1 U23514 ( .A(top_core_KE_new_sboxw_192_30_), .Y(n6409) );
  OAI221XL U23515 ( .A0(top_core_KE_n2100), .A1(n2238), .B0(n2246), .B1(n6991), 
        .C0(top_core_KE_n2101), .Y(top_core_KE_n4768) );
  AOI222X1 U23516 ( .A0(n2260), .A1(n1339), .B0(top_core_KE_n1876), .B1(
        top_core_KE_CipherKey0_151_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_87_), .Y(top_core_KE_n2101) );
  XNOR2X1 U23517 ( .A(top_core_KE_n2102), .B(n6708), .Y(top_core_KE_n2100) );
  INVX1 U23518 ( .A(top_core_KE_new_sboxw_192_15_), .Y(n6708) );
  OAI221XL U23519 ( .A0(top_core_KE_n2169), .A1(n2236), .B0(n2244), .B1(n6979), 
        .C0(top_core_KE_n2170), .Y(top_core_KE_n4791) );
  AOI222X1 U23520 ( .A0(n2254), .A1(n1831), .B0(n2264), .B1(
        top_core_KE_CipherKey0_128_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_64_), .Y(top_core_KE_n2170) );
  XNOR2X1 U23521 ( .A(top_core_KE_n2171), .B(n6427), .Y(top_core_KE_n2169) );
  INVX1 U23522 ( .A(top_core_KE_new_sboxw_192_24_), .Y(n6427) );
  OAI221XL U23523 ( .A0(top_core_KE_n2166), .A1(n2236), .B0(n2244), .B1(n6969), 
        .C0(top_core_KE_n2167), .Y(top_core_KE_n4790) );
  AOI222X1 U23524 ( .A0(n2254), .A1(n1824), .B0(n2264), .B1(
        top_core_KE_CipherKey0_129_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_65_), .Y(top_core_KE_n2167) );
  XNOR2X1 U23525 ( .A(top_core_KE_n2168), .B(n6424), .Y(top_core_KE_n2166) );
  INVX1 U23526 ( .A(top_core_KE_new_sboxw_192_25_), .Y(n6424) );
  OAI221XL U23527 ( .A0(top_core_KE_n2139), .A1(n2236), .B0(n2244), .B1(n6963), 
        .C0(top_core_KE_n2140), .Y(top_core_KE_n4781) );
  AOI222X1 U23528 ( .A0(n2254), .A1(n1344), .B0(n2264), .B1(
        top_core_KE_CipherKey0_138_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_74_), .Y(top_core_KE_n2140) );
  XNOR2X1 U23529 ( .A(top_core_KE_n2141), .B(n6760), .Y(top_core_KE_n2139) );
  INVX1 U23530 ( .A(top_core_KE_new_sboxw_192_2_), .Y(n6760) );
  OAI221XL U23531 ( .A0(top_core_KE_n2163), .A1(n2236), .B0(n2244), .B1(n6957), 
        .C0(top_core_KE_n2164), .Y(top_core_KE_n4789) );
  AOI222X1 U23532 ( .A0(n2254), .A1(n1345), .B0(n2264), .B1(
        top_core_KE_CipherKey0_130_), .C0(n2274), .C1(
        top_core_KE_CipherKey0_66_), .Y(top_core_KE_n2164) );
  XNOR2X1 U23533 ( .A(top_core_KE_n2165), .B(n6416), .Y(top_core_KE_n2163) );
  INVX1 U23534 ( .A(top_core_KE_new_sboxw_192_26_), .Y(n6416) );
  OAI221XL U23535 ( .A0(top_core_KE_n2136), .A1(n2237), .B0(n2245), .B1(n6947), 
        .C0(top_core_KE_n2137), .Y(top_core_KE_n4780) );
  AOI222X1 U23536 ( .A0(n2255), .A1(n1346), .B0(n2268), .B1(
        top_core_KE_CipherKey0_139_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_75_), .Y(top_core_KE_n2137) );
  XNOR2X1 U23537 ( .A(top_core_KE_n2138), .B(n6757), .Y(top_core_KE_n2136) );
  INVX1 U23538 ( .A(top_core_KE_new_sboxw_192_3_), .Y(n6757) );
  OAI221XL U23539 ( .A0(top_core_KE_n2133), .A1(n2237), .B0(n2245), .B1(n6902), 
        .C0(top_core_KE_n2134), .Y(top_core_KE_n4779) );
  AOI222X1 U23540 ( .A0(n2255), .A1(n1350), .B0(n2264), .B1(
        top_core_KE_CipherKey0_140_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_76_), .Y(top_core_KE_n2134) );
  XNOR2X1 U23541 ( .A(top_core_KE_n2135), .B(n6754), .Y(top_core_KE_n2133) );
  INVX1 U23542 ( .A(top_core_KE_new_sboxw_192_4_), .Y(n6754) );
  OAI221XL U23543 ( .A0(top_core_KE_n2130), .A1(n2237), .B0(n2245), .B1(n6822), 
        .C0(top_core_KE_n2131), .Y(top_core_KE_n4778) );
  AOI222X1 U23544 ( .A0(n2255), .A1(n1801), .B0(n2266), .B1(
        top_core_KE_CipherKey0_141_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_77_), .Y(top_core_KE_n2131) );
  XNOR2X1 U23545 ( .A(top_core_KE_n2132), .B(n6751), .Y(top_core_KE_n2130) );
  INVX1 U23546 ( .A(top_core_KE_new_sboxw_192_5_), .Y(n6751) );
  OAI221XL U23547 ( .A0(top_core_KE_n2127), .A1(n2237), .B0(n2245), .B1(n6720), 
        .C0(top_core_KE_n2128), .Y(top_core_KE_n4777) );
  AOI222X1 U23548 ( .A0(n2255), .A1(n1354), .B0(n2267), .B1(
        top_core_KE_CipherKey0_142_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_78_), .Y(top_core_KE_n2128) );
  XNOR2X1 U23549 ( .A(top_core_KE_n2129), .B(n6750), .Y(top_core_KE_n2127) );
  INVX1 U23550 ( .A(top_core_KE_new_sboxw_192_6_), .Y(n6750) );
  OAI221XL U23551 ( .A0(top_core_KE_n2097), .A1(n2238), .B0(n2245), .B1(n6697), 
        .C0(top_core_KE_n2098), .Y(top_core_KE_n4767) );
  AOI222X1 U23552 ( .A0(n2261), .A1(n1768), .B0(top_core_KE_n1876), .B1(
        top_core_KE_CipherKey0_152_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_88_), .Y(top_core_KE_n2098) );
  XNOR2X1 U23553 ( .A(top_core_KE_n2099), .B(n6466), .Y(top_core_KE_n2097) );
  OAI221XL U23554 ( .A0(top_core_KE_n2121), .A1(n2237), .B0(n2245), .B1(n6691), 
        .C0(top_core_KE_n2122), .Y(top_core_KE_n4775) );
  AOI222X1 U23555 ( .A0(n2255), .A1(n1789), .B0(n2271), .B1(
        top_core_KE_CipherKey0_144_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_80_), .Y(top_core_KE_n2122) );
  XNOR2X1 U23556 ( .A(top_core_KE_n2123), .B(n6710), .Y(top_core_KE_n2121) );
  INVX1 U23557 ( .A(top_core_KE_new_sboxw_192_8_), .Y(n6710) );
  OAI221XL U23558 ( .A0(top_core_KE_n2118), .A1(n2237), .B0(n2245), .B1(n6684), 
        .C0(top_core_KE_n2119), .Y(top_core_KE_n4774) );
  AOI222X1 U23559 ( .A0(n2255), .A1(n1782), .B0(n2268), .B1(
        top_core_KE_CipherKey0_145_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_81_), .Y(top_core_KE_n2119) );
  XNOR2X1 U23560 ( .A(top_core_KE_n2120), .B(n6709), .Y(top_core_KE_n2118) );
  INVX1 U23561 ( .A(top_core_KE_new_sboxw_192_9_), .Y(n6709) );
  OAI221XL U23562 ( .A0(top_core_KE_n2091), .A1(n2238), .B0(n2249), .B1(n6676), 
        .C0(top_core_KE_n2092), .Y(top_core_KE_n4765) );
  AOI222X1 U23563 ( .A0(n2254), .A1(n1358), .B0(top_core_KE_n1876), .B1(
        top_core_KE_CipherKey0_154_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_90_), .Y(top_core_KE_n2092) );
  XNOR2X1 U23564 ( .A(top_core_KE_n2093), .B(n6461), .Y(top_core_KE_n2091) );
  OAI221XL U23565 ( .A0(top_core_KE_n2115), .A1(n2237), .B0(n2245), .B1(n6669), 
        .C0(top_core_KE_n2116), .Y(top_core_KE_n4773) );
  AOI222X1 U23566 ( .A0(n2255), .A1(n1359), .B0(n2265), .B1(
        top_core_KE_CipherKey0_146_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_82_), .Y(top_core_KE_n2116) );
  XNOR2X1 U23567 ( .A(top_core_KE_n2117), .B(n6705), .Y(top_core_KE_n2115) );
  INVX1 U23568 ( .A(top_core_KE_new_sboxw_192_10_), .Y(n6705) );
  OAI221XL U23569 ( .A0(top_core_KE_n2088), .A1(n2238), .B0(n2247), .B1(n6657), 
        .C0(top_core_KE_n2089), .Y(top_core_KE_n4764) );
  AOI222X1 U23570 ( .A0(n2257), .A1(n1360), .B0(n2265), .B1(
        top_core_KE_CipherKey0_155_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_91_), .Y(top_core_KE_n2089) );
  XNOR2X1 U23571 ( .A(top_core_KE_n2090), .B(n6458), .Y(top_core_KE_n2088) );
  OAI221XL U23572 ( .A0(top_core_KE_n2112), .A1(n2237), .B0(n2245), .B1(n6641), 
        .C0(top_core_KE_n2113), .Y(top_core_KE_n4772) );
  AOI222X1 U23573 ( .A0(n2255), .A1(n1362), .B0(n2270), .B1(
        top_core_KE_CipherKey0_147_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_83_), .Y(top_core_KE_n2113) );
  XNOR2X1 U23574 ( .A(top_core_KE_n2114), .B(n6707), .Y(top_core_KE_n2112) );
  INVX1 U23575 ( .A(top_core_KE_new_sboxw_192_11_), .Y(n6707) );
  OAI221XL U23576 ( .A0(top_core_KE_n2085), .A1(n2238), .B0(n2251), .B1(n6609), 
        .C0(top_core_KE_n2086), .Y(top_core_KE_n4763) );
  AOI222X1 U23577 ( .A0(n2255), .A1(n1364), .B0(top_core_KE_n1876), .B1(
        top_core_KE_CipherKey0_156_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_92_), .Y(top_core_KE_n2086) );
  XNOR2X1 U23578 ( .A(top_core_KE_n2087), .B(n6455), .Y(top_core_KE_n2085) );
  OAI221XL U23579 ( .A0(top_core_KE_n2109), .A1(n2237), .B0(n2245), .B1(n6562), 
        .C0(top_core_KE_n2110), .Y(top_core_KE_n4771) );
  AOI222X1 U23580 ( .A0(n2255), .A1(n1366), .B0(n2269), .B1(
        top_core_KE_CipherKey0_148_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_84_), .Y(top_core_KE_n2110) );
  XNOR2X1 U23581 ( .A(top_core_KE_n2111), .B(n6704), .Y(top_core_KE_n2109) );
  INVX1 U23582 ( .A(top_core_KE_new_sboxw_192_12_), .Y(n6704) );
  OAI221XL U23583 ( .A0(top_core_KE_n2082), .A1(n2238), .B0(n2246), .B1(n6526), 
        .C0(top_core_KE_n2083), .Y(top_core_KE_n4762) );
  AOI222X1 U23584 ( .A0(n2258), .A1(n1755), .B0(n2270), .B1(
        top_core_KE_CipherKey0_157_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_93_), .Y(top_core_KE_n2083) );
  XNOR2X1 U23585 ( .A(top_core_KE_n2084), .B(n6452), .Y(top_core_KE_n2082) );
  OAI221XL U23586 ( .A0(top_core_KE_n2106), .A1(n2237), .B0(n2245), .B1(n6482), 
        .C0(top_core_KE_n2107), .Y(top_core_KE_n4770) );
  AOI222X1 U23587 ( .A0(n2255), .A1(n1780), .B0(n2264), .B1(
        top_core_KE_CipherKey0_149_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_85_), .Y(top_core_KE_n2107) );
  XNOR2X1 U23588 ( .A(top_core_KE_n2108), .B(n6703), .Y(top_core_KE_n2106) );
  INVX1 U23589 ( .A(top_core_KE_new_sboxw_192_13_), .Y(n6703) );
  OAI221XL U23590 ( .A0(top_core_KE_n2079), .A1(n2238), .B0(n2245), .B1(n6438), 
        .C0(top_core_KE_n2080), .Y(top_core_KE_n4761) );
  AOI222X1 U23591 ( .A0(n2259), .A1(n1368), .B0(top_core_KE_n1876), .B1(
        top_core_KE_CipherKey0_158_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_94_), .Y(top_core_KE_n2080) );
  XNOR2X1 U23592 ( .A(top_core_KE_n2081), .B(n6449), .Y(top_core_KE_n2079) );
  OAI221XL U23593 ( .A0(top_core_KE_n2103), .A1(n2237), .B0(n2245), .B1(n6404), 
        .C0(top_core_KE_n2104), .Y(top_core_KE_n4769) );
  AOI222X1 U23594 ( .A0(n2255), .A1(n1357), .B0(n2266), .B1(
        top_core_KE_CipherKey0_150_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_86_), .Y(top_core_KE_n2104) );
  XNOR2X1 U23595 ( .A(top_core_KE_n2105), .B(n6702), .Y(top_core_KE_n2103) );
  INVX1 U23596 ( .A(top_core_KE_new_sboxw_192_14_), .Y(n6702) );
  OAI221XL U23597 ( .A0(top_core_KE_n2076), .A1(n2238), .B0(n2250), .B1(n6345), 
        .C0(top_core_KE_n2077), .Y(top_core_KE_n4760) );
  AOI222X1 U23598 ( .A0(n2256), .A1(n1370), .B0(n2269), .B1(
        top_core_KE_CipherKey0_159_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_95_), .Y(top_core_KE_n2077) );
  XNOR2X1 U23599 ( .A(top_core_KE_n2078), .B(n6448), .Y(top_core_KE_n2076) );
  OAI221XL U23600 ( .A0(top_core_KE_n2124), .A1(n2237), .B0(n2245), .B1(n6331), 
        .C0(top_core_KE_n2125), .Y(top_core_KE_n4776) );
  AOI222X1 U23601 ( .A0(n2255), .A1(n1338), .B0(n2267), .B1(
        top_core_KE_CipherKey0_143_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_79_), .Y(top_core_KE_n2125) );
  XNOR2X1 U23602 ( .A(top_core_KE_n2126), .B(n6749), .Y(top_core_KE_n2124) );
  INVX1 U23603 ( .A(top_core_KE_new_sboxw_192_7_), .Y(n6749) );
  OAI221XL U23604 ( .A0(top_core_KE_n2094), .A1(n2238), .B0(n2248), .B1(n6318), 
        .C0(top_core_KE_n2095), .Y(top_core_KE_n4766) );
  AOI222X1 U23605 ( .A0(n2260), .A1(n1761), .B0(n2264), .B1(
        top_core_KE_CipherKey0_153_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_89_), .Y(top_core_KE_n2095) );
  XNOR2X1 U23606 ( .A(top_core_KE_n2096), .B(n6463), .Y(top_core_KE_n2094) );
  OAI221XL U23607 ( .A0(top_core_KE_n1629), .A1(n2349), .B0(n2288), .B1(n1753), 
        .C0(top_core_KE_n2568), .Y(top_core_KE_n4890) );
  AOI222X1 U23608 ( .A0(n2342), .A1(top_core_KE_n1633), .B0(n2323), .B1(
        top_core_KE_CipherKey0_29_), .C0(n2332), .C1(top_core_KE_n1631), .Y(
        top_core_KE_n2568) );
  OAI221XL U23609 ( .A0(top_core_KE_n1773), .A1(n2347), .B0(n2290), .B1(n1209), 
        .C0(top_core_KE_n2646), .Y(top_core_KE_n4908) );
  AOI222X1 U23610 ( .A0(n2343), .A1(top_core_KE_n1777), .B0(n2324), .B1(
        top_core_KE_CipherKey0_11_), .C0(n2333), .C1(top_core_KE_n1775), .Y(
        top_core_KE_n2646) );
  OAI221XL U23611 ( .A0(top_core_KE_n1837), .A1(n2347), .B0(n2290), .B1(n1207), 
        .C0(top_core_KE_n2678), .Y(top_core_KE_n4916) );
  AOI222X1 U23612 ( .A0(n2344), .A1(top_core_KE_n1841), .B0(n2320), .B1(
        top_core_KE_CipherKey0_3_), .C0(n2334), .C1(top_core_KE_n1839), .Y(
        top_core_KE_n2678) );
  OAI221XL U23613 ( .A0(top_core_KE_n1709), .A1(n2348), .B0(n2289), .B1(n1167), 
        .C0(top_core_KE_n2614), .Y(top_core_KE_n4900) );
  AOI222X1 U23614 ( .A0(n2343), .A1(top_core_KE_n1713), .B0(n2324), .B1(
        top_core_KE_CipherKey0_19_), .C0(n2333), .C1(top_core_KE_n1711), .Y(
        top_core_KE_n2614) );
  OAI221XL U23615 ( .A0(top_core_KE_n1781), .A1(n2347), .B0(n2290), .B1(n1211), 
        .C0(top_core_KE_n2650), .Y(top_core_KE_n4909) );
  AOI222X1 U23616 ( .A0(n2343), .A1(top_core_KE_n1785), .B0(n2324), .B1(
        top_core_KE_CipherKey0_10_), .C0(n2333), .C1(top_core_KE_n1783), .Y(
        top_core_KE_n2650) );
  OAI221XL U23617 ( .A0(top_core_KE_n1845), .A1(n2347), .B0(n2290), .B1(n1210), 
        .C0(top_core_KE_n2682), .Y(top_core_KE_n4917) );
  AOI222X1 U23618 ( .A0(n2344), .A1(top_core_KE_n1849), .B0(n2319), .B1(
        top_core_KE_CipherKey0_2_), .C0(n2334), .C1(top_core_KE_n1847), .Y(
        top_core_KE_n2682) );
  OAI221XL U23619 ( .A0(top_core_KE_n1717), .A1(n2348), .B0(n2289), .B1(n1170), 
        .C0(top_core_KE_n2618), .Y(top_core_KE_n4901) );
  AOI222X1 U23620 ( .A0(n2343), .A1(top_core_KE_n1721), .B0(n2324), .B1(
        top_core_KE_CipherKey0_18_), .C0(n2333), .C1(top_core_KE_n1719), .Y(
        top_core_KE_n2618) );
  OAI221XL U23621 ( .A0(top_core_KE_n1358), .A1(n2347), .B0(n2305), .B1(n6338), 
        .C0(top_core_KE_n2511), .Y(top_core_KE_n4856) );
  AOI222X1 U23622 ( .A0(n2340), .A1(top_core_KE_n1361), .B0(n2321), .B1(
        top_core_KE_CipherKey0_63_), .C0(n2330), .C1(top_core_KE_n1359), .Y(
        top_core_KE_n2511) );
  OAI221XL U23623 ( .A0(top_core_KE_n1645), .A1(n2349), .B0(n2289), .B1(n1169), 
        .C0(top_core_KE_n2578), .Y(top_core_KE_n4892) );
  AOI222X1 U23624 ( .A0(n2342), .A1(top_core_KE_n1649), .B0(n2323), .B1(
        top_core_KE_CipherKey0_27_), .C0(n2332), .C1(top_core_KE_n1647), .Y(
        top_core_KE_n2578) );
  OAI221XL U23625 ( .A0(top_core_KE_n1813), .A1(n2347), .B0(n2290), .B1(n1224), 
        .C0(top_core_KE_n2666), .Y(top_core_KE_n4913) );
  AOI222X1 U23626 ( .A0(n2343), .A1(top_core_KE_n1817), .B0(n2324), .B1(
        top_core_KE_CipherKey0_6_), .C0(n2333), .C1(top_core_KE_n1815), .Y(
        top_core_KE_n2666) );
  OAI221XL U23627 ( .A0(top_core_KE_n1765), .A1(n2348), .B0(n2290), .B1(n1204), 
        .C0(top_core_KE_n2642), .Y(top_core_KE_n4907) );
  AOI222X1 U23628 ( .A0(n2343), .A1(top_core_KE_n1769), .B0(n2324), .B1(
        top_core_KE_CipherKey0_12_), .C0(n2333), .C1(top_core_KE_n1767), .Y(
        top_core_KE_n2642) );
  OAI221XL U23629 ( .A0(top_core_KE_n1829), .A1(n2347), .B0(n2288), .B1(n1195), 
        .C0(top_core_KE_n2674), .Y(top_core_KE_n4915) );
  AOI222X1 U23630 ( .A0(n2344), .A1(top_core_KE_n1833), .B0(n2317), .B1(
        top_core_KE_CipherKey0_4_), .C0(n2334), .C1(top_core_KE_n1831), .Y(
        top_core_KE_n2674) );
  OAI221XL U23631 ( .A0(top_core_KE_n1749), .A1(n2348), .B0(n2290), .B1(n1187), 
        .C0(top_core_KE_n2634), .Y(top_core_KE_n4905) );
  AOI222X1 U23632 ( .A0(n2343), .A1(top_core_KE_n1753), .B0(n2324), .B1(
        top_core_KE_CipherKey0_14_), .C0(n2333), .C1(top_core_KE_n1751), .Y(
        top_core_KE_n2634) );
  OAI221XL U23633 ( .A0(top_core_KE_n1685), .A1(n2348), .B0(n2289), .B1(n1184), 
        .C0(top_core_KE_n2602), .Y(top_core_KE_n4897) );
  AOI222X1 U23634 ( .A0(n2342), .A1(top_core_KE_n1689), .B0(n2323), .B1(
        top_core_KE_CipherKey0_22_), .C0(n2332), .C1(top_core_KE_n1687), .Y(
        top_core_KE_n2602) );
  OAI221XL U23635 ( .A0(top_core_KE_n1701), .A1(n2348), .B0(n2289), .B1(n1155), 
        .C0(top_core_KE_n2610), .Y(top_core_KE_n4899) );
  AOI222X1 U23636 ( .A0(n2343), .A1(top_core_KE_n1705), .B0(n2324), .B1(
        top_core_KE_CipherKey0_20_), .C0(n2333), .C1(top_core_KE_n1703), .Y(
        top_core_KE_n2610) );
  OAI221XL U23637 ( .A0(top_core_KE_n1637), .A1(n2349), .B0(n2288), .B1(n1164), 
        .C0(top_core_KE_n2573), .Y(top_core_KE_n4891) );
  AOI222X1 U23638 ( .A0(n2342), .A1(top_core_KE_n1641), .B0(n2323), .B1(
        top_core_KE_CipherKey0_28_), .C0(n2332), .C1(top_core_KE_n1639), .Y(
        top_core_KE_n2573) );
  OAI221XL U23639 ( .A0(top_core_KE_n1621), .A1(n2349), .B0(n2288), .B1(n1147), 
        .C0(top_core_KE_n2563), .Y(top_core_KE_n4889) );
  AOI222X1 U23640 ( .A0(n2342), .A1(top_core_KE_n1625), .B0(n2323), .B1(
        top_core_KE_CipherKey0_30_), .C0(n2332), .C1(top_core_KE_n1623), .Y(
        top_core_KE_n2563) );
  OAI221XL U23641 ( .A0(top_core_KE_n1413), .A1(n2347), .B0(n2305), .B1(n6693), 
        .C0(top_core_KE_n2531), .Y(top_core_KE_n4863) );
  INVX1 U23642 ( .A(top_core_KE_prev_key1_reg_56_), .Y(n6693) );
  AOI222X1 U23643 ( .A0(n2340), .A1(top_core_KE_n1417), .B0(n2321), .B1(
        top_core_KE_CipherKey0_56_), .C0(n2330), .C1(top_core_KE_n1415), .Y(
        top_core_KE_n2531) );
  OAI221XL U23644 ( .A0(top_core_KE_n1397), .A1(n2348), .B0(n2305), .B1(n6672), 
        .C0(top_core_KE_n2525), .Y(top_core_KE_n4861) );
  INVX1 U23645 ( .A(top_core_KE_prev_key1_reg_58_), .Y(n6672) );
  AOI222X1 U23646 ( .A0(n2340), .A1(top_core_KE_n1401), .B0(n2321), .B1(
        top_core_KE_CipherKey0_58_), .C0(n2330), .C1(top_core_KE_n1399), .Y(
        top_core_KE_n2525) );
  OAI221XL U23647 ( .A0(top_core_KE_n1389), .A1(n2349), .B0(n2287), .B1(n6648), 
        .C0(top_core_KE_n2522), .Y(top_core_KE_n4860) );
  INVX1 U23648 ( .A(top_core_KE_prev_key1_reg_59_), .Y(n6648) );
  AOI222X1 U23649 ( .A0(n2340), .A1(top_core_KE_n1393), .B0(n2321), .B1(
        top_core_KE_CipherKey0_59_), .C0(n2330), .C1(top_core_KE_n1391), .Y(
        top_core_KE_n2522) );
  OAI221XL U23650 ( .A0(top_core_KE_n1381), .A1(n2348), .B0(n2287), .B1(n6584), 
        .C0(top_core_KE_n2519), .Y(top_core_KE_n4859) );
  INVX1 U23651 ( .A(top_core_KE_prev_key1_reg_60_), .Y(n6584) );
  AOI222X1 U23652 ( .A0(n2340), .A1(top_core_KE_n1385), .B0(n2321), .B1(
        top_core_KE_CipherKey0_60_), .C0(n2330), .C1(top_core_KE_n1383), .Y(
        top_core_KE_n2519) );
  OAI221XL U23653 ( .A0(top_core_KE_n1373), .A1(n2349), .B0(n2288), .B1(n6514), 
        .C0(top_core_KE_n2516), .Y(top_core_KE_n4858) );
  INVX1 U23654 ( .A(top_core_KE_prev_key1_reg_61_), .Y(n6514) );
  AOI222X1 U23655 ( .A0(n2340), .A1(top_core_KE_n1377), .B0(n2321), .B1(
        top_core_KE_CipherKey0_61_), .C0(n2330), .C1(top_core_KE_n1375), .Y(
        top_core_KE_n2516) );
  OAI221XL U23656 ( .A0(top_core_KE_n1365), .A1(n2350), .B0(n2287), .B1(n6406), 
        .C0(top_core_KE_n2513), .Y(top_core_KE_n4857) );
  INVX1 U23657 ( .A(top_core_KE_prev_key1_reg_62_), .Y(n6406) );
  AOI222X1 U23658 ( .A0(n2340), .A1(top_core_KE_n1369), .B0(n2321), .B1(
        top_core_KE_CipherKey0_62_), .C0(n2330), .C1(top_core_KE_n1367), .Y(
        top_core_KE_n2513) );
  OAI221XL U23659 ( .A0(top_core_KE_n1405), .A1(n2350), .B0(n2290), .B1(n6311), 
        .C0(top_core_KE_n2528), .Y(top_core_KE_n4862) );
  INVX1 U23660 ( .A(top_core_KE_prev_key1_reg_57_), .Y(n6311) );
  AOI222X1 U23661 ( .A0(n2340), .A1(top_core_KE_n1409), .B0(n2321), .B1(
        top_core_KE_CipherKey0_57_), .C0(n2330), .C1(top_core_KE_n1407), .Y(
        top_core_KE_n2528) );
  OAI221XL U23662 ( .A0(n6313), .A1(n2242), .B0(n2250), .B1(n6998), .C0(
        top_core_KE_n1920), .Y(top_core_KE_n4702) );
  INVX1 U23663 ( .A(top_core_KE_n1666), .Y(n6313) );
  INVX1 U23664 ( .A(top_core_KE_prev_key0_reg_89_), .Y(n6998) );
  AOI222X1 U23665 ( .A0(n2260), .A1(n1652), .B0(n2269), .B1(
        top_core_KE_CipherKey0_217_), .C0(n2281), .C1(
        top_core_KE_CipherKey0_153_), .Y(top_core_KE_n1920) );
  OAI221XL U23666 ( .A0(top_core_KE_n1661), .A1(n2349), .B0(n2289), .B1(n1765), 
        .C0(top_core_KE_n2588), .Y(top_core_KE_n4894) );
  AOI222X1 U23667 ( .A0(n2342), .A1(top_core_KE_n1665), .B0(n2323), .B1(
        top_core_KE_CipherKey0_25_), .C0(n2332), .C1(top_core_KE_n1663), .Y(
        top_core_KE_n2588) );
  OAI221XL U23668 ( .A0(top_core_KE_n1797), .A1(n2347), .B0(n2290), .B1(n1813), 
        .C0(top_core_KE_n2658), .Y(top_core_KE_n4911) );
  AOI222X1 U23669 ( .A0(n2343), .A1(top_core_KE_n1801), .B0(n2324), .B1(
        top_core_KE_CipherKey0_8_), .C0(n2333), .C1(top_core_KE_n1799), .Y(
        top_core_KE_n2658) );
  OAI221XL U23670 ( .A0(top_core_KE_n1541), .A1(n2350), .B0(n2287), .B1(n6981), 
        .C0(top_core_KE_n2549), .Y(top_core_KE_n4879) );
  INVX1 U23671 ( .A(top_core_KE_prev_key1_reg_40_), .Y(n6981) );
  AOI222X1 U23672 ( .A0(n2341), .A1(top_core_KE_n1545), .B0(n2322), .B1(
        top_core_KE_CipherKey0_40_), .C0(n2331), .C1(top_core_KE_n1543), .Y(
        top_core_KE_n2549) );
  OAI221XL U23673 ( .A0(top_core_KE_n1605), .A1(n2349), .B0(n2288), .B1(n6976), 
        .C0(top_core_KE_n2557), .Y(top_core_KE_n4887) );
  INVX1 U23674 ( .A(top_core_KE_prev_key1_reg_32_), .Y(n6976) );
  AOI222X1 U23675 ( .A0(n2342), .A1(top_core_KE_n1609), .B0(n2323), .B1(
        top_core_KE_CipherKey0_32_), .C0(n2332), .C1(top_core_KE_n1607), .Y(
        top_core_KE_n2557) );
  OAI221XL U23676 ( .A0(top_core_KE_n1789), .A1(n2347), .B0(n2290), .B1(n1806), 
        .C0(top_core_KE_n2654), .Y(top_core_KE_n4910) );
  AOI222X1 U23677 ( .A0(n2343), .A1(top_core_KE_n1793), .B0(n2324), .B1(
        top_core_KE_CipherKey0_9_), .C0(n2333), .C1(top_core_KE_n1791), .Y(
        top_core_KE_n2654) );
  OAI221XL U23678 ( .A0(top_core_KE_n1533), .A1(n2350), .B0(n2287), .B1(n6971), 
        .C0(top_core_KE_n2548), .Y(top_core_KE_n4878) );
  INVX1 U23679 ( .A(top_core_KE_prev_key1_reg_41_), .Y(n6971) );
  AOI222X1 U23680 ( .A0(n2341), .A1(top_core_KE_n1537), .B0(n2322), .B1(
        top_core_KE_CipherKey0_41_), .C0(n2331), .C1(top_core_KE_n1535), .Y(
        top_core_KE_n2548) );
  OAI221XL U23681 ( .A0(top_core_KE_n1597), .A1(n2349), .B0(n2288), .B1(n6966), 
        .C0(top_core_KE_n2556), .Y(top_core_KE_n4886) );
  INVX1 U23682 ( .A(top_core_KE_prev_key1_reg_33_), .Y(n6966) );
  AOI222X1 U23683 ( .A0(n2342), .A1(top_core_KE_n1601), .B0(n2323), .B1(
        top_core_KE_CipherKey0_33_), .C0(n2332), .C1(top_core_KE_n1599), .Y(
        top_core_KE_n2556) );
  OAI221XL U23684 ( .A0(top_core_KE_n1525), .A1(n2350), .B0(n2287), .B1(n6960), 
        .C0(top_core_KE_n2547), .Y(top_core_KE_n4877) );
  INVX1 U23685 ( .A(top_core_KE_prev_key1_reg_42_), .Y(n6960) );
  AOI222X1 U23686 ( .A0(n2341), .A1(top_core_KE_n1529), .B0(n2322), .B1(
        top_core_KE_CipherKey0_42_), .C0(n2331), .C1(top_core_KE_n1527), .Y(
        top_core_KE_n2547) );
  OAI221XL U23687 ( .A0(top_core_KE_n1589), .A1(n2349), .B0(n2288), .B1(n6954), 
        .C0(top_core_KE_n2555), .Y(top_core_KE_n4885) );
  INVX1 U23688 ( .A(top_core_KE_prev_key1_reg_34_), .Y(n6954) );
  AOI222X1 U23689 ( .A0(n2342), .A1(top_core_KE_n1593), .B0(n2323), .B1(
        top_core_KE_CipherKey0_34_), .C0(n2332), .C1(top_core_KE_n1591), .Y(
        top_core_KE_n2555) );
  OAI221XL U23690 ( .A0(top_core_KE_n1517), .A1(n2350), .B0(n2287), .B1(n6939), 
        .C0(top_core_KE_n2546), .Y(top_core_KE_n4876) );
  INVX1 U23691 ( .A(top_core_KE_prev_key1_reg_43_), .Y(n6939) );
  AOI222X1 U23692 ( .A0(n2341), .A1(top_core_KE_n1521), .B0(n2322), .B1(
        top_core_KE_CipherKey0_43_), .C0(n2331), .C1(top_core_KE_n1519), .Y(
        top_core_KE_n2546) );
  OAI221XL U23693 ( .A0(top_core_KE_n1581), .A1(n2349), .B0(n2288), .B1(n6924), 
        .C0(top_core_KE_n2554), .Y(top_core_KE_n4884) );
  INVX1 U23694 ( .A(top_core_KE_prev_key1_reg_35_), .Y(n6924) );
  AOI222X1 U23695 ( .A0(n2342), .A1(top_core_KE_n1585), .B0(n2323), .B1(
        top_core_KE_CipherKey0_35_), .C0(n2332), .C1(top_core_KE_n1583), .Y(
        top_core_KE_n2554) );
  OAI221XL U23696 ( .A0(top_core_KE_n1509), .A1(n2350), .B0(n2287), .B1(n6878), 
        .C0(top_core_KE_n2545), .Y(top_core_KE_n4875) );
  INVX1 U23697 ( .A(top_core_KE_prev_key1_reg_44_), .Y(n6878) );
  AOI222X1 U23698 ( .A0(n2341), .A1(top_core_KE_n1513), .B0(n2322), .B1(
        top_core_KE_CipherKey0_44_), .C0(n2331), .C1(top_core_KE_n1511), .Y(
        top_core_KE_n2545) );
  OAI221XL U23699 ( .A0(top_core_KE_n1573), .A1(n2350), .B0(n2288), .B1(n6832), 
        .C0(top_core_KE_n2553), .Y(top_core_KE_n4883) );
  INVX1 U23700 ( .A(top_core_KE_prev_key1_reg_36_), .Y(n6832) );
  AOI222X1 U23701 ( .A0(n2342), .A1(top_core_KE_n1577), .B0(n2323), .B1(
        top_core_KE_CipherKey0_36_), .C0(n2332), .C1(top_core_KE_n1575), .Y(
        top_core_KE_n2553) );
  OAI221XL U23702 ( .A0(top_core_KE_n1501), .A1(n2350), .B0(n2287), .B1(n6811), 
        .C0(top_core_KE_n2544), .Y(top_core_KE_n4874) );
  INVX1 U23703 ( .A(top_core_KE_prev_key1_reg_45_), .Y(n6811) );
  AOI222X1 U23704 ( .A0(n2341), .A1(top_core_KE_n1505), .B0(n2322), .B1(
        top_core_KE_CipherKey0_45_), .C0(n2331), .C1(top_core_KE_n1503), .Y(
        top_core_KE_n2544) );
  OAI221XL U23705 ( .A0(top_core_KE_n1565), .A1(n2350), .B0(n2288), .B1(n6748), 
        .C0(top_core_KE_n2552), .Y(top_core_KE_n4882) );
  INVX1 U23706 ( .A(top_core_KE_prev_key1_reg_37_), .Y(n6748) );
  AOI222X1 U23707 ( .A0(n2341), .A1(top_core_KE_n1569), .B0(n2322), .B1(
        top_core_KE_CipherKey0_37_), .C0(n2331), .C1(top_core_KE_n1567), .Y(
        top_core_KE_n2552) );
  OAI221XL U23708 ( .A0(top_core_KE_n1669), .A1(n2349), .B0(n2289), .B1(n1772), 
        .C0(top_core_KE_n2593), .Y(top_core_KE_n4895) );
  AOI222X1 U23709 ( .A0(n2342), .A1(top_core_KE_n1673), .B0(n2323), .B1(
        top_core_KE_CipherKey0_24_), .C0(n2332), .C1(top_core_KE_n1671), .Y(
        top_core_KE_n2593) );
  OAI221XL U23710 ( .A0(n6465), .A1(n2242), .B0(n2250), .B1(n6694), .C0(
        top_core_KE_n1922), .Y(top_core_KE_n4703) );
  INVX1 U23711 ( .A(top_core_KE_n1674), .Y(n6465) );
  INVX1 U23712 ( .A(top_core_KE_prev_key0_reg_88_), .Y(n6694) );
  AOI222X1 U23713 ( .A0(n2260), .A1(n1659), .B0(n2269), .B1(
        top_core_KE_CipherKey0_216_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_152_), .Y(top_core_KE_n1922) );
  OAI221XL U23714 ( .A0(top_core_KE_n1733), .A1(n2348), .B0(n2289), .B1(n1792), 
        .C0(top_core_KE_n2626), .Y(top_core_KE_n4903) );
  AOI222X1 U23715 ( .A0(n2343), .A1(top_core_KE_n1737), .B0(n2324), .B1(
        top_core_KE_CipherKey0_16_), .C0(n2333), .C1(top_core_KE_n1735), .Y(
        top_core_KE_n2626) );
  OAI221XL U23716 ( .A0(top_core_KE_n1477), .A1(n2347), .B0(n2288), .B1(n6686), 
        .C0(top_core_KE_n2541), .Y(top_core_KE_n4871) );
  INVX1 U23717 ( .A(top_core_KE_prev_key1_reg_48_), .Y(n6686) );
  AOI222X1 U23718 ( .A0(n2341), .A1(top_core_KE_n1481), .B0(n2322), .B1(
        top_core_KE_CipherKey0_48_), .C0(n2331), .C1(top_core_KE_n1479), .Y(
        top_core_KE_n2541) );
  OAI221XL U23719 ( .A0(top_core_KE_n1725), .A1(n2348), .B0(n2289), .B1(n1785), 
        .C0(top_core_KE_n2622), .Y(top_core_KE_n4902) );
  AOI222X1 U23720 ( .A0(n2343), .A1(top_core_KE_n1729), .B0(n2324), .B1(
        top_core_KE_CipherKey0_17_), .C0(n2333), .C1(top_core_KE_n1727), .Y(
        top_core_KE_n2622) );
  OAI221XL U23721 ( .A0(top_core_KE_n1469), .A1(n2348), .B0(n2287), .B1(n6679), 
        .C0(top_core_KE_n2540), .Y(top_core_KE_n4870) );
  INVX1 U23722 ( .A(top_core_KE_prev_key1_reg_49_), .Y(n6679) );
  AOI222X1 U23723 ( .A0(n2341), .A1(top_core_KE_n1473), .B0(n2322), .B1(
        top_core_KE_CipherKey0_49_), .C0(n2331), .C1(top_core_KE_n1471), .Y(
        top_core_KE_n2540) );
  OAI221XL U23724 ( .A0(n6460), .A1(n2242), .B0(n2250), .B1(n6673), .C0(
        top_core_KE_n1918), .Y(top_core_KE_n4701) );
  INVX1 U23725 ( .A(top_core_KE_n1658), .Y(n6460) );
  INVX1 U23726 ( .A(top_core_KE_prev_key0_reg_90_), .Y(n6673) );
  AOI222X1 U23727 ( .A0(n2260), .A1(n1646), .B0(n2269), .B1(
        top_core_KE_CipherKey0_218_), .C0(n2275), .C1(
        top_core_KE_CipherKey0_154_), .Y(top_core_KE_n1918) );
  OAI221XL U23728 ( .A0(top_core_KE_n1461), .A1(n2349), .B0(n2287), .B1(n6664), 
        .C0(top_core_KE_n2539), .Y(top_core_KE_n4869) );
  INVX1 U23729 ( .A(top_core_KE_prev_key1_reg_50_), .Y(n6664) );
  AOI222X1 U23730 ( .A0(n2341), .A1(top_core_KE_n1465), .B0(n2322), .B1(
        top_core_KE_CipherKey0_50_), .C0(n2331), .C1(top_core_KE_n1463), .Y(
        top_core_KE_n2539) );
  OAI221XL U23731 ( .A0(n6457), .A1(n2242), .B0(n2250), .B1(n6649), .C0(
        top_core_KE_n1916), .Y(top_core_KE_n4700) );
  INVX1 U23732 ( .A(top_core_KE_n1650), .Y(n6457) );
  INVX1 U23733 ( .A(top_core_KE_prev_key0_reg_91_), .Y(n6649) );
  AOI222X1 U23734 ( .A0(n2260), .A1(n1361), .B0(n2269), .B1(
        top_core_KE_CipherKey0_219_), .C0(n2279), .C1(
        top_core_KE_CipherKey0_155_), .Y(top_core_KE_n1916) );
  OAI221XL U23735 ( .A0(top_core_KE_n1453), .A1(n2350), .B0(n2287), .B1(n6631), 
        .C0(top_core_KE_n2538), .Y(top_core_KE_n4868) );
  INVX1 U23736 ( .A(top_core_KE_prev_key1_reg_51_), .Y(n6631) );
  AOI222X1 U23737 ( .A0(n2341), .A1(top_core_KE_n1457), .B0(n2322), .B1(
        top_core_KE_CipherKey0_51_), .C0(n2331), .C1(top_core_KE_n1455), .Y(
        top_core_KE_n2538) );
  OAI221XL U23738 ( .A0(n6454), .A1(n2242), .B0(n2250), .B1(n6585), .C0(
        top_core_KE_n1914), .Y(top_core_KE_n4699) );
  INVX1 U23739 ( .A(top_core_KE_n1642), .Y(n6454) );
  INVX1 U23740 ( .A(top_core_KE_prev_key0_reg_92_), .Y(n6585) );
  AOI222X1 U23741 ( .A0(n2260), .A1(n1365), .B0(n2269), .B1(
        top_core_KE_CipherKey0_220_), .C0(n2280), .C1(
        top_core_KE_CipherKey0_156_), .Y(top_core_KE_n1914) );
  OAI221XL U23742 ( .A0(top_core_KE_n1445), .A1(n2347), .B0(n2288), .B1(n6536), 
        .C0(top_core_KE_n2537), .Y(top_core_KE_n4867) );
  INVX1 U23743 ( .A(top_core_KE_prev_key1_reg_52_), .Y(n6536) );
  AOI222X1 U23744 ( .A0(n2341), .A1(top_core_KE_n1449), .B0(n2322), .B1(
        top_core_KE_CipherKey0_52_), .C0(n2331), .C1(top_core_KE_n1447), .Y(
        top_core_KE_n2537) );
  OAI221XL U23745 ( .A0(n6451), .A1(n2242), .B0(n2250), .B1(n6515), .C0(
        top_core_KE_n1912), .Y(top_core_KE_n4698) );
  INVX1 U23746 ( .A(top_core_KE_n1634), .Y(n6451) );
  INVX1 U23747 ( .A(top_core_KE_prev_key0_reg_93_), .Y(n6515) );
  AOI222X1 U23748 ( .A0(n2260), .A1(top_core_KE_prev_key1_reg_93_), .B0(n2269), 
        .B1(top_core_KE_CipherKey0_221_), .C0(n2276), .C1(
        top_core_KE_CipherKey0_157_), .Y(top_core_KE_n1912) );
  OAI221XL U23749 ( .A0(top_core_KE_n1437), .A1(n2348), .B0(n2287), .B1(n6445), 
        .C0(top_core_KE_n2536), .Y(top_core_KE_n4866) );
  INVX1 U23750 ( .A(top_core_KE_prev_key1_reg_53_), .Y(n6445) );
  AOI222X1 U23751 ( .A0(n2340), .A1(top_core_KE_n1441), .B0(n2321), .B1(
        top_core_KE_CipherKey0_53_), .C0(n2330), .C1(top_core_KE_n1439), .Y(
        top_core_KE_n2536) );
  OAI221XL U23752 ( .A0(n6408), .A1(n2242), .B0(n2250), .B1(n6407), .C0(
        top_core_KE_n1910), .Y(top_core_KE_n4697) );
  INVX1 U23753 ( .A(top_core_KE_n1626), .Y(n6408) );
  INVX1 U23754 ( .A(top_core_KE_prev_key0_reg_94_), .Y(n6407) );
  AOI222X1 U23755 ( .A0(n2260), .A1(n1369), .B0(n2269), .B1(
        top_core_KE_CipherKey0_222_), .C0(n2277), .C1(
        top_core_KE_CipherKey0_158_), .Y(top_core_KE_n1910) );
  OAI221XL U23756 ( .A0(top_core_KE_n1429), .A1(n2349), .B0(n2290), .B1(n6397), 
        .C0(top_core_KE_n2535), .Y(top_core_KE_n4865) );
  INVX1 U23757 ( .A(top_core_KE_prev_key1_reg_54_), .Y(n6397) );
  AOI222X1 U23758 ( .A0(n2340), .A1(top_core_KE_n1433), .B0(n2321), .B1(
        top_core_KE_CipherKey0_54_), .C0(n2330), .C1(top_core_KE_n1431), .Y(
        top_core_KE_n2535) );
  OAI221XL U23759 ( .A0(top_core_KE_n1493), .A1(n2350), .B0(n2287), .B1(n6389), 
        .C0(top_core_KE_n2543), .Y(top_core_KE_n4873) );
  INVX1 U23760 ( .A(top_core_KE_prev_key1_reg_46_), .Y(n6389) );
  AOI222X1 U23761 ( .A0(n2341), .A1(top_core_KE_n1497), .B0(n2322), .B1(
        top_core_KE_CipherKey0_46_), .C0(n2331), .C1(top_core_KE_n1495), .Y(
        top_core_KE_n2543) );
  OAI221XL U23762 ( .A0(top_core_KE_n1557), .A1(n2350), .B0(n2288), .B1(n6381), 
        .C0(top_core_KE_n2551), .Y(top_core_KE_n4881) );
  INVX1 U23763 ( .A(top_core_KE_prev_key1_reg_38_), .Y(n6381) );
  AOI222X1 U23764 ( .A0(n2341), .A1(top_core_KE_n1561), .B0(n2322), .B1(
        top_core_KE_CipherKey0_38_), .C0(n2331), .C1(top_core_KE_n1559), .Y(
        top_core_KE_n2551) );
  OAI221XL U23765 ( .A0(n6340), .A1(n2242), .B0(n2246), .B1(n6375), .C0(
        top_core_KE_n1908), .Y(top_core_KE_n4696) );
  INVX1 U23766 ( .A(top_core_KE_n1618), .Y(n6340) );
  INVX1 U23767 ( .A(top_core_KE_prev_key0_reg_95_), .Y(n6375) );
  AOI222X1 U23768 ( .A0(n2258), .A1(n1341), .B0(n2270), .B1(
        top_core_KE_CipherKey0_223_), .C0(n2278), .C1(
        top_core_KE_CipherKey0_159_), .Y(top_core_KE_n1908) );
  OAI221XL U23769 ( .A0(top_core_KE_n1421), .A1(n2350), .B0(n2288), .B1(n6333), 
        .C0(top_core_KE_n2534), .Y(top_core_KE_n4864) );
  INVX1 U23770 ( .A(top_core_KE_prev_key1_reg_55_), .Y(n6333) );
  AOI222X1 U23771 ( .A0(n2340), .A1(top_core_KE_n1425), .B0(n2321), .B1(
        top_core_KE_CipherKey0_55_), .C0(n2330), .C1(top_core_KE_n1423), .Y(
        top_core_KE_n2534) );
  OAI221XL U23772 ( .A0(top_core_KE_n1485), .A1(n2350), .B0(n2287), .B1(n6324), 
        .C0(top_core_KE_n2542), .Y(top_core_KE_n4872) );
  INVX1 U23773 ( .A(top_core_KE_prev_key1_reg_47_), .Y(n6324) );
  AOI222X1 U23774 ( .A0(n2341), .A1(top_core_KE_n1489), .B0(n2322), .B1(
        top_core_KE_CipherKey0_47_), .C0(n2331), .C1(top_core_KE_n1487), .Y(
        top_core_KE_n2542) );
  OAI221XL U23775 ( .A0(top_core_KE_n1549), .A1(n2350), .B0(n2287), .B1(n6320), 
        .C0(top_core_KE_n2550), .Y(top_core_KE_n4880) );
  INVX1 U23776 ( .A(top_core_KE_prev_key1_reg_39_), .Y(n6320) );
  AOI222X1 U23777 ( .A0(n2341), .A1(top_core_KE_n1553), .B0(n2322), .B1(
        top_core_KE_CipherKey0_39_), .C0(n2331), .C1(top_core_KE_n1551), .Y(
        top_core_KE_n2550) );
  OAI221XL U23778 ( .A0(top_core_KE_n1861), .A1(n2347), .B0(n2290), .B1(n1834), 
        .C0(top_core_KE_n2690), .Y(top_core_KE_n4919) );
  AOI222X1 U23779 ( .A0(n2344), .A1(top_core_KE_n1868), .B0(n2318), .B1(
        top_core_KE_CipherKey0_0_), .C0(n2334), .C1(top_core_KE_n1863), .Y(
        top_core_KE_n2690) );
  OAI221XL U23780 ( .A0(top_core_KE_n1853), .A1(n2347), .B0(n2288), .B1(n1827), 
        .C0(top_core_KE_n2686), .Y(top_core_KE_n4918) );
  AOI222X1 U23781 ( .A0(n2344), .A1(top_core_KE_n1857), .B0(n2320), .B1(
        top_core_KE_CipherKey0_1_), .C0(n2334), .C1(top_core_KE_n1855), .Y(
        top_core_KE_n2686) );
  NAND2X1 U23782 ( .A(top_core_KE_n1864), .B(top_core_KE_n728), .Y(
        top_core_KE_n900) );
  NAND3X1 U23783 ( .A(top_core_KE_n875), .B(top_core_KE_n728), .C(n1333), .Y(
        top_core_KE_n880) );
  NAND3X1 U23784 ( .A(top_core_KE_n878), .B(top_core_KE_n728), .C(n1334), .Y(
        top_core_KE_n889) );
  XNOR2X1 U23785 ( .A(top_core_KE_prev_key1_reg_127_), .B(n6989), .Y(
        top_core_KE_n2344) );
  XNOR2X1 U23786 ( .A(top_core_KE_prev_key1_reg_126_), .B(n1146), .Y(
        top_core_KE_n2350) );
  XNOR2X1 U23787 ( .A(top_core_KE_prev_key1_reg_125_), .B(n1635), .Y(
        top_core_KE_n2356) );
  XNOR2X1 U23788 ( .A(top_core_KE_prev_key1_reg_124_), .B(n1159), .Y(
        top_core_KE_n2362) );
  XNOR2X1 U23789 ( .A(top_core_KE_prev_key1_reg_123_), .B(n1168), .Y(
        top_core_KE_n2368) );
  XNOR2X1 U23790 ( .A(top_core_KE_prev_key1_reg_122_), .B(n1643), .Y(
        top_core_KE_n2374) );
  XNOR2X1 U23791 ( .A(top_core_KE_prev_key1_reg_121_), .B(n1653), .Y(
        top_core_KE_n2380) );
  XNOR2X1 U23792 ( .A(top_core_KE_prev_key1_reg_120_), .B(n1664), .Y(
        top_core_KE_n2386) );
  XNOR2X1 U23795 ( .A(top_core_EC_rounds_2_), .B(n3976), .Y(top_core_EC_n1033)
         );
  NAND2X1 U23796 ( .A(top_core_Key[128]), .B(top_core_Core_Full), .Y(
        top_core_EC_n946) );
  NAND3X1 U23797 ( .A(n1333), .B(top_core_KE_n728), .C(top_core_KE_n887), .Y(
        top_core_KE_n891) );
  NAND3X1 U23798 ( .A(top_core_KE_n883), .B(top_core_KE_n728), .C(
        top_core_KE_n884), .Y(top_core_KE_n882) );
  OAI211X1 U23799 ( .A0(top_core_KE_n2725), .A1(n7018), .B0(top_core_KE_n2722), 
        .C0(top_core_KE_n2721), .Y(top_core_KE_n4933) );
  NAND3X1 U23800 ( .A(n7018), .B(n7017), .C(n3687), .Y(top_core_KE_n2722) );
  INVX1 U23801 ( .A(top_core_KE_key_mem_ctrl_reg_0_), .Y(n7018) );
  NOR2X1 U23802 ( .A(n7247), .B(top_core_EC_rounds_3_), .Y(top_core_EC_N577)
         );
  XNOR2X1 U23803 ( .A(top_core_KE_n2600), .B(top_core_KE_n969), .Y(
        top_core_KE_n1425) );
  XNOR2X1 U23804 ( .A(top_core_KE_prev_key1_reg_55_), .B(n1340), .Y(
        top_core_KE_n2600) );
  XNOR2X1 U23805 ( .A(top_core_KE_n2608), .B(top_core_KE_n983), .Y(
        top_core_KE_n1441) );
  XNOR2X1 U23806 ( .A(top_core_KE_prev_key1_reg_53_), .B(n1666), .Y(
        top_core_KE_n2608) );
  XNOR2X1 U23807 ( .A(top_core_KE_n2620), .B(top_core_KE_n1004), .Y(
        top_core_KE_n1465) );
  XNOR2X1 U23808 ( .A(top_core_KE_prev_key1_reg_50_), .B(n1673), .Y(
        top_core_KE_n2620) );
  XNOR2X1 U23809 ( .A(top_core_KE_n2632), .B(top_core_KE_n1025), .Y(
        top_core_KE_n1489) );
  XNOR2X1 U23810 ( .A(top_core_KE_prev_key1_reg_47_), .B(n1337), .Y(
        top_core_KE_n2632) );
  XNOR2X1 U23811 ( .A(top_core_KE_n2640), .B(top_core_KE_n1039), .Y(
        top_core_KE_n1505) );
  XNOR2X1 U23812 ( .A(top_core_KE_prev_key1_reg_45_), .B(n1695), .Y(
        top_core_KE_n2640) );
  XNOR2X1 U23813 ( .A(top_core_KE_n2652), .B(top_core_KE_n1060), .Y(
        top_core_KE_n1529) );
  XNOR2X1 U23814 ( .A(top_core_KE_prev_key1_reg_42_), .B(n1702), .Y(
        top_core_KE_n2652) );
  XNOR2X1 U23815 ( .A(top_core_KE_n2664), .B(top_core_KE_n1081), .Y(
        top_core_KE_n1553) );
  XNOR2X1 U23816 ( .A(top_core_KE_prev_key1_reg_39_), .B(n1336), .Y(
        top_core_KE_n2664) );
  XNOR2X1 U23817 ( .A(top_core_KE_n2672), .B(top_core_KE_n1095), .Y(
        top_core_KE_n1569) );
  XNOR2X1 U23818 ( .A(top_core_KE_prev_key1_reg_37_), .B(n1724), .Y(
        top_core_KE_n2672) );
  XNOR2X1 U23819 ( .A(top_core_KE_n2684), .B(top_core_KE_n1116), .Y(
        top_core_KE_n1593) );
  XNOR2X1 U23820 ( .A(top_core_KE_prev_key1_reg_34_), .B(n1731), .Y(
        top_core_KE_n2684) );
  XNOR2X1 U23821 ( .A(top_core_KE_n2604), .B(top_core_KE_n976), .Y(
        top_core_KE_n1433) );
  XNOR2X1 U23822 ( .A(top_core_KE_prev_key1_reg_54_), .B(n1356), .Y(
        top_core_KE_n2604) );
  XNOR2X1 U23823 ( .A(top_core_KE_n2612), .B(top_core_KE_n990), .Y(
        top_core_KE_n1449) );
  XNOR2X1 U23824 ( .A(top_core_KE_prev_key1_reg_52_), .B(n1367), .Y(
        top_core_KE_n2612) );
  XNOR2X1 U23825 ( .A(top_core_KE_n2616), .B(top_core_KE_n997), .Y(
        top_core_KE_n1457) );
  XNOR2X1 U23826 ( .A(top_core_KE_prev_key1_reg_51_), .B(n1363), .Y(
        top_core_KE_n2616) );
  XNOR2X1 U23827 ( .A(top_core_KE_n2624), .B(top_core_KE_n1011), .Y(
        top_core_KE_n1473) );
  XNOR2X1 U23828 ( .A(top_core_KE_prev_key1_reg_49_), .B(n1680), .Y(
        top_core_KE_n2624) );
  XNOR2X1 U23829 ( .A(top_core_KE_n2628), .B(top_core_KE_n1018), .Y(
        top_core_KE_n1481) );
  XNOR2X1 U23830 ( .A(top_core_KE_prev_key1_reg_48_), .B(n1687), .Y(
        top_core_KE_n2628) );
  XNOR2X1 U23831 ( .A(top_core_KE_n2636), .B(top_core_KE_n1032), .Y(
        top_core_KE_n1497) );
  XNOR2X1 U23832 ( .A(top_core_KE_prev_key1_reg_46_), .B(n1355), .Y(
        top_core_KE_n2636) );
  XNOR2X1 U23833 ( .A(top_core_KE_n2644), .B(top_core_KE_n1046), .Y(
        top_core_KE_n1513) );
  XNOR2X1 U23834 ( .A(top_core_KE_prev_key1_reg_44_), .B(n1351), .Y(
        top_core_KE_n2644) );
  XNOR2X1 U23835 ( .A(top_core_KE_n2648), .B(top_core_KE_n1053), .Y(
        top_core_KE_n1521) );
  XNOR2X1 U23836 ( .A(top_core_KE_prev_key1_reg_43_), .B(n1347), .Y(
        top_core_KE_n2648) );
  XNOR2X1 U23837 ( .A(top_core_KE_n2656), .B(top_core_KE_n1067), .Y(
        top_core_KE_n1537) );
  XNOR2X1 U23838 ( .A(top_core_KE_prev_key1_reg_41_), .B(n1709), .Y(
        top_core_KE_n2656) );
  XNOR2X1 U23839 ( .A(top_core_KE_n2660), .B(top_core_KE_n1074), .Y(
        top_core_KE_n1545) );
  XNOR2X1 U23840 ( .A(top_core_KE_prev_key1_reg_40_), .B(n1716), .Y(
        top_core_KE_n2660) );
  XNOR2X1 U23841 ( .A(top_core_KE_n2668), .B(top_core_KE_n1088), .Y(
        top_core_KE_n1561) );
  XNOR2X1 U23842 ( .A(top_core_KE_prev_key1_reg_38_), .B(n1342), .Y(
        top_core_KE_n2668) );
  XNOR2X1 U23843 ( .A(top_core_KE_n2676), .B(top_core_KE_n1102), .Y(
        top_core_KE_n1577) );
  XNOR2X1 U23844 ( .A(top_core_KE_prev_key1_reg_36_), .B(n1353), .Y(
        top_core_KE_n2676) );
  XNOR2X1 U23845 ( .A(top_core_KE_n2680), .B(top_core_KE_n1109), .Y(
        top_core_KE_n1585) );
  XNOR2X1 U23846 ( .A(top_core_KE_prev_key1_reg_35_), .B(n1349), .Y(
        top_core_KE_n2680) );
  XNOR2X1 U23847 ( .A(top_core_KE_n2688), .B(top_core_KE_n1123), .Y(
        top_core_KE_n1601) );
  XNOR2X1 U23848 ( .A(top_core_KE_prev_key1_reg_33_), .B(n1738), .Y(
        top_core_KE_n2688) );
  XNOR2X1 U23849 ( .A(top_core_KE_n2694), .B(top_core_KE_n1130), .Y(
        top_core_KE_n1609) );
  XNOR2X1 U23850 ( .A(top_core_KE_prev_key1_reg_32_), .B(n1745), .Y(
        top_core_KE_n2694) );
  INVX1 U23851 ( .A(top_core_KE_rcon_reg_7_), .Y(n7006) );
  NAND2X1 U23853 ( .A(top_core_io_inter_ok), .B(top_core_io_NK_0_), .Y(
        top_core_io_n653) );
  NAND3X1 U23854 ( .A(top_core_EC_n863), .B(top_core_EC_n864), .C(
        top_core_EC_n865), .Y(top_core_EC_n861) );
  NOR3X1 U23856 ( .A(top_core_EC_n866), .B(top_core_EC_N577), .C(
        top_core_EC_n867), .Y(top_core_EC_n865) );
  INVX1 U23857 ( .A(top_core_KE_key_mem_ctrl_reg_1_), .Y(n7017) );
  XNOR2X1 U23858 ( .A(top_core_KE_n2601), .B(top_core_KE_n1925), .Y(
        top_core_KE_n2599) );
  XNOR2X1 U23859 ( .A(top_core_KE_prev_key0_reg_23_), .B(
        top_core_KE_prev_key0_reg_55_), .Y(top_core_KE_n2601) );
  XNOR2X1 U23860 ( .A(top_core_KE_n2605), .B(top_core_KE_n1927), .Y(
        top_core_KE_n2603) );
  XNOR2X1 U23861 ( .A(top_core_KE_prev_key0_reg_22_), .B(
        top_core_KE_prev_key0_reg_54_), .Y(top_core_KE_n2605) );
  XNOR2X1 U23862 ( .A(top_core_KE_n2609), .B(top_core_KE_n1929), .Y(
        top_core_KE_n2607) );
  XNOR2X1 U23863 ( .A(top_core_KE_prev_key0_reg_21_), .B(
        top_core_KE_prev_key0_reg_53_), .Y(top_core_KE_n2609) );
  XNOR2X1 U23864 ( .A(top_core_KE_n2613), .B(top_core_KE_n1931), .Y(
        top_core_KE_n2611) );
  XNOR2X1 U23865 ( .A(top_core_KE_prev_key0_reg_20_), .B(
        top_core_KE_prev_key0_reg_52_), .Y(top_core_KE_n2613) );
  XNOR2X1 U23866 ( .A(top_core_KE_n2617), .B(top_core_KE_n1933), .Y(
        top_core_KE_n2615) );
  XNOR2X1 U23867 ( .A(top_core_KE_prev_key0_reg_19_), .B(
        top_core_KE_prev_key0_reg_51_), .Y(top_core_KE_n2617) );
  XNOR2X1 U23868 ( .A(top_core_KE_n2621), .B(top_core_KE_n1935), .Y(
        top_core_KE_n2619) );
  XNOR2X1 U23869 ( .A(top_core_KE_prev_key0_reg_18_), .B(
        top_core_KE_prev_key0_reg_50_), .Y(top_core_KE_n2621) );
  XNOR2X1 U23870 ( .A(top_core_KE_n2625), .B(top_core_KE_n1937), .Y(
        top_core_KE_n2623) );
  XNOR2X1 U23871 ( .A(top_core_KE_prev_key0_reg_17_), .B(
        top_core_KE_prev_key0_reg_49_), .Y(top_core_KE_n2625) );
  XNOR2X1 U23872 ( .A(top_core_KE_n2629), .B(top_core_KE_n1939), .Y(
        top_core_KE_n2627) );
  XNOR2X1 U23873 ( .A(top_core_KE_prev_key0_reg_16_), .B(
        top_core_KE_prev_key0_reg_48_), .Y(top_core_KE_n2629) );
  XNOR2X1 U23874 ( .A(top_core_KE_n2633), .B(top_core_KE_n1941), .Y(
        top_core_KE_n2631) );
  XNOR2X1 U23875 ( .A(top_core_KE_prev_key0_reg_15_), .B(
        top_core_KE_prev_key0_reg_47_), .Y(top_core_KE_n2633) );
  XNOR2X1 U23876 ( .A(top_core_KE_n2637), .B(top_core_KE_n1943), .Y(
        top_core_KE_n2635) );
  XNOR2X1 U23877 ( .A(top_core_KE_prev_key0_reg_14_), .B(
        top_core_KE_prev_key0_reg_46_), .Y(top_core_KE_n2637) );
  XNOR2X1 U23878 ( .A(top_core_KE_n2641), .B(top_core_KE_n1945), .Y(
        top_core_KE_n2639) );
  XNOR2X1 U23879 ( .A(top_core_KE_prev_key0_reg_13_), .B(
        top_core_KE_prev_key0_reg_45_), .Y(top_core_KE_n2641) );
  XNOR2X1 U23880 ( .A(top_core_KE_n2645), .B(top_core_KE_n1947), .Y(
        top_core_KE_n2643) );
  XNOR2X1 U23881 ( .A(top_core_KE_prev_key0_reg_12_), .B(
        top_core_KE_prev_key0_reg_44_), .Y(top_core_KE_n2645) );
  XNOR2X1 U23882 ( .A(top_core_KE_n2649), .B(top_core_KE_n1949), .Y(
        top_core_KE_n2647) );
  XNOR2X1 U23883 ( .A(top_core_KE_prev_key0_reg_11_), .B(
        top_core_KE_prev_key0_reg_43_), .Y(top_core_KE_n2649) );
  XNOR2X1 U23884 ( .A(top_core_KE_n2653), .B(top_core_KE_n1951), .Y(
        top_core_KE_n2651) );
  XNOR2X1 U23885 ( .A(top_core_KE_prev_key0_reg_10_), .B(
        top_core_KE_prev_key0_reg_42_), .Y(top_core_KE_n2653) );
  XNOR2X1 U23886 ( .A(top_core_KE_n2657), .B(top_core_KE_n1953), .Y(
        top_core_KE_n2655) );
  XNOR2X1 U23887 ( .A(top_core_KE_prev_key0_reg_41_), .B(
        top_core_KE_prev_key0_reg_9_), .Y(top_core_KE_n2657) );
  XNOR2X1 U23888 ( .A(top_core_KE_n2661), .B(top_core_KE_n1955), .Y(
        top_core_KE_n2659) );
  XNOR2X1 U23889 ( .A(top_core_KE_prev_key0_reg_40_), .B(
        top_core_KE_prev_key0_reg_8_), .Y(top_core_KE_n2661) );
  XNOR2X1 U23890 ( .A(top_core_KE_n2665), .B(top_core_KE_n1957), .Y(
        top_core_KE_n2663) );
  XNOR2X1 U23891 ( .A(top_core_KE_prev_key0_reg_39_), .B(
        top_core_KE_prev_key0_reg_7_), .Y(top_core_KE_n2665) );
  XNOR2X1 U23892 ( .A(top_core_KE_n2669), .B(top_core_KE_n1959), .Y(
        top_core_KE_n2667) );
  XNOR2X1 U23893 ( .A(top_core_KE_prev_key0_reg_38_), .B(
        top_core_KE_prev_key0_reg_6_), .Y(top_core_KE_n2669) );
  XNOR2X1 U23894 ( .A(top_core_KE_n2673), .B(top_core_KE_n1961), .Y(
        top_core_KE_n2671) );
  XNOR2X1 U23895 ( .A(top_core_KE_prev_key0_reg_37_), .B(
        top_core_KE_prev_key0_reg_5_), .Y(top_core_KE_n2673) );
  XNOR2X1 U23896 ( .A(top_core_KE_n2677), .B(top_core_KE_n1963), .Y(
        top_core_KE_n2675) );
  XNOR2X1 U23897 ( .A(top_core_KE_prev_key0_reg_36_), .B(
        top_core_KE_prev_key0_reg_4_), .Y(top_core_KE_n2677) );
  XNOR2X1 U23898 ( .A(top_core_KE_n2681), .B(top_core_KE_n1965), .Y(
        top_core_KE_n2679) );
  XNOR2X1 U23899 ( .A(top_core_KE_prev_key0_reg_35_), .B(
        top_core_KE_prev_key0_reg_3_), .Y(top_core_KE_n2681) );
  XNOR2X1 U23900 ( .A(top_core_KE_n2685), .B(top_core_KE_n1967), .Y(
        top_core_KE_n2683) );
  XNOR2X1 U23901 ( .A(top_core_KE_prev_key0_reg_2_), .B(
        top_core_KE_prev_key0_reg_34_), .Y(top_core_KE_n2685) );
  XNOR2X1 U23902 ( .A(top_core_KE_n2689), .B(top_core_KE_n1969), .Y(
        top_core_KE_n2687) );
  XNOR2X1 U23903 ( .A(top_core_KE_prev_key0_reg_1_), .B(
        top_core_KE_prev_key0_reg_33_), .Y(top_core_KE_n2689) );
  XNOR2X1 U23904 ( .A(top_core_KE_n2697), .B(top_core_KE_n1971), .Y(
        top_core_KE_n2691) );
  XNOR2X1 U23905 ( .A(top_core_KE_prev_key0_reg_0_), .B(
        top_core_KE_prev_key0_reg_32_), .Y(top_core_KE_n2697) );
  XNOR2X1 U23906 ( .A(top_core_KE_n2562), .B(top_core_KE_n1909), .Y(
        top_core_KE_n2559) );
  XNOR2X1 U23907 ( .A(top_core_KE_prev_key0_reg_31_), .B(
        top_core_KE_prev_key0_reg_63_), .Y(top_core_KE_n2562) );
  XNOR2X1 U23908 ( .A(top_core_KE_n2567), .B(top_core_KE_n1911), .Y(
        top_core_KE_n2564) );
  XNOR2X1 U23909 ( .A(top_core_KE_prev_key0_reg_30_), .B(
        top_core_KE_prev_key0_reg_62_), .Y(top_core_KE_n2567) );
  XNOR2X1 U23910 ( .A(top_core_KE_n2572), .B(top_core_KE_n1913), .Y(
        top_core_KE_n2569) );
  XNOR2X1 U23911 ( .A(top_core_KE_prev_key0_reg_29_), .B(
        top_core_KE_prev_key0_reg_61_), .Y(top_core_KE_n2572) );
  XNOR2X1 U23912 ( .A(top_core_KE_n2577), .B(top_core_KE_n1915), .Y(
        top_core_KE_n2574) );
  XNOR2X1 U23913 ( .A(top_core_KE_prev_key0_reg_28_), .B(
        top_core_KE_prev_key0_reg_60_), .Y(top_core_KE_n2577) );
  XNOR2X1 U23914 ( .A(top_core_KE_n2582), .B(top_core_KE_n1917), .Y(
        top_core_KE_n2579) );
  XNOR2X1 U23915 ( .A(top_core_KE_prev_key0_reg_27_), .B(
        top_core_KE_prev_key0_reg_59_), .Y(top_core_KE_n2582) );
  XNOR2X1 U23916 ( .A(top_core_KE_n2587), .B(top_core_KE_n1919), .Y(
        top_core_KE_n2584) );
  XNOR2X1 U23917 ( .A(top_core_KE_prev_key0_reg_26_), .B(
        top_core_KE_prev_key0_reg_58_), .Y(top_core_KE_n2587) );
  XNOR2X1 U23918 ( .A(top_core_KE_n2592), .B(top_core_KE_n1921), .Y(
        top_core_KE_n2589) );
  XNOR2X1 U23919 ( .A(top_core_KE_prev_key0_reg_25_), .B(
        top_core_KE_prev_key0_reg_57_), .Y(top_core_KE_n2592) );
  XNOR2X1 U23920 ( .A(top_core_KE_n2597), .B(top_core_KE_n1923), .Y(
        top_core_KE_n2594) );
  XNOR2X1 U23921 ( .A(top_core_KE_prev_key0_reg_24_), .B(
        top_core_KE_prev_key0_reg_56_), .Y(top_core_KE_n2597) );
  OAI21XL U23922 ( .A0(n6305), .A1(top_core_EC_n25), .B0(n1), .Y(
        top_core_EC_n1026) );
  XNOR2X1 U23923 ( .A(top_core_KE_prev_key0_reg_127_), .B(top_core_KE_n2183), 
        .Y(top_core_KE_n903) );
  XNOR2XL U23924 ( .A(top_core_KE_prev_key0_reg_106_), .B(
        top_core_KE_new_sboxw_10_), .Y(top_core_KE_n1056) );
  XNOR2XL U23925 ( .A(top_core_KE_prev_key0_reg_98_), .B(
        top_core_KE_new_sboxw_2_), .Y(top_core_KE_n1112) );
  XNOR2XL U23926 ( .A(top_core_KE_prev_key0_reg_109_), .B(
        top_core_KE_new_sboxw_13_), .Y(top_core_KE_n1035) );
  XNOR2XL U23927 ( .A(top_core_KE_prev_key0_reg_101_), .B(
        top_core_KE_new_sboxw_5_), .Y(top_core_KE_n1091) );
  XNOR2XL U23928 ( .A(top_core_KE_prev_key0_reg_103_), .B(
        top_core_KE_new_sboxw_7_), .Y(top_core_KE_n1077) );
  XNOR2XL U23929 ( .A(top_core_KE_prev_key0_reg_111_), .B(
        top_core_KE_new_sboxw_15_), .Y(top_core_KE_n1021) );
  XNOR2XL U23930 ( .A(top_core_KE_prev_key0_reg_122_), .B(
        top_core_KE_new_sboxw_26_), .Y(top_core_KE_n944) );
  XNOR2XL U23931 ( .A(top_core_KE_prev_key0_reg_125_), .B(
        top_core_KE_new_sboxw_29_), .Y(top_core_KE_n923) );
  BUFX4 U23932 ( .A(top_core_KE_prev_key1_reg_28_), .Y(n1364) );
  NAND2X1 U23933 ( .A(n7017), .B(top_core_KE_key_mem_ctrl_reg_0_), .Y(
        top_core_KE_n2720) );
  BUFX4 U23934 ( .A(top_core_KE_prev_key1_reg_70_), .Y(n1342) );
  BUFX4 U23935 ( .A(top_core_KE_prev_key1_reg_78_), .Y(n1355) );
  BUFX4 U23936 ( .A(top_core_KE_prev_key1_reg_86_), .Y(n1356) );
  XNOR2X1 U23937 ( .A(top_core_KE_prev_key0_reg_104_), .B(
        top_core_KE_new_sboxw_8_), .Y(top_core_KE_n1070) );
  XNOR2X1 U23938 ( .A(top_core_KE_prev_key0_reg_96_), .B(
        top_core_KE_new_sboxw_0_), .Y(top_core_KE_n1126) );
  XNOR2X1 U23939 ( .A(top_core_KE_prev_key0_reg_110_), .B(
        top_core_KE_new_sboxw_14_), .Y(top_core_KE_n1028) );
  XNOR2X1 U23940 ( .A(top_core_KE_prev_key0_reg_102_), .B(
        top_core_KE_new_sboxw_6_), .Y(top_core_KE_n1084) );
  XNOR2X1 U23941 ( .A(top_core_KE_prev_key0_reg_120_), .B(
        top_core_KE_new_sboxw_24_), .Y(top_core_KE_n958) );
  XNOR2X1 U23942 ( .A(top_core_KE_prev_key0_reg_126_), .B(
        top_core_KE_new_sboxw_30_), .Y(top_core_KE_n913) );
  XNOR2X1 U23943 ( .A(top_core_KE_prev_key0_reg_105_), .B(
        top_core_KE_new_sboxw_9_), .Y(top_core_KE_n1063) );
  XNOR2X1 U23944 ( .A(top_core_KE_prev_key0_reg_97_), .B(
        top_core_KE_new_sboxw_1_), .Y(top_core_KE_n1119) );
  XNOR2X1 U23945 ( .A(top_core_KE_prev_key0_reg_121_), .B(
        top_core_KE_new_sboxw_25_), .Y(top_core_KE_n951) );
  XNOR2X1 U23946 ( .A(top_core_KE_prev_key0_reg_107_), .B(
        top_core_KE_new_sboxw_11_), .Y(top_core_KE_n1049) );
  XNOR2X1 U23947 ( .A(top_core_KE_prev_key0_reg_99_), .B(
        top_core_KE_new_sboxw_3_), .Y(top_core_KE_n1105) );
  XNOR2X1 U23948 ( .A(top_core_KE_prev_key0_reg_108_), .B(
        top_core_KE_new_sboxw_12_), .Y(top_core_KE_n1042) );
  XNOR2X1 U23949 ( .A(top_core_KE_prev_key0_reg_100_), .B(
        top_core_KE_new_sboxw_4_), .Y(top_core_KE_n1098) );
  XNOR2X1 U23950 ( .A(top_core_KE_prev_key0_reg_123_), .B(
        top_core_KE_new_sboxw_27_), .Y(top_core_KE_n937) );
  XNOR2X1 U23951 ( .A(top_core_KE_prev_key0_reg_124_), .B(
        top_core_KE_new_sboxw_28_), .Y(top_core_KE_n930) );
  INVX1 U23952 ( .A(top_core_KE_prev_key0_reg_127_), .Y(n6341) );
  XNOR2X1 U23953 ( .A(top_core_KE_rcon_reg_0_), .B(top_core_KE_rcon_reg_7_), 
        .Y(top_core_KE_n2711) );
  XNOR2X1 U23954 ( .A(top_core_KE_rcon_reg_3_), .B(top_core_KE_rcon_reg_7_), 
        .Y(top_core_KE_n2708) );
  INVX1 U23955 ( .A(top_core_KE_Nk0_2_), .Y(n7023) );
  XNOR2X1 U23956 ( .A(top_core_KE_prev_key0_reg_5_), .B(top_core_KE_n2060), 
        .Y(top_core_KE_n2156) );
  XNOR2X1 U23957 ( .A(top_core_KE_prev_key0_reg_7_), .B(top_core_KE_n2054), 
        .Y(top_core_KE_n2150) );
  XNOR2X1 U23958 ( .A(top_core_KE_prev_key0_reg_8_), .B(top_core_KE_n2051), 
        .Y(top_core_KE_n2147) );
  XNOR2X1 U23959 ( .A(top_core_KE_prev_key0_reg_9_), .B(top_core_KE_n2048), 
        .Y(top_core_KE_n2144) );
  XNOR2X1 U23960 ( .A(top_core_KE_prev_key0_reg_3_), .B(top_core_KE_n2066), 
        .Y(top_core_KE_n2162) );
  XNOR2X1 U23961 ( .A(top_core_KE_prev_key0_reg_4_), .B(top_core_KE_n2063), 
        .Y(top_core_KE_n2159) );
  XNOR2X1 U23962 ( .A(top_core_KE_prev_key0_reg_6_), .B(top_core_KE_n2057), 
        .Y(top_core_KE_n2153) );
  XNOR2X1 U23963 ( .A(top_core_KE_prev_key0_reg_10_), .B(top_core_KE_n2045), 
        .Y(top_core_KE_n2141) );
  XNOR2X1 U23964 ( .A(top_core_KE_prev_key0_reg_2_), .B(top_core_KE_n2069), 
        .Y(top_core_KE_n2165) );
  XNOR2X1 U23965 ( .A(top_core_KE_prev_key0_reg_13_), .B(top_core_KE_n2036), 
        .Y(top_core_KE_n2132) );
  XNOR2X1 U23966 ( .A(top_core_KE_prev_key0_reg_24_), .B(top_core_KE_n2003), 
        .Y(top_core_KE_n2099) );
  XNOR2X1 U23967 ( .A(top_core_KE_prev_key0_reg_26_), .B(top_core_KE_n1995), 
        .Y(top_core_KE_n2093) );
  XNOR2X1 U23968 ( .A(top_core_KE_prev_key0_reg_18_), .B(top_core_KE_n2021), 
        .Y(top_core_KE_n2117) );
  XNOR2X1 U23969 ( .A(top_core_KE_prev_key0_reg_27_), .B(top_core_KE_n1991), 
        .Y(top_core_KE_n2090) );
  XNOR2X1 U23970 ( .A(top_core_KE_prev_key0_reg_28_), .B(top_core_KE_n1987), 
        .Y(top_core_KE_n2087) );
  XNOR2X1 U23971 ( .A(top_core_KE_prev_key0_reg_29_), .B(top_core_KE_n1983), 
        .Y(top_core_KE_n2084) );
  XNOR2X1 U23972 ( .A(top_core_KE_prev_key0_reg_21_), .B(top_core_KE_n2012), 
        .Y(top_core_KE_n2108) );
  XNOR2X1 U23973 ( .A(top_core_KE_prev_key0_reg_30_), .B(top_core_KE_n1979), 
        .Y(top_core_KE_n2081) );
  XNOR2X1 U23974 ( .A(top_core_KE_prev_key0_reg_23_), .B(top_core_KE_n2006), 
        .Y(top_core_KE_n2102) );
  XNOR2X1 U23975 ( .A(top_core_KE_prev_key0_reg_31_), .B(top_core_KE_n1975), 
        .Y(top_core_KE_n2078) );
  XNOR2X1 U23976 ( .A(top_core_KE_prev_key0_reg_15_), .B(top_core_KE_n2030), 
        .Y(top_core_KE_n2126) );
  XNOR2X1 U23977 ( .A(top_core_KE_prev_key0_reg_25_), .B(top_core_KE_n1999), 
        .Y(top_core_KE_n2096) );
  XNOR2X1 U23978 ( .A(top_core_KE_prev_key0_reg_0_), .B(top_core_KE_n2075), 
        .Y(top_core_KE_n2171) );
  XNOR2X1 U23979 ( .A(top_core_KE_prev_key0_reg_1_), .B(top_core_KE_n2072), 
        .Y(top_core_KE_n2168) );
  XNOR2X1 U23980 ( .A(top_core_KE_prev_key0_reg_11_), .B(top_core_KE_n2042), 
        .Y(top_core_KE_n2138) );
  XNOR2X1 U23981 ( .A(top_core_KE_prev_key0_reg_12_), .B(top_core_KE_n2039), 
        .Y(top_core_KE_n2135) );
  XNOR2X1 U23982 ( .A(top_core_KE_prev_key0_reg_14_), .B(top_core_KE_n2033), 
        .Y(top_core_KE_n2129) );
  XNOR2X1 U23983 ( .A(top_core_KE_prev_key0_reg_16_), .B(top_core_KE_n2027), 
        .Y(top_core_KE_n2123) );
  XNOR2X1 U23984 ( .A(top_core_KE_prev_key0_reg_17_), .B(top_core_KE_n2024), 
        .Y(top_core_KE_n2120) );
  XNOR2X1 U23985 ( .A(top_core_KE_prev_key0_reg_19_), .B(top_core_KE_n2018), 
        .Y(top_core_KE_n2114) );
  XNOR2X1 U23986 ( .A(top_core_KE_prev_key0_reg_20_), .B(top_core_KE_n2015), 
        .Y(top_core_KE_n2111) );
  XNOR2X1 U23987 ( .A(top_core_KE_prev_key0_reg_22_), .B(top_core_KE_n2009), 
        .Y(top_core_KE_n2105) );
  INVX1 U23988 ( .A(top_core_KE_Nk0_1_), .Y(n7022) );
  BUFX4 U23989 ( .A(top_core_KE_prev_key1_reg_12_), .Y(n1350) );
  BUFX4 U23990 ( .A(top_core_KE_prev_key1_reg_4_), .Y(n1352) );
  BUFX4 U23991 ( .A(top_core_KE_prev_key1_reg_20_), .Y(n1366) );
  INVX1 U23992 ( .A(top_core_KE_prev_key1_reg_127_), .Y(n6344) );
  INVX1 U23993 ( .A(top_core_KE_prev_key1_reg_126_), .Y(n6437) );
  INVX1 U23994 ( .A(top_core_KE_prev_key1_reg_125_), .Y(n6525) );
  INVX1 U23995 ( .A(top_core_KE_prev_key1_reg_124_), .Y(n6608) );
  INVX1 U23996 ( .A(top_core_KE_prev_key1_reg_123_), .Y(n6656) );
  INVX1 U23997 ( .A(top_core_KE_prev_key1_reg_122_), .Y(n6675) );
  INVX1 U23998 ( .A(top_core_KE_prev_key1_reg_121_), .Y(n6317) );
  INVX1 U23999 ( .A(top_core_KE_prev_key1_reg_120_), .Y(n6696) );
  OAI2BB1X1 U24000 ( .A0N(n7017), .A1N(n3704), .B0(top_core_KE_n2726), .Y(
        top_core_KE_n2725) );
  AOI31X1 U24001 ( .A0(top_core_KE_n2723), .A1(top_core_KE_key_mem_ctrl_reg_1_), .A2(top_core_KE_n2724), .B0(top_core_KE_key_mem_ctrl_reg_0_), .Y(
        top_core_KE_n2726) );
  BUFX4 U24002 ( .A(top_core_KE_prev_key1_reg_94_), .Y(n1369) );
  XNOR2X1 U24003 ( .A(top_core_KE_prev_key0_reg_126_), .B(n6449), .Y(
        top_core_KE_n1370) );
  XNOR2X1 U24004 ( .A(top_core_KE_prev_key0_reg_125_), .B(n6452), .Y(
        top_core_KE_n1378) );
  XNOR2X1 U24005 ( .A(top_core_KE_prev_key0_reg_124_), .B(n6455), .Y(
        top_core_KE_n1386) );
  XNOR2X1 U24006 ( .A(top_core_KE_prev_key0_reg_123_), .B(n6458), .Y(
        top_core_KE_n1394) );
  XNOR2X1 U24007 ( .A(top_core_KE_prev_key0_reg_122_), .B(n6461), .Y(
        top_core_KE_n1402) );
  XNOR2X1 U24008 ( .A(top_core_KE_prev_key0_reg_121_), .B(n6463), .Y(
        top_core_KE_n1410) );
  XNOR2X1 U24009 ( .A(top_core_KE_prev_key0_reg_120_), .B(n6466), .Y(
        top_core_KE_n1418) );
  INVX1 U24010 ( .A(top_core_KE_prev_key0_reg_111_), .Y(n6328) );
  INVX1 U24011 ( .A(top_core_KE_prev_key0_reg_110_), .Y(n6717) );
  INVX1 U24012 ( .A(top_core_KE_prev_key0_reg_109_), .Y(n6820) );
  INVX1 U24013 ( .A(top_core_KE_prev_key0_reg_108_), .Y(n6900) );
  INVX1 U24014 ( .A(top_core_KE_prev_key0_reg_107_), .Y(n6945) );
  INVX1 U24015 ( .A(top_core_KE_prev_key0_reg_106_), .Y(n6961) );
  INVX1 U24016 ( .A(top_core_KE_prev_key0_reg_105_), .Y(n6972) );
  INVX1 U24017 ( .A(top_core_KE_prev_key0_reg_104_), .Y(n6982) );
  INVX1 U24018 ( .A(top_core_KE_prev_key0_reg_103_), .Y(n6377) );
  INVX1 U24019 ( .A(top_core_KE_prev_key0_reg_102_), .Y(n6384) );
  INVX1 U24020 ( .A(top_core_KE_prev_key0_reg_101_), .Y(n6781) );
  INVX1 U24021 ( .A(top_core_KE_prev_key0_reg_100_), .Y(n6854) );
  INVX1 U24022 ( .A(top_core_KE_prev_key0_reg_99_), .Y(n6930) );
  INVX1 U24023 ( .A(top_core_KE_prev_key0_reg_98_), .Y(n6955) );
  INVX1 U24024 ( .A(top_core_KE_prev_key0_reg_97_), .Y(n6967) );
  INVX1 U24025 ( .A(top_core_KE_prev_key0_reg_96_), .Y(n6977) );
  XNOR2X1 U24026 ( .A(top_core_KE_prev_key0_reg_127_), .B(n6448), .Y(
        top_core_KE_n1362) );
  INVX1 U24027 ( .A(top_core_KE_prev_key0_reg_63_), .Y(n6337) );
  INVX1 U24028 ( .A(top_core_KE_prev_key0_reg_121_), .Y(n6314) );
  INVX1 U24029 ( .A(top_core_KE_prev_key0_reg_120_), .Y(n6695) );
  INVX1 U24030 ( .A(top_core_KE_prev_key0_reg_122_), .Y(n6674) );
  INVX1 U24031 ( .A(top_core_KE_prev_key0_reg_123_), .Y(n6655) );
  INVX1 U24032 ( .A(top_core_KE_prev_key0_reg_124_), .Y(n6607) );
  INVX1 U24033 ( .A(top_core_KE_prev_key0_reg_125_), .Y(n6524) );
  INVX1 U24034 ( .A(top_core_KE_prev_key0_reg_126_), .Y(n6435) );
  INVX1 U24035 ( .A(top_core_KE_rcon_reg_4_), .Y(n7001) );
  INVX1 U24036 ( .A(top_core_KE_rcon_reg_5_), .Y(n7000) );
  AOI22X1 U24037 ( .A0(n1626), .A1(top_core_KE_n1044), .B0(
        top_core_KE_prev_key0_reg_108_), .B1(n2227), .Y(top_core_KE_n1043) );
  AOI22X1 U24038 ( .A0(n1626), .A1(top_core_KE_n1051), .B0(
        top_core_KE_prev_key0_reg_107_), .B1(n2227), .Y(top_core_KE_n1050) );
  AOI22X1 U24039 ( .A0(n1627), .A1(top_core_KE_n1058), .B0(
        top_core_KE_prev_key0_reg_106_), .B1(n2227), .Y(top_core_KE_n1057) );
  AOI22X1 U24040 ( .A0(n1627), .A1(top_core_KE_n1065), .B0(
        top_core_KE_prev_key0_reg_105_), .B1(n2227), .Y(top_core_KE_n1064) );
  AOI22X1 U24041 ( .A0(n1627), .A1(top_core_KE_n1072), .B0(
        top_core_KE_prev_key0_reg_104_), .B1(n2227), .Y(top_core_KE_n1071) );
  AOI22X1 U24042 ( .A0(n1627), .A1(top_core_KE_n1079), .B0(
        top_core_KE_prev_key0_reg_103_), .B1(n2227), .Y(top_core_KE_n1078) );
  AOI22X1 U24043 ( .A0(n1627), .A1(top_core_KE_n1086), .B0(
        top_core_KE_prev_key0_reg_102_), .B1(n2227), .Y(top_core_KE_n1085) );
  AOI22X1 U24044 ( .A0(n1627), .A1(top_core_KE_n1093), .B0(
        top_core_KE_prev_key0_reg_101_), .B1(n2227), .Y(top_core_KE_n1092) );
  AOI22X1 U24045 ( .A0(n1627), .A1(top_core_KE_n1100), .B0(
        top_core_KE_prev_key0_reg_100_), .B1(n2227), .Y(top_core_KE_n1099) );
  AOI22X1 U24046 ( .A0(n1627), .A1(top_core_KE_n1107), .B0(
        top_core_KE_prev_key0_reg_99_), .B1(n2227), .Y(top_core_KE_n1106) );
  AOI22X1 U24047 ( .A0(n1627), .A1(top_core_KE_n1114), .B0(
        top_core_KE_prev_key0_reg_98_), .B1(n2227), .Y(top_core_KE_n1113) );
  AOI22X1 U24048 ( .A0(n1627), .A1(top_core_KE_n1121), .B0(
        top_core_KE_prev_key0_reg_97_), .B1(n2227), .Y(top_core_KE_n1120) );
  AOI22X1 U24049 ( .A0(n1627), .A1(top_core_KE_n1128), .B0(
        top_core_KE_prev_key0_reg_96_), .B1(n2226), .Y(top_core_KE_n1127) );
  AOI22X1 U24050 ( .A0(n1627), .A1(top_core_KE_n1135), .B0(
        top_core_KE_prev_key0_reg_95_), .B1(n2226), .Y(top_core_KE_n1134) );
  AOI22X1 U24051 ( .A0(n1628), .A1(top_core_KE_n1142), .B0(
        top_core_KE_prev_key0_reg_94_), .B1(n2226), .Y(top_core_KE_n1141) );
  AOI22X1 U24052 ( .A0(n1628), .A1(top_core_KE_n1149), .B0(
        top_core_KE_prev_key0_reg_93_), .B1(n2226), .Y(top_core_KE_n1148) );
  AOI22X1 U24053 ( .A0(n1628), .A1(top_core_KE_n1156), .B0(
        top_core_KE_prev_key0_reg_92_), .B1(n2226), .Y(top_core_KE_n1155) );
  AOI22X1 U24054 ( .A0(n1628), .A1(top_core_KE_n1163), .B0(
        top_core_KE_prev_key0_reg_91_), .B1(n2226), .Y(top_core_KE_n1162) );
  AOI22X1 U24055 ( .A0(n1628), .A1(top_core_KE_n1170), .B0(
        top_core_KE_prev_key0_reg_90_), .B1(n2226), .Y(top_core_KE_n1169) );
  AOI22X1 U24056 ( .A0(n1628), .A1(top_core_KE_n1177), .B0(
        top_core_KE_prev_key0_reg_89_), .B1(n2226), .Y(top_core_KE_n1176) );
  AOI22X1 U24057 ( .A0(n1628), .A1(top_core_KE_n1184), .B0(
        top_core_KE_prev_key0_reg_88_), .B1(n2226), .Y(top_core_KE_n1183) );
  AOI22X1 U24058 ( .A0(n1628), .A1(top_core_KE_n1367), .B0(
        top_core_KE_prev_key0_reg_62_), .B1(n2226), .Y(top_core_KE_n1366) );
  AOI22X1 U24059 ( .A0(n1628), .A1(top_core_KE_n1375), .B0(
        top_core_KE_prev_key0_reg_61_), .B1(n2226), .Y(top_core_KE_n1374) );
  AOI22X1 U24060 ( .A0(n1628), .A1(top_core_KE_n1383), .B0(
        top_core_KE_prev_key0_reg_60_), .B1(n2226), .Y(top_core_KE_n1382) );
  AOI22X1 U24061 ( .A0(n1628), .A1(top_core_KE_n1391), .B0(
        top_core_KE_prev_key0_reg_59_), .B1(n2226), .Y(top_core_KE_n1390) );
  AOI22X1 U24062 ( .A0(n1628), .A1(top_core_KE_n1399), .B0(
        top_core_KE_prev_key0_reg_58_), .B1(n2226), .Y(top_core_KE_n1398) );
  AOI22X1 U24063 ( .A0(n1631), .A1(top_core_KE_n1407), .B0(
        top_core_KE_prev_key0_reg_57_), .B1(n2224), .Y(top_core_KE_n1406) );
  AOI22X1 U24064 ( .A0(n1627), .A1(top_core_KE_n1415), .B0(
        top_core_KE_prev_key0_reg_56_), .B1(n2223), .Y(top_core_KE_n1414) );
  AOI22X1 U24065 ( .A0(n1629), .A1(top_core_KE_n1423), .B0(
        top_core_KE_prev_key0_reg_55_), .B1(n2225), .Y(top_core_KE_n1422) );
  AOI22X1 U24066 ( .A0(n1630), .A1(top_core_KE_n1431), .B0(
        top_core_KE_prev_key0_reg_54_), .B1(n2222), .Y(top_core_KE_n1430) );
  AOI22X1 U24067 ( .A0(n1628), .A1(top_core_KE_n1439), .B0(
        top_core_KE_prev_key0_reg_53_), .B1(n2227), .Y(top_core_KE_n1438) );
  AOI22X1 U24068 ( .A0(n1626), .A1(top_core_KE_n1447), .B0(
        top_core_KE_prev_key0_reg_52_), .B1(n2226), .Y(top_core_KE_n1446) );
  AOI22X1 U24069 ( .A0(n1631), .A1(top_core_KE_n1455), .B0(
        top_core_KE_prev_key0_reg_51_), .B1(n2224), .Y(top_core_KE_n1454) );
  AOI22X1 U24070 ( .A0(n1627), .A1(top_core_KE_n1463), .B0(
        top_core_KE_prev_key0_reg_50_), .B1(n2223), .Y(top_core_KE_n1462) );
  AOI22X1 U24071 ( .A0(n1629), .A1(top_core_KE_n1471), .B0(
        top_core_KE_prev_key0_reg_49_), .B1(n2225), .Y(top_core_KE_n1470) );
  AOI22X1 U24072 ( .A0(n1630), .A1(top_core_KE_n1479), .B0(
        top_core_KE_prev_key0_reg_48_), .B1(n2222), .Y(top_core_KE_n1478) );
  AOI22X1 U24073 ( .A0(n1628), .A1(top_core_KE_n1487), .B0(
        top_core_KE_prev_key0_reg_47_), .B1(n2225), .Y(top_core_KE_n1486) );
  AOI22X1 U24074 ( .A0(n1629), .A1(top_core_KE_n1495), .B0(
        top_core_KE_prev_key0_reg_46_), .B1(n2225), .Y(top_core_KE_n1494) );
  AOI22X1 U24075 ( .A0(n1629), .A1(top_core_KE_n1503), .B0(
        top_core_KE_prev_key0_reg_45_), .B1(n2225), .Y(top_core_KE_n1502) );
  AOI22X1 U24076 ( .A0(n1629), .A1(top_core_KE_n1511), .B0(
        top_core_KE_prev_key0_reg_44_), .B1(n2225), .Y(top_core_KE_n1510) );
  AOI22X1 U24077 ( .A0(n1629), .A1(top_core_KE_n1519), .B0(
        top_core_KE_prev_key0_reg_43_), .B1(n2225), .Y(top_core_KE_n1518) );
  AOI22X1 U24078 ( .A0(n1629), .A1(top_core_KE_n1527), .B0(
        top_core_KE_prev_key0_reg_42_), .B1(n2225), .Y(top_core_KE_n1526) );
  AOI22X1 U24079 ( .A0(n1629), .A1(top_core_KE_n1535), .B0(
        top_core_KE_prev_key0_reg_41_), .B1(n2225), .Y(top_core_KE_n1534) );
  AOI22X1 U24080 ( .A0(n1629), .A1(top_core_KE_n1543), .B0(
        top_core_KE_prev_key0_reg_40_), .B1(n2225), .Y(top_core_KE_n1542) );
  AOI22X1 U24081 ( .A0(n1629), .A1(top_core_KE_n1551), .B0(
        top_core_KE_prev_key0_reg_39_), .B1(n2225), .Y(top_core_KE_n1550) );
  AOI22X1 U24082 ( .A0(n1629), .A1(top_core_KE_n1559), .B0(
        top_core_KE_prev_key0_reg_38_), .B1(n2225), .Y(top_core_KE_n1558) );
  AOI22X1 U24083 ( .A0(n1629), .A1(top_core_KE_n1567), .B0(
        top_core_KE_prev_key0_reg_37_), .B1(n2225), .Y(top_core_KE_n1566) );
  AOI22X1 U24084 ( .A0(n1629), .A1(top_core_KE_n1575), .B0(
        top_core_KE_prev_key0_reg_36_), .B1(n2225), .Y(top_core_KE_n1574) );
  AOI22X1 U24085 ( .A0(n1629), .A1(top_core_KE_n1583), .B0(
        top_core_KE_prev_key0_reg_35_), .B1(n2224), .Y(top_core_KE_n1582) );
  AOI22X1 U24086 ( .A0(n1630), .A1(top_core_KE_n1591), .B0(
        top_core_KE_prev_key0_reg_34_), .B1(n2224), .Y(top_core_KE_n1590) );
  AOI22X1 U24087 ( .A0(n1630), .A1(top_core_KE_n1599), .B0(
        top_core_KE_prev_key0_reg_33_), .B1(n2224), .Y(top_core_KE_n1598) );
  AOI22X1 U24088 ( .A0(n1630), .A1(top_core_KE_n1607), .B0(
        top_core_KE_prev_key0_reg_32_), .B1(n2224), .Y(top_core_KE_n1606) );
  AOI22X1 U24089 ( .A0(n1630), .A1(top_core_KE_n1615), .B0(
        top_core_KE_prev_key0_reg_31_), .B1(n2224), .Y(top_core_KE_n1614) );
  AOI22X1 U24090 ( .A0(n1631), .A1(top_core_KE_n1623), .B0(
        top_core_KE_prev_key0_reg_30_), .B1(n2224), .Y(top_core_KE_n1622) );
  AOI22X1 U24091 ( .A0(n1630), .A1(top_core_KE_n1631), .B0(
        top_core_KE_prev_key0_reg_29_), .B1(n2224), .Y(top_core_KE_n1630) );
  AOI22X1 U24092 ( .A0(n1631), .A1(top_core_KE_n1639), .B0(
        top_core_KE_prev_key0_reg_28_), .B1(n2224), .Y(top_core_KE_n1638) );
  AOI22X1 U24093 ( .A0(n1630), .A1(top_core_KE_n1647), .B0(
        top_core_KE_prev_key0_reg_27_), .B1(n2224), .Y(top_core_KE_n1646) );
  AOI22X1 U24094 ( .A0(n1631), .A1(top_core_KE_n1655), .B0(
        top_core_KE_prev_key0_reg_26_), .B1(n2224), .Y(top_core_KE_n1654) );
  AOI22X1 U24095 ( .A0(n1630), .A1(top_core_KE_n1663), .B0(
        top_core_KE_prev_key0_reg_25_), .B1(n2224), .Y(top_core_KE_n1662) );
  AOI22X1 U24096 ( .A0(n1631), .A1(top_core_KE_n1671), .B0(
        top_core_KE_prev_key0_reg_24_), .B1(n2224), .Y(top_core_KE_n1670) );
  AOI22X1 U24097 ( .A0(n1630), .A1(top_core_KE_n1679), .B0(
        top_core_KE_prev_key0_reg_23_), .B1(n2223), .Y(top_core_KE_n1678) );
  AOI22X1 U24098 ( .A0(n1631), .A1(top_core_KE_n1687), .B0(
        top_core_KE_prev_key0_reg_22_), .B1(n2223), .Y(top_core_KE_n1686) );
  AOI22X1 U24099 ( .A0(n1631), .A1(top_core_KE_n1695), .B0(
        top_core_KE_prev_key0_reg_21_), .B1(n2223), .Y(top_core_KE_n1694) );
  AOI22X1 U24100 ( .A0(n1627), .A1(top_core_KE_n1703), .B0(
        top_core_KE_prev_key0_reg_20_), .B1(n2223), .Y(top_core_KE_n1702) );
  AOI22X1 U24101 ( .A0(n1631), .A1(top_core_KE_n1711), .B0(
        top_core_KE_prev_key0_reg_19_), .B1(n2223), .Y(top_core_KE_n1710) );
  AOI22X1 U24102 ( .A0(n1629), .A1(top_core_KE_n1719), .B0(
        top_core_KE_prev_key0_reg_18_), .B1(n2223), .Y(top_core_KE_n1718) );
  AOI22X1 U24103 ( .A0(n1630), .A1(top_core_KE_n1727), .B0(
        top_core_KE_prev_key0_reg_17_), .B1(n2223), .Y(top_core_KE_n1726) );
  AOI22X1 U24104 ( .A0(n1630), .A1(top_core_KE_n1735), .B0(
        top_core_KE_prev_key0_reg_16_), .B1(n2223), .Y(top_core_KE_n1734) );
  AOI22X1 U24105 ( .A0(n1631), .A1(top_core_KE_n1743), .B0(
        top_core_KE_prev_key0_reg_15_), .B1(n2223), .Y(top_core_KE_n1742) );
  AOI22X1 U24106 ( .A0(n1628), .A1(top_core_KE_n1751), .B0(
        top_core_KE_prev_key0_reg_14_), .B1(n2223), .Y(top_core_KE_n1750) );
  AOI22X1 U24107 ( .A0(n1631), .A1(top_core_KE_n1759), .B0(
        top_core_KE_prev_key0_reg_13_), .B1(n2223), .Y(top_core_KE_n1758) );
  AOI22X1 U24108 ( .A0(n1632), .A1(top_core_KE_n1767), .B0(
        top_core_KE_prev_key0_reg_12_), .B1(n2223), .Y(top_core_KE_n1766) );
  AOI22X1 U24109 ( .A0(n1630), .A1(top_core_KE_n1775), .B0(
        top_core_KE_prev_key0_reg_11_), .B1(n2222), .Y(top_core_KE_n1774) );
  AOI22X1 U24110 ( .A0(n1633), .A1(top_core_KE_n1783), .B0(
        top_core_KE_prev_key0_reg_10_), .B1(n2222), .Y(top_core_KE_n1782) );
  AOI22X1 U24111 ( .A0(n1631), .A1(top_core_KE_n1791), .B0(
        top_core_KE_prev_key0_reg_9_), .B1(n2222), .Y(top_core_KE_n1790) );
  AOI22X1 U24112 ( .A0(n1631), .A1(top_core_KE_n1799), .B0(
        top_core_KE_prev_key0_reg_8_), .B1(n2222), .Y(top_core_KE_n1798) );
  AOI22X1 U24113 ( .A0(n1630), .A1(top_core_KE_n1807), .B0(
        top_core_KE_prev_key0_reg_7_), .B1(n2222), .Y(top_core_KE_n1806) );
  AOI22X1 U24114 ( .A0(n1626), .A1(top_core_KE_n1815), .B0(
        top_core_KE_prev_key0_reg_6_), .B1(n2222), .Y(top_core_KE_n1814) );
  AOI22X1 U24115 ( .A0(n1631), .A1(top_core_KE_n1823), .B0(
        top_core_KE_prev_key0_reg_5_), .B1(n2222), .Y(top_core_KE_n1822) );
  AOI22X1 U24116 ( .A0(n1631), .A1(top_core_KE_n1831), .B0(
        top_core_KE_prev_key0_reg_4_), .B1(n2222), .Y(top_core_KE_n1830) );
  AOI22X1 U24117 ( .A0(n1631), .A1(top_core_KE_n1839), .B0(
        top_core_KE_prev_key0_reg_3_), .B1(n2222), .Y(top_core_KE_n1838) );
  AOI22X1 U24118 ( .A0(n1627), .A1(top_core_KE_n1847), .B0(
        top_core_KE_prev_key0_reg_2_), .B1(n2222), .Y(top_core_KE_n1846) );
  AOI22X1 U24119 ( .A0(n1630), .A1(top_core_KE_n1855), .B0(
        top_core_KE_prev_key0_reg_1_), .B1(n2222), .Y(top_core_KE_n1854) );
  AOI22X1 U24120 ( .A0(n1626), .A1(top_core_KE_n1863), .B0(
        top_core_KE_prev_key0_reg_0_), .B1(n2222), .Y(top_core_KE_n1862) );
  AOI22X1 U24121 ( .A0(n1626), .A1(top_core_KE_n1023), .B0(
        top_core_KE_prev_key0_reg_111_), .B1(n2223), .Y(top_core_KE_n1022) );
  AOI22X1 U24122 ( .A0(n1626), .A1(top_core_KE_n1037), .B0(
        top_core_KE_prev_key0_reg_109_), .B1(n2224), .Y(top_core_KE_n1036) );
  AOI22X1 U24123 ( .A0(n1633), .A1(top_core_KE_n917), .B0(
        top_core_KE_prev_key0_reg_126_), .B1(top_core_KE_n918), .Y(
        top_core_KE_n916) );
  AOI22X1 U24124 ( .A0(n1626), .A1(top_core_KE_n925), .B0(
        top_core_KE_prev_key0_reg_125_), .B1(n2225), .Y(top_core_KE_n924) );
  AOI22X1 U24125 ( .A0(n1626), .A1(top_core_KE_n932), .B0(
        top_core_KE_prev_key0_reg_124_), .B1(n2227), .Y(top_core_KE_n931) );
  AOI22X1 U24126 ( .A0(n1626), .A1(top_core_KE_n939), .B0(
        top_core_KE_prev_key0_reg_123_), .B1(n2224), .Y(top_core_KE_n938) );
  AOI22X1 U24127 ( .A0(n1626), .A1(top_core_KE_n946), .B0(
        top_core_KE_prev_key0_reg_122_), .B1(n2223), .Y(top_core_KE_n945) );
  AOI22X1 U24128 ( .A0(n1626), .A1(top_core_KE_n953), .B0(
        top_core_KE_prev_key0_reg_121_), .B1(n2225), .Y(top_core_KE_n952) );
  AOI22X1 U24129 ( .A0(n1626), .A1(top_core_KE_n960), .B0(
        top_core_KE_prev_key0_reg_120_), .B1(n2222), .Y(top_core_KE_n959) );
  AOI22X1 U24130 ( .A0(n1626), .A1(top_core_KE_n1030), .B0(
        top_core_KE_prev_key0_reg_110_), .B1(n2227), .Y(top_core_KE_n1029) );
  AOI22X1 U24131 ( .A0(n2202), .A1(top_core_KE_n902), .B0(
        top_core_KE_CipherKey0_127_), .B1(n2219), .Y(top_core_KE_n901) );
  INVX1 U24132 ( .A(top_core_KE_rcon_reg_1_), .Y(n7004) );
  INVX1 U24133 ( .A(top_core_KE_rcon_reg_6_), .Y(n6999) );
  AOI221X1 U24134 ( .A0(n7022), .A1(n1332), .B0(n7023), .B1(n1333), .C0(
        top_core_KE_n2727), .Y(top_core_KE_n2724) );
  OAI221XL U24135 ( .A0(top_core_KE_n883), .A1(top_core_KE_Nk0_0_), .B0(n7019), 
        .B1(top_core_KE_n2728), .C0(top_core_KE_n728), .Y(top_core_KE_n2727)
         );
  AOI22X1 U24136 ( .A0(n1226), .A1(top_core_KE_Nk0_2_), .B0(n7014), .B1(
        top_core_KE_Nk0_1_), .Y(top_core_KE_n2728) );
  INVX1 U24137 ( .A(top_core_KE_prev_key1_reg_119_), .Y(n6395) );
  INVX1 U24138 ( .A(top_core_KE_prev_key1_reg_118_), .Y(n6403) );
  INVX1 U24139 ( .A(top_core_KE_prev_key1_reg_117_), .Y(n6481) );
  INVX1 U24140 ( .A(top_core_KE_prev_key1_reg_116_), .Y(n6561) );
  INVX1 U24141 ( .A(top_core_KE_prev_key1_reg_115_), .Y(n6640) );
  INVX1 U24142 ( .A(top_core_KE_prev_key1_reg_114_), .Y(n6668) );
  INVX1 U24143 ( .A(top_core_KE_prev_key1_reg_113_), .Y(n6683) );
  INVX1 U24144 ( .A(top_core_KE_prev_key1_reg_112_), .Y(n6690) );
  INVX1 U24145 ( .A(top_core_KE_prev_key1_reg_111_), .Y(n6330) );
  INVX1 U24146 ( .A(top_core_KE_prev_key1_reg_110_), .Y(n6719) );
  INVX1 U24147 ( .A(top_core_KE_prev_key1_reg_109_), .Y(n6821) );
  INVX1 U24148 ( .A(top_core_KE_prev_key1_reg_108_), .Y(n6901) );
  INVX1 U24149 ( .A(top_core_KE_prev_key1_reg_107_), .Y(n6946) );
  INVX1 U24150 ( .A(top_core_KE_prev_key1_reg_106_), .Y(n6962) );
  INVX1 U24151 ( .A(top_core_KE_prev_key1_reg_105_), .Y(n6973) );
  INVX1 U24152 ( .A(top_core_KE_prev_key1_reg_104_), .Y(n6983) );
  INVX1 U24153 ( .A(top_core_KE_prev_key1_reg_103_), .Y(n6379) );
  INVX1 U24154 ( .A(top_core_KE_prev_key1_reg_102_), .Y(n6386) );
  INVX1 U24155 ( .A(top_core_KE_prev_key1_reg_101_), .Y(n6783) );
  INVX1 U24156 ( .A(top_core_KE_prev_key1_reg_100_), .Y(n6855) );
  INVX1 U24157 ( .A(top_core_KE_prev_key1_reg_99_), .Y(n6931) );
  INVX1 U24158 ( .A(top_core_KE_prev_key1_reg_98_), .Y(n6956) );
  INVX1 U24159 ( .A(top_core_KE_prev_key1_reg_97_), .Y(n6968) );
  INVX1 U24160 ( .A(top_core_KE_prev_key1_reg_96_), .Y(n6978) );
  OAI2BB2X1 U24161 ( .B0(n1840), .B1(n1427), .A0N(top_core_KE_key_mem_0__72_), 
        .A1N(n1851), .Y(top_core_KE_n2786) );
  OAI2BB2X1 U24162 ( .B0(n1841), .B1(n1435), .A0N(top_core_KE_key_mem_0__64_), 
        .A1N(n1839), .Y(top_core_KE_n2794) );
  OAI2BB2X1 U24163 ( .B0(n1840), .B1(n1426), .A0N(top_core_KE_key_mem_0__73_), 
        .A1N(n1851), .Y(top_core_KE_n2785) );
  OAI2BB2X1 U24164 ( .B0(n1841), .B1(n1434), .A0N(top_core_KE_key_mem_0__65_), 
        .A1N(n1837), .Y(top_core_KE_n2793) );
  OAI2BB2X1 U24165 ( .B0(n1840), .B1(n1425), .A0N(top_core_KE_key_mem_0__74_), 
        .A1N(n1851), .Y(top_core_KE_n2784) );
  OAI2BB2X1 U24166 ( .B0(n1841), .B1(n1433), .A0N(top_core_KE_key_mem_0__66_), 
        .A1N(n1844), .Y(top_core_KE_n2792) );
  OAI2BB2X1 U24167 ( .B0(n1840), .B1(n1424), .A0N(top_core_KE_key_mem_0__75_), 
        .A1N(n1851), .Y(top_core_KE_n2783) );
  OAI2BB2X1 U24168 ( .B0(n1841), .B1(n1432), .A0N(top_core_KE_key_mem_0__67_), 
        .A1N(n1841), .Y(top_core_KE_n2791) );
  OAI2BB2X1 U24169 ( .B0(n1840), .B1(n1423), .A0N(top_core_KE_key_mem_0__76_), 
        .A1N(n1851), .Y(top_core_KE_n2782) );
  OAI2BB2X1 U24170 ( .B0(n1840), .B1(n1431), .A0N(top_core_KE_key_mem_0__68_), 
        .A1N(n1850), .Y(top_core_KE_n2790) );
  OAI2BB2X1 U24171 ( .B0(n1840), .B1(n1422), .A0N(top_core_KE_key_mem_0__77_), 
        .A1N(n1851), .Y(top_core_KE_n2781) );
  OAI2BB2X1 U24172 ( .B0(n1840), .B1(n1430), .A0N(top_core_KE_key_mem_0__69_), 
        .A1N(n1851), .Y(top_core_KE_n2789) );
  OAI2BB2X1 U24173 ( .B0(n1839), .B1(n1419), .A0N(top_core_KE_key_mem_0__80_), 
        .A1N(n1850), .Y(top_core_KE_n2778) );
  OAI2BB2X1 U24174 ( .B0(n1843), .B1(n1387), .A0N(top_core_KE_key_mem_0__112_), 
        .A1N(n1847), .Y(top_core_KE_n2746) );
  OAI2BB2X1 U24175 ( .B0(n1839), .B1(n1418), .A0N(top_core_KE_key_mem_0__81_), 
        .A1N(n1850), .Y(top_core_KE_n2777) );
  OAI2BB2X1 U24176 ( .B0(n1838), .B1(n1386), .A0N(top_core_KE_key_mem_0__113_), 
        .A1N(n1848), .Y(top_core_KE_n2745) );
  OAI2BB2X1 U24177 ( .B0(n1839), .B1(n1417), .A0N(top_core_KE_key_mem_0__82_), 
        .A1N(n1850), .Y(top_core_KE_n2776) );
  OAI2BB2X1 U24178 ( .B0(n1839), .B1(n1385), .A0N(top_core_KE_key_mem_0__114_), 
        .A1N(n1848), .Y(top_core_KE_n2744) );
  OAI2BB2X1 U24179 ( .B0(n1839), .B1(n1416), .A0N(top_core_KE_key_mem_0__83_), 
        .A1N(n1850), .Y(top_core_KE_n2775) );
  OAI2BB2X1 U24180 ( .B0(n1837), .B1(n1384), .A0N(top_core_KE_key_mem_0__115_), 
        .A1N(n1848), .Y(top_core_KE_n2743) );
  OAI2BB2X1 U24181 ( .B0(n1839), .B1(n1415), .A0N(top_core_KE_key_mem_0__84_), 
        .A1N(n1850), .Y(top_core_KE_n2774) );
  OAI2BB2X1 U24182 ( .B0(n1837), .B1(n1383), .A0N(top_core_KE_key_mem_0__116_), 
        .A1N(n1848), .Y(top_core_KE_n2742) );
  OAI2BB2X1 U24183 ( .B0(n1839), .B1(n1414), .A0N(top_core_KE_key_mem_0__85_), 
        .A1N(n1850), .Y(top_core_KE_n2773) );
  OAI2BB2X1 U24184 ( .B0(n1837), .B1(n1382), .A0N(top_core_KE_key_mem_0__117_), 
        .A1N(n1848), .Y(top_core_KE_n2741) );
  OAI2BB2X1 U24185 ( .B0(n1839), .B1(n1413), .A0N(top_core_KE_key_mem_0__86_), 
        .A1N(n1850), .Y(top_core_KE_n2772) );
  OAI2BB2X1 U24186 ( .B0(n1837), .B1(n1381), .A0N(top_core_KE_key_mem_0__118_), 
        .A1N(n1848), .Y(top_core_KE_n2740) );
  OAI2BB2X1 U24187 ( .B0(n1840), .B1(n1421), .A0N(top_core_KE_key_mem_0__78_), 
        .A1N(n1851), .Y(top_core_KE_n2780) );
  OAI2BB2X1 U24188 ( .B0(n1840), .B1(n1429), .A0N(top_core_KE_key_mem_0__70_), 
        .A1N(n1851), .Y(top_core_KE_n2788) );
  OAI2BB2X1 U24189 ( .B0(n1837), .B1(n1372), .A0N(top_core_KE_key_mem_0__127_), 
        .A1N(n1849), .Y(top_core_KE_n2731) );
  OAI2BB2X1 U24190 ( .B0(n1839), .B1(n1412), .A0N(top_core_KE_key_mem_0__87_), 
        .A1N(n1850), .Y(top_core_KE_n2771) );
  OAI2BB2X1 U24191 ( .B0(n1837), .B1(n1380), .A0N(top_core_KE_key_mem_0__119_), 
        .A1N(n1848), .Y(top_core_KE_n2739) );
  OAI2BB2X1 U24192 ( .B0(n1840), .B1(n1420), .A0N(top_core_KE_key_mem_0__79_), 
        .A1N(n1850), .Y(top_core_KE_n2779) );
  OAI2BB2X1 U24193 ( .B0(n1840), .B1(n1428), .A0N(top_core_KE_key_mem_0__71_), 
        .A1N(n1851), .Y(top_core_KE_n2787) );
  OAI2BB2X1 U24194 ( .B0(n1837), .B1(n1373), .A0N(top_core_KE_key_mem_0__126_), 
        .A1N(n1849), .Y(top_core_KE_n2732) );
  OAI2BB2X1 U24195 ( .B0(n1837), .B1(n1374), .A0N(top_core_KE_key_mem_0__125_), 
        .A1N(n1849), .Y(top_core_KE_n2733) );
  OAI2BB2X1 U24196 ( .B0(n1837), .B1(n1375), .A0N(top_core_KE_key_mem_0__124_), 
        .A1N(n1849), .Y(top_core_KE_n2734) );
  OAI2BB2X1 U24197 ( .B0(n1837), .B1(n1376), .A0N(top_core_KE_key_mem_0__123_), 
        .A1N(n1849), .Y(top_core_KE_n2735) );
  OAI2BB2X1 U24198 ( .B0(n1837), .B1(n1377), .A0N(top_core_KE_key_mem_0__122_), 
        .A1N(n1848), .Y(top_core_KE_n2736) );
  OAI2BB2X1 U24199 ( .B0(n1837), .B1(n1378), .A0N(top_core_KE_key_mem_0__121_), 
        .A1N(n1848), .Y(top_core_KE_n2737) );
  OAI2BB2X1 U24200 ( .B0(n1837), .B1(n1379), .A0N(top_core_KE_key_mem_0__120_), 
        .A1N(n1847), .Y(top_core_KE_n2738) );
  OAI2BB2X1 U24201 ( .B0(n1841), .B1(n1388), .A0N(top_core_KE_key_mem_0__111_), 
        .A1N(n1847), .Y(top_core_KE_n2747) );
  OAI2BB2X1 U24202 ( .B0(n1844), .B1(n1389), .A0N(top_core_KE_key_mem_0__110_), 
        .A1N(n1847), .Y(top_core_KE_n2748) );
  OAI2BB2X1 U24203 ( .B0(n1852), .B1(n1390), .A0N(top_core_KE_key_mem_0__109_), 
        .A1N(n1847), .Y(top_core_KE_n2749) );
  OAI2BB2X1 U24204 ( .B0(n1846), .B1(n1391), .A0N(top_core_KE_key_mem_0__108_), 
        .A1N(n1847), .Y(top_core_KE_n2750) );
  OAI2BB2X1 U24205 ( .B0(n1847), .B1(n1392), .A0N(top_core_KE_key_mem_0__107_), 
        .A1N(n1847), .Y(top_core_KE_n2751) );
  OAI2BB2X1 U24206 ( .B0(n1851), .B1(n1393), .A0N(top_core_KE_key_mem_0__106_), 
        .A1N(n1847), .Y(top_core_KE_n2752) );
  OAI2BB2X1 U24207 ( .B0(n1849), .B1(n1394), .A0N(top_core_KE_key_mem_0__105_), 
        .A1N(n1847), .Y(top_core_KE_n2753) );
  OAI2BB2X1 U24208 ( .B0(n1848), .B1(n1395), .A0N(top_core_KE_key_mem_0__104_), 
        .A1N(n1847), .Y(top_core_KE_n2754) );
  OAI2BB2X1 U24209 ( .B0(n1838), .B1(n1396), .A0N(top_core_KE_key_mem_0__103_), 
        .A1N(n1846), .Y(top_core_KE_n2755) );
  OAI2BB2X1 U24210 ( .B0(n1838), .B1(n1397), .A0N(top_core_KE_key_mem_0__102_), 
        .A1N(n1846), .Y(top_core_KE_n2756) );
  OAI2BB2X1 U24211 ( .B0(n1838), .B1(n1398), .A0N(top_core_KE_key_mem_0__101_), 
        .A1N(n1846), .Y(top_core_KE_n2757) );
  OAI2BB2X1 U24212 ( .B0(n1838), .B1(n1399), .A0N(top_core_KE_key_mem_0__100_), 
        .A1N(n1846), .Y(top_core_KE_n2758) );
  OAI2BB2X1 U24213 ( .B0(n1838), .B1(n1400), .A0N(top_core_KE_key_mem_0__99_), 
        .A1N(n1846), .Y(top_core_KE_n2759) );
  OAI2BB2X1 U24214 ( .B0(n1838), .B1(n1401), .A0N(top_core_KE_key_mem_0__98_), 
        .A1N(n1846), .Y(top_core_KE_n2760) );
  OAI2BB2X1 U24215 ( .B0(n1838), .B1(n1402), .A0N(top_core_KE_key_mem_0__97_), 
        .A1N(n1846), .Y(top_core_KE_n2761) );
  OAI2BB2X1 U24216 ( .B0(n1838), .B1(n1403), .A0N(top_core_KE_key_mem_0__96_), 
        .A1N(n1846), .Y(top_core_KE_n2762) );
  OAI2BB2X1 U24217 ( .B0(n1838), .B1(n1404), .A0N(top_core_KE_key_mem_0__95_), 
        .A1N(n1846), .Y(top_core_KE_n2763) );
  OAI2BB2X1 U24218 ( .B0(n1838), .B1(n1405), .A0N(top_core_KE_key_mem_0__94_), 
        .A1N(n1846), .Y(top_core_KE_n2764) );
  OAI2BB2X1 U24219 ( .B0(n1838), .B1(n1406), .A0N(top_core_KE_key_mem_0__93_), 
        .A1N(n1845), .Y(top_core_KE_n2765) );
  OAI2BB2X1 U24220 ( .B0(n1838), .B1(n1407), .A0N(top_core_KE_key_mem_0__92_), 
        .A1N(n1849), .Y(top_core_KE_n2766) );
  OAI2BB2X1 U24221 ( .B0(n1839), .B1(n1408), .A0N(top_core_KE_key_mem_0__91_), 
        .A1N(n1849), .Y(top_core_KE_n2767) );
  OAI2BB2X1 U24222 ( .B0(n1839), .B1(n1409), .A0N(top_core_KE_key_mem_0__90_), 
        .A1N(n1849), .Y(top_core_KE_n2768) );
  OAI2BB2X1 U24223 ( .B0(n1839), .B1(n1410), .A0N(top_core_KE_key_mem_0__89_), 
        .A1N(n1849), .Y(top_core_KE_n2769) );
  OAI2BB2X1 U24224 ( .B0(n1839), .B1(n1411), .A0N(top_core_KE_key_mem_0__88_), 
        .A1N(n1850), .Y(top_core_KE_n2770) );
  OAI2BB2X1 U24225 ( .B0(n1845), .B1(n1436), .A0N(top_core_KE_key_mem_0__63_), 
        .A1N(n1849), .Y(top_core_KE_n2795) );
  OAI2BB2X1 U24226 ( .B0(n1841), .B1(n1437), .A0N(top_core_KE_key_mem_0__62_), 
        .A1N(n1852), .Y(top_core_KE_n2796) );
  OAI2BB2X1 U24227 ( .B0(n1841), .B1(n1438), .A0N(top_core_KE_key_mem_0__61_), 
        .A1N(n1846), .Y(top_core_KE_n2797) );
  OAI2BB2X1 U24228 ( .B0(n1841), .B1(n1439), .A0N(top_core_KE_key_mem_0__60_), 
        .A1N(n1851), .Y(top_core_KE_n2798) );
  OAI2BB2X1 U24229 ( .B0(n1841), .B1(n1440), .A0N(top_core_KE_key_mem_0__59_), 
        .A1N(n1849), .Y(top_core_KE_n2799) );
  OAI2BB2X1 U24230 ( .B0(n1841), .B1(n1441), .A0N(top_core_KE_key_mem_0__58_), 
        .A1N(n1848), .Y(top_core_KE_n2800) );
  OAI2BB2X1 U24231 ( .B0(n1841), .B1(n1442), .A0N(top_core_KE_key_mem_0__57_), 
        .A1N(n1852), .Y(top_core_KE_n2801) );
  OAI2BB2X1 U24232 ( .B0(n1841), .B1(n1443), .A0N(top_core_KE_key_mem_0__56_), 
        .A1N(n1852), .Y(top_core_KE_n2802) );
  OAI2BB2X1 U24233 ( .B0(n1842), .B1(n1444), .A0N(top_core_KE_key_mem_0__55_), 
        .A1N(n1852), .Y(top_core_KE_n2803) );
  OAI2BB2X1 U24234 ( .B0(n1842), .B1(n1445), .A0N(top_core_KE_key_mem_0__54_), 
        .A1N(n1852), .Y(top_core_KE_n2804) );
  OAI2BB2X1 U24235 ( .B0(n1842), .B1(n1446), .A0N(top_core_KE_key_mem_0__53_), 
        .A1N(n1852), .Y(top_core_KE_n2805) );
  OAI2BB2X1 U24236 ( .B0(n1842), .B1(n1447), .A0N(top_core_KE_key_mem_0__52_), 
        .A1N(n1852), .Y(top_core_KE_n2806) );
  OAI2BB2X1 U24237 ( .B0(n1842), .B1(n1448), .A0N(top_core_KE_key_mem_0__51_), 
        .A1N(n1852), .Y(top_core_KE_n2807) );
  OAI2BB2X1 U24238 ( .B0(n1842), .B1(n1449), .A0N(top_core_KE_key_mem_0__50_), 
        .A1N(n1852), .Y(top_core_KE_n2808) );
  OAI2BB2X1 U24239 ( .B0(n1842), .B1(n1450), .A0N(top_core_KE_key_mem_0__49_), 
        .A1N(n1852), .Y(top_core_KE_n2809) );
  OAI2BB2X1 U24240 ( .B0(n1842), .B1(n1451), .A0N(top_core_KE_key_mem_0__48_), 
        .A1N(n1852), .Y(top_core_KE_n2810) );
  OAI2BB2X1 U24241 ( .B0(n1842), .B1(n1452), .A0N(top_core_KE_key_mem_0__47_), 
        .A1N(n1842), .Y(top_core_KE_n2811) );
  OAI2BB2X1 U24242 ( .B0(n1842), .B1(n1453), .A0N(top_core_KE_key_mem_0__46_), 
        .A1N(n1843), .Y(top_core_KE_n2812) );
  OAI2BB2X1 U24243 ( .B0(n1842), .B1(n1454), .A0N(top_core_KE_key_mem_0__45_), 
        .A1N(n1837), .Y(top_core_KE_n2813) );
  OAI2BB2X1 U24244 ( .B0(n1842), .B1(n1455), .A0N(top_core_KE_key_mem_0__44_), 
        .A1N(n1850), .Y(top_core_KE_n2814) );
  OAI2BB2X1 U24245 ( .B0(n1842), .B1(n1456), .A0N(top_core_KE_key_mem_0__43_), 
        .A1N(n1838), .Y(top_core_KE_n2815) );
  OAI2BB2X1 U24246 ( .B0(n1843), .B1(n1457), .A0N(top_core_KE_key_mem_0__42_), 
        .A1N(n1845), .Y(top_core_KE_n2816) );
  OAI2BB2X1 U24247 ( .B0(n1838), .B1(n1458), .A0N(top_core_KE_key_mem_0__41_), 
        .A1N(n1839), .Y(top_core_KE_n2817) );
  OAI2BB2X1 U24248 ( .B0(n1839), .B1(n1459), .A0N(top_core_KE_key_mem_0__40_), 
        .A1N(n1840), .Y(top_core_KE_n2818) );
  OAI2BB2X1 U24249 ( .B0(n1837), .B1(n1460), .A0N(top_core_KE_key_mem_0__39_), 
        .A1N(n1852), .Y(top_core_KE_n2819) );
  OAI2BB2X1 U24250 ( .B0(n1843), .B1(n1461), .A0N(top_core_KE_key_mem_0__38_), 
        .A1N(n1852), .Y(top_core_KE_n2820) );
  OAI2BB2X1 U24251 ( .B0(top_core_KE_n743), .B1(n1462), .A0N(
        top_core_KE_key_mem_0__37_), .A1N(n1852), .Y(top_core_KE_n2821) );
  OAI2BB2X1 U24252 ( .B0(n1843), .B1(n1463), .A0N(top_core_KE_key_mem_0__36_), 
        .A1N(n1852), .Y(top_core_KE_n2822) );
  OAI2BB2X1 U24253 ( .B0(n1844), .B1(n1464), .A0N(top_core_KE_key_mem_0__35_), 
        .A1N(n1852), .Y(top_core_KE_n2823) );
  OAI2BB2X1 U24254 ( .B0(n1844), .B1(n1465), .A0N(top_core_KE_key_mem_0__34_), 
        .A1N(n1842), .Y(top_core_KE_n2824) );
  OAI2BB2X1 U24255 ( .B0(n1844), .B1(n1466), .A0N(top_core_KE_key_mem_0__33_), 
        .A1N(n1843), .Y(top_core_KE_n2825) );
  OAI2BB2X1 U24256 ( .B0(n1843), .B1(n1467), .A0N(top_core_KE_key_mem_0__32_), 
        .A1N(n1838), .Y(top_core_KE_n2826) );
  OAI2BB2X1 U24257 ( .B0(n1845), .B1(n1468), .A0N(top_core_KE_key_mem_0__31_), 
        .A1N(n1845), .Y(top_core_KE_n2827) );
  OAI2BB2X1 U24258 ( .B0(n1845), .B1(n1469), .A0N(top_core_KE_key_mem_0__30_), 
        .A1N(n1840), .Y(top_core_KE_n2828) );
  OAI2BB2X1 U24259 ( .B0(n1844), .B1(n1470), .A0N(top_core_KE_key_mem_0__29_), 
        .A1N(n1851), .Y(top_core_KE_n2829) );
  OAI2BB2X1 U24260 ( .B0(n1845), .B1(n1471), .A0N(top_core_KE_key_mem_0__28_), 
        .A1N(n1851), .Y(top_core_KE_n2830) );
  OAI2BB2X1 U24261 ( .B0(n1844), .B1(n1472), .A0N(top_core_KE_key_mem_0__27_), 
        .A1N(n1851), .Y(top_core_KE_n2831) );
  OAI2BB2X1 U24262 ( .B0(n1845), .B1(n1473), .A0N(top_core_KE_key_mem_0__26_), 
        .A1N(n1851), .Y(top_core_KE_n2832) );
  OAI2BB2X1 U24263 ( .B0(n1845), .B1(n1474), .A0N(top_core_KE_key_mem_0__25_), 
        .A1N(n1851), .Y(top_core_KE_n2833) );
  OAI2BB2X1 U24264 ( .B0(n1844), .B1(n1475), .A0N(top_core_KE_key_mem_0__24_), 
        .A1N(n1850), .Y(top_core_KE_n2834) );
  OAI2BB2X1 U24265 ( .B0(n1844), .B1(n1476), .A0N(top_core_KE_key_mem_0__23_), 
        .A1N(n1850), .Y(top_core_KE_n2835) );
  OAI2BB2X1 U24266 ( .B0(n1843), .B1(n1477), .A0N(top_core_KE_key_mem_0__22_), 
        .A1N(n1850), .Y(top_core_KE_n2836) );
  OAI2BB2X1 U24267 ( .B0(n1843), .B1(n1478), .A0N(top_core_KE_key_mem_0__21_), 
        .A1N(n1850), .Y(top_core_KE_n2837) );
  OAI2BB2X1 U24268 ( .B0(n1843), .B1(n1479), .A0N(top_core_KE_key_mem_0__20_), 
        .A1N(n1850), .Y(top_core_KE_n2838) );
  OAI2BB2X1 U24269 ( .B0(n1843), .B1(n1480), .A0N(top_core_KE_key_mem_0__19_), 
        .A1N(n1849), .Y(top_core_KE_n2839) );
  OAI2BB2X1 U24270 ( .B0(n1844), .B1(n1481), .A0N(top_core_KE_key_mem_0__18_), 
        .A1N(n1849), .Y(top_core_KE_n2840) );
  OAI2BB2X1 U24271 ( .B0(n1843), .B1(n1482), .A0N(top_core_KE_key_mem_0__17_), 
        .A1N(n1846), .Y(top_core_KE_n2841) );
  OAI2BB2X1 U24272 ( .B0(n1841), .B1(n1483), .A0N(top_core_KE_key_mem_0__16_), 
        .A1N(n1847), .Y(top_core_KE_n2842) );
  OAI2BB2X1 U24273 ( .B0(n1843), .B1(n1484), .A0N(top_core_KE_key_mem_0__15_), 
        .A1N(n1846), .Y(top_core_KE_n2843) );
  OAI2BB2X1 U24274 ( .B0(n1843), .B1(n1485), .A0N(top_core_KE_key_mem_0__14_), 
        .A1N(n1846), .Y(top_core_KE_n2844) );
  OAI2BB2X1 U24275 ( .B0(n1844), .B1(n1486), .A0N(top_core_KE_key_mem_0__13_), 
        .A1N(n1846), .Y(top_core_KE_n2845) );
  OAI2BB2X1 U24276 ( .B0(n1844), .B1(n1487), .A0N(top_core_KE_key_mem_0__12_), 
        .A1N(n1846), .Y(top_core_KE_n2846) );
  OAI2BB2X1 U24277 ( .B0(n1845), .B1(n1488), .A0N(top_core_KE_key_mem_0__11_), 
        .A1N(n1847), .Y(top_core_KE_n2847) );
  OAI2BB2X1 U24278 ( .B0(n1845), .B1(n1489), .A0N(top_core_KE_key_mem_0__10_), 
        .A1N(n1847), .Y(top_core_KE_n2848) );
  OAI2BB2X1 U24279 ( .B0(n1844), .B1(n1490), .A0N(top_core_KE_key_mem_0__9_), 
        .A1N(n1847), .Y(top_core_KE_n2849) );
  OAI2BB2X1 U24280 ( .B0(n1845), .B1(n1491), .A0N(top_core_KE_key_mem_0__8_), 
        .A1N(n1847), .Y(top_core_KE_n2850) );
  OAI2BB2X1 U24281 ( .B0(n1844), .B1(n1492), .A0N(top_core_KE_key_mem_0__7_), 
        .A1N(n1848), .Y(top_core_KE_n2851) );
  OAI2BB2X1 U24282 ( .B0(n1845), .B1(n1493), .A0N(top_core_KE_key_mem_0__6_), 
        .A1N(n1848), .Y(top_core_KE_n2852) );
  OAI2BB2X1 U24283 ( .B0(n1844), .B1(n1494), .A0N(top_core_KE_key_mem_0__5_), 
        .A1N(n1848), .Y(top_core_KE_n2853) );
  OAI2BB2X1 U24284 ( .B0(n1843), .B1(n1495), .A0N(top_core_KE_key_mem_0__4_), 
        .A1N(n1848), .Y(top_core_KE_n2854) );
  OAI2BB2X1 U24285 ( .B0(n1845), .B1(n1496), .A0N(top_core_KE_key_mem_0__3_), 
        .A1N(n1848), .Y(top_core_KE_n2855) );
  OAI2BB2X1 U24286 ( .B0(n1843), .B1(n1497), .A0N(top_core_KE_key_mem_0__2_), 
        .A1N(n1848), .Y(top_core_KE_n2856) );
  OAI2BB2X1 U24287 ( .B0(n1840), .B1(n1498), .A0N(top_core_KE_key_mem_0__1_), 
        .A1N(n1849), .Y(top_core_KE_n2857) );
  OAI2BB2X1 U24288 ( .B0(n1842), .B1(n1499), .A0N(top_core_KE_key_mem_0__0_), 
        .A1N(n1849), .Y(top_core_KE_n2858) );
  OAI2BB2X1 U24289 ( .B0(n1841), .B1(n1371), .A0N(top_core_KE_key_mem_0__128_), 
        .A1N(n1849), .Y(top_core_KE_n2730) );
  OAI2BB2X1 U24290 ( .B0(n1427), .B1(n1860), .A0N(top_core_KE_key_mem_1__72_), 
        .A1N(n1871), .Y(top_core_KE_n2915) );
  OAI2BB2X1 U24291 ( .B0(n1427), .B1(n1878), .A0N(top_core_KE_key_mem_2__72_), 
        .A1N(n1889), .Y(top_core_KE_n3044) );
  OAI2BB2X1 U24292 ( .B0(n1427), .B1(n1898), .A0N(top_core_KE_key_mem_3__72_), 
        .A1N(n1908), .Y(top_core_KE_n3173) );
  OAI2BB2X1 U24293 ( .B0(n1427), .B1(n1918), .A0N(top_core_KE_key_mem_4__72_), 
        .A1N(n1929), .Y(top_core_KE_n3302) );
  OAI2BB2X1 U24294 ( .B0(n1427), .B1(n1952), .A0N(top_core_KE_key_mem_5__72_), 
        .A1N(n1948), .Y(top_core_KE_n3431) );
  OAI2BB2X1 U24295 ( .B0(n1427), .B1(n1958), .A0N(top_core_KE_key_mem_6__72_), 
        .A1N(n1968), .Y(top_core_KE_n3560) );
  OAI2BB2X1 U24296 ( .B0(n1427), .B1(n1977), .A0N(top_core_KE_key_mem_7__72_), 
        .A1N(n1988), .Y(top_core_KE_n3689) );
  OAI2BB2X1 U24297 ( .B0(n1427), .B1(n2038), .A0N(top_core_KE_key_mem_10__72_), 
        .A1N(n2047), .Y(top_core_KE_n4076) );
  OAI2BB2X1 U24298 ( .B0(n1427), .B1(n2057), .A0N(top_core_KE_key_mem_11__72_), 
        .A1N(n2068), .Y(top_core_KE_n4205) );
  OAI2BB2X1 U24299 ( .B0(n1427), .B1(n2092), .A0N(top_core_KE_key_mem_12__72_), 
        .A1N(n2088), .Y(top_core_KE_n4334) );
  OAI2BB2X1 U24300 ( .B0(n1427), .B1(n2097), .A0N(top_core_KE_key_mem_13__72_), 
        .A1N(n2108), .Y(top_core_KE_n4463) );
  OAI2BB2X1 U24301 ( .B0(n1427), .B1(n2117), .A0N(top_core_KE_key_mem_14__72_), 
        .A1N(n2128), .Y(top_core_KE_n4592) );
  OAI2BB2X1 U24302 ( .B0(n1435), .B1(n1860), .A0N(top_core_KE_key_mem_1__64_), 
        .A1N(n1872), .Y(top_core_KE_n2923) );
  OAI2BB2X1 U24303 ( .B0(n1435), .B1(n1879), .A0N(top_core_KE_key_mem_2__64_), 
        .A1N(n1890), .Y(top_core_KE_n3052) );
  OAI2BB2X1 U24304 ( .B0(n1435), .B1(n1905), .A0N(top_core_KE_key_mem_3__64_), 
        .A1N(n1909), .Y(top_core_KE_n3181) );
  OAI2BB2X1 U24305 ( .B0(n1435), .B1(n1919), .A0N(top_core_KE_key_mem_4__64_), 
        .A1N(n1927), .Y(top_core_KE_n3310) );
  OAI2BB2X1 U24306 ( .B0(n1435), .B1(n1938), .A0N(top_core_KE_key_mem_5__64_), 
        .A1N(n1949), .Y(top_core_KE_n3439) );
  OAI2BB2X1 U24307 ( .B0(n1435), .B1(n1959), .A0N(top_core_KE_key_mem_6__64_), 
        .A1N(n1969), .Y(top_core_KE_n3568) );
  OAI2BB2X1 U24308 ( .B0(n1435), .B1(n1978), .A0N(top_core_KE_key_mem_7__64_), 
        .A1N(n1989), .Y(top_core_KE_n3697) );
  OAI2BB2X1 U24309 ( .B0(n1435), .B1(n2039), .A0N(top_core_KE_key_mem_10__64_), 
        .A1N(n2049), .Y(top_core_KE_n4084) );
  OAI2BB2X1 U24310 ( .B0(n1435), .B1(n2058), .A0N(top_core_KE_key_mem_11__64_), 
        .A1N(n2069), .Y(top_core_KE_n4213) );
  OAI2BB2X1 U24311 ( .B0(n1435), .B1(n2078), .A0N(top_core_KE_key_mem_12__64_), 
        .A1N(n2089), .Y(top_core_KE_n4342) );
  OAI2BB2X1 U24312 ( .B0(n1435), .B1(n2098), .A0N(top_core_KE_key_mem_13__64_), 
        .A1N(n2109), .Y(top_core_KE_n4471) );
  OAI2BB2X1 U24313 ( .B0(n1435), .B1(n2118), .A0N(top_core_KE_key_mem_14__64_), 
        .A1N(n2129), .Y(top_core_KE_n4600) );
  OAI2BB2X1 U24314 ( .B0(n1426), .B1(n1860), .A0N(top_core_KE_key_mem_1__73_), 
        .A1N(n1871), .Y(top_core_KE_n2914) );
  OAI2BB2X1 U24315 ( .B0(n1426), .B1(n1878), .A0N(top_core_KE_key_mem_2__73_), 
        .A1N(n1889), .Y(top_core_KE_n3043) );
  OAI2BB2X1 U24316 ( .B0(n1426), .B1(n1898), .A0N(top_core_KE_key_mem_3__73_), 
        .A1N(n1908), .Y(top_core_KE_n3172) );
  OAI2BB2X1 U24317 ( .B0(n1426), .B1(n1918), .A0N(top_core_KE_key_mem_4__73_), 
        .A1N(n1929), .Y(top_core_KE_n3301) );
  OAI2BB2X1 U24318 ( .B0(n1426), .B1(n1946), .A0N(top_core_KE_key_mem_5__73_), 
        .A1N(n1948), .Y(top_core_KE_n3430) );
  OAI2BB2X1 U24319 ( .B0(n1426), .B1(n1958), .A0N(top_core_KE_key_mem_6__73_), 
        .A1N(n1968), .Y(top_core_KE_n3559) );
  OAI2BB2X1 U24320 ( .B0(n1426), .B1(n1977), .A0N(top_core_KE_key_mem_7__73_), 
        .A1N(n1988), .Y(top_core_KE_n3688) );
  OAI2BB2X1 U24321 ( .B0(n1426), .B1(n2038), .A0N(top_core_KE_key_mem_10__73_), 
        .A1N(n2048), .Y(top_core_KE_n4075) );
  OAI2BB2X1 U24322 ( .B0(n1426), .B1(n2057), .A0N(top_core_KE_key_mem_11__73_), 
        .A1N(n2068), .Y(top_core_KE_n4204) );
  OAI2BB2X1 U24323 ( .B0(n1426), .B1(n2086), .A0N(top_core_KE_key_mem_12__73_), 
        .A1N(n2088), .Y(top_core_KE_n4333) );
  OAI2BB2X1 U24324 ( .B0(n1426), .B1(n2097), .A0N(top_core_KE_key_mem_13__73_), 
        .A1N(n2108), .Y(top_core_KE_n4462) );
  OAI2BB2X1 U24325 ( .B0(n1426), .B1(n2117), .A0N(top_core_KE_key_mem_14__73_), 
        .A1N(n2128), .Y(top_core_KE_n4591) );
  OAI2BB2X1 U24326 ( .B0(n1434), .B1(n1860), .A0N(top_core_KE_key_mem_1__65_), 
        .A1N(n1872), .Y(top_core_KE_n2922) );
  OAI2BB2X1 U24327 ( .B0(n1434), .B1(n1879), .A0N(top_core_KE_key_mem_2__65_), 
        .A1N(n1890), .Y(top_core_KE_n3051) );
  OAI2BB2X1 U24328 ( .B0(n1434), .B1(n1910), .A0N(top_core_KE_key_mem_3__65_), 
        .A1N(n1909), .Y(top_core_KE_n3180) );
  OAI2BB2X1 U24329 ( .B0(n1434), .B1(n1919), .A0N(top_core_KE_key_mem_4__65_), 
        .A1N(n1928), .Y(top_core_KE_n3309) );
  OAI2BB2X1 U24330 ( .B0(n1434), .B1(n1938), .A0N(top_core_KE_key_mem_5__65_), 
        .A1N(n1949), .Y(top_core_KE_n3438) );
  OAI2BB2X1 U24331 ( .B0(n1434), .B1(n1959), .A0N(top_core_KE_key_mem_6__65_), 
        .A1N(n1969), .Y(top_core_KE_n3567) );
  OAI2BB2X1 U24332 ( .B0(n1434), .B1(n1978), .A0N(top_core_KE_key_mem_7__65_), 
        .A1N(n1989), .Y(top_core_KE_n3696) );
  OAI2BB2X1 U24333 ( .B0(n1434), .B1(n2039), .A0N(top_core_KE_key_mem_10__65_), 
        .A1N(n2049), .Y(top_core_KE_n4083) );
  OAI2BB2X1 U24334 ( .B0(n1434), .B1(n2058), .A0N(top_core_KE_key_mem_11__65_), 
        .A1N(n2069), .Y(top_core_KE_n4212) );
  OAI2BB2X1 U24335 ( .B0(n1434), .B1(n2078), .A0N(top_core_KE_key_mem_12__65_), 
        .A1N(n2089), .Y(top_core_KE_n4341) );
  OAI2BB2X1 U24336 ( .B0(n1434), .B1(n2098), .A0N(top_core_KE_key_mem_13__65_), 
        .A1N(n2109), .Y(top_core_KE_n4470) );
  OAI2BB2X1 U24337 ( .B0(n1434), .B1(n2118), .A0N(top_core_KE_key_mem_14__65_), 
        .A1N(n2129), .Y(top_core_KE_n4599) );
  OAI2BB2X1 U24338 ( .B0(n1425), .B1(n1860), .A0N(top_core_KE_key_mem_1__74_), 
        .A1N(n1871), .Y(top_core_KE_n2913) );
  OAI2BB2X1 U24339 ( .B0(n1425), .B1(n1878), .A0N(top_core_KE_key_mem_2__74_), 
        .A1N(n1889), .Y(top_core_KE_n3042) );
  OAI2BB2X1 U24340 ( .B0(n1425), .B1(n1898), .A0N(top_core_KE_key_mem_3__74_), 
        .A1N(n1908), .Y(top_core_KE_n3171) );
  OAI2BB2X1 U24341 ( .B0(n1425), .B1(n1918), .A0N(top_core_KE_key_mem_4__74_), 
        .A1N(n1929), .Y(top_core_KE_n3300) );
  OAI2BB2X1 U24342 ( .B0(n1425), .B1(n1947), .A0N(top_core_KE_key_mem_5__74_), 
        .A1N(n1948), .Y(top_core_KE_n3429) );
  OAI2BB2X1 U24343 ( .B0(n1425), .B1(n1958), .A0N(top_core_KE_key_mem_6__74_), 
        .A1N(n1968), .Y(top_core_KE_n3558) );
  OAI2BB2X1 U24344 ( .B0(n1425), .B1(n1977), .A0N(top_core_KE_key_mem_7__74_), 
        .A1N(n1988), .Y(top_core_KE_n3687) );
  OAI2BB2X1 U24345 ( .B0(n1425), .B1(n2038), .A0N(top_core_KE_key_mem_10__74_), 
        .A1N(n2046), .Y(top_core_KE_n4074) );
  OAI2BB2X1 U24346 ( .B0(n1425), .B1(n2057), .A0N(top_core_KE_key_mem_11__74_), 
        .A1N(n2068), .Y(top_core_KE_n4203) );
  OAI2BB2X1 U24347 ( .B0(n1425), .B1(n2087), .A0N(top_core_KE_key_mem_12__74_), 
        .A1N(n2088), .Y(top_core_KE_n4332) );
  OAI2BB2X1 U24348 ( .B0(n1425), .B1(n2097), .A0N(top_core_KE_key_mem_13__74_), 
        .A1N(n2108), .Y(top_core_KE_n4461) );
  OAI2BB2X1 U24349 ( .B0(n1425), .B1(n2117), .A0N(top_core_KE_key_mem_14__74_), 
        .A1N(n2128), .Y(top_core_KE_n4590) );
  OAI2BB2X1 U24350 ( .B0(n1433), .B1(n1860), .A0N(top_core_KE_key_mem_1__66_), 
        .A1N(n1872), .Y(top_core_KE_n2921) );
  OAI2BB2X1 U24351 ( .B0(n1433), .B1(n1879), .A0N(top_core_KE_key_mem_2__66_), 
        .A1N(n1890), .Y(top_core_KE_n3050) );
  OAI2BB2X1 U24352 ( .B0(n1433), .B1(n1911), .A0N(top_core_KE_key_mem_3__66_), 
        .A1N(n1909), .Y(top_core_KE_n3179) );
  OAI2BB2X1 U24353 ( .B0(n1433), .B1(n1919), .A0N(top_core_KE_key_mem_4__66_), 
        .A1N(n1926), .Y(top_core_KE_n3308) );
  OAI2BB2X1 U24354 ( .B0(n1433), .B1(n1938), .A0N(top_core_KE_key_mem_5__66_), 
        .A1N(n1949), .Y(top_core_KE_n3437) );
  OAI2BB2X1 U24355 ( .B0(n1433), .B1(n1959), .A0N(top_core_KE_key_mem_6__66_), 
        .A1N(n1969), .Y(top_core_KE_n3566) );
  OAI2BB2X1 U24356 ( .B0(n1433), .B1(n1978), .A0N(top_core_KE_key_mem_7__66_), 
        .A1N(n1989), .Y(top_core_KE_n3695) );
  OAI2BB2X1 U24357 ( .B0(n1433), .B1(n2039), .A0N(top_core_KE_key_mem_10__66_), 
        .A1N(n2049), .Y(top_core_KE_n4082) );
  OAI2BB2X1 U24358 ( .B0(n1433), .B1(n2058), .A0N(top_core_KE_key_mem_11__66_), 
        .A1N(n2069), .Y(top_core_KE_n4211) );
  OAI2BB2X1 U24359 ( .B0(n1433), .B1(n2078), .A0N(top_core_KE_key_mem_12__66_), 
        .A1N(n2089), .Y(top_core_KE_n4340) );
  OAI2BB2X1 U24360 ( .B0(n1433), .B1(n2098), .A0N(top_core_KE_key_mem_13__66_), 
        .A1N(n2109), .Y(top_core_KE_n4469) );
  OAI2BB2X1 U24361 ( .B0(n1433), .B1(n2118), .A0N(top_core_KE_key_mem_14__66_), 
        .A1N(n2129), .Y(top_core_KE_n4598) );
  OAI2BB2X1 U24362 ( .B0(n1424), .B1(n1860), .A0N(top_core_KE_key_mem_1__75_), 
        .A1N(n1871), .Y(top_core_KE_n2912) );
  OAI2BB2X1 U24363 ( .B0(n1424), .B1(n1878), .A0N(top_core_KE_key_mem_2__75_), 
        .A1N(n1889), .Y(top_core_KE_n3041) );
  OAI2BB2X1 U24364 ( .B0(n1424), .B1(n1898), .A0N(top_core_KE_key_mem_3__75_), 
        .A1N(n1908), .Y(top_core_KE_n3170) );
  OAI2BB2X1 U24365 ( .B0(n1424), .B1(n1918), .A0N(top_core_KE_key_mem_4__75_), 
        .A1N(n1929), .Y(top_core_KE_n3299) );
  OAI2BB2X1 U24366 ( .B0(n1424), .B1(n1950), .A0N(top_core_KE_key_mem_5__75_), 
        .A1N(n1948), .Y(top_core_KE_n3428) );
  OAI2BB2X1 U24367 ( .B0(n1424), .B1(n1958), .A0N(top_core_KE_key_mem_6__75_), 
        .A1N(n1968), .Y(top_core_KE_n3557) );
  OAI2BB2X1 U24368 ( .B0(n1424), .B1(n1977), .A0N(top_core_KE_key_mem_7__75_), 
        .A1N(n1988), .Y(top_core_KE_n3686) );
  OAI2BB2X1 U24369 ( .B0(n1424), .B1(n2038), .A0N(top_core_KE_key_mem_10__75_), 
        .A1N(n2050), .Y(top_core_KE_n4073) );
  OAI2BB2X1 U24370 ( .B0(n1424), .B1(n2057), .A0N(top_core_KE_key_mem_11__75_), 
        .A1N(n2068), .Y(top_core_KE_n4202) );
  OAI2BB2X1 U24371 ( .B0(n1424), .B1(n2090), .A0N(top_core_KE_key_mem_12__75_), 
        .A1N(n2088), .Y(top_core_KE_n4331) );
  OAI2BB2X1 U24372 ( .B0(n1424), .B1(n2097), .A0N(top_core_KE_key_mem_13__75_), 
        .A1N(n2108), .Y(top_core_KE_n4460) );
  OAI2BB2X1 U24373 ( .B0(n1424), .B1(n2117), .A0N(top_core_KE_key_mem_14__75_), 
        .A1N(n2128), .Y(top_core_KE_n4589) );
  OAI2BB2X1 U24374 ( .B0(n1432), .B1(n1860), .A0N(top_core_KE_key_mem_1__67_), 
        .A1N(n1872), .Y(top_core_KE_n2920) );
  OAI2BB2X1 U24375 ( .B0(n1432), .B1(n1879), .A0N(top_core_KE_key_mem_2__67_), 
        .A1N(n1889), .Y(top_core_KE_n3049) );
  OAI2BB2X1 U24376 ( .B0(n1432), .B1(n1912), .A0N(top_core_KE_key_mem_3__67_), 
        .A1N(n1908), .Y(top_core_KE_n3178) );
  OAI2BB2X1 U24377 ( .B0(n1432), .B1(n1919), .A0N(top_core_KE_key_mem_4__67_), 
        .A1N(n1929), .Y(top_core_KE_n3307) );
  OAI2BB2X1 U24378 ( .B0(n1432), .B1(n1938), .A0N(top_core_KE_key_mem_5__67_), 
        .A1N(n1948), .Y(top_core_KE_n3436) );
  OAI2BB2X1 U24379 ( .B0(n1432), .B1(n1959), .A0N(top_core_KE_key_mem_6__67_), 
        .A1N(n1968), .Y(top_core_KE_n3565) );
  OAI2BB2X1 U24380 ( .B0(n1432), .B1(n1978), .A0N(top_core_KE_key_mem_7__67_), 
        .A1N(n1988), .Y(top_core_KE_n3694) );
  OAI2BB2X1 U24381 ( .B0(n1432), .B1(n2039), .A0N(top_core_KE_key_mem_10__67_), 
        .A1N(n2051), .Y(top_core_KE_n4081) );
  OAI2BB2X1 U24382 ( .B0(n1432), .B1(n2058), .A0N(top_core_KE_key_mem_11__67_), 
        .A1N(n2068), .Y(top_core_KE_n4210) );
  OAI2BB2X1 U24383 ( .B0(n1432), .B1(n2078), .A0N(top_core_KE_key_mem_12__67_), 
        .A1N(n2088), .Y(top_core_KE_n4339) );
  OAI2BB2X1 U24384 ( .B0(n1432), .B1(n2098), .A0N(top_core_KE_key_mem_13__67_), 
        .A1N(n2108), .Y(top_core_KE_n4468) );
  OAI2BB2X1 U24385 ( .B0(n1432), .B1(n2118), .A0N(top_core_KE_key_mem_14__67_), 
        .A1N(n2128), .Y(top_core_KE_n4597) );
  OAI2BB2X1 U24386 ( .B0(n1423), .B1(n1860), .A0N(top_core_KE_key_mem_1__76_), 
        .A1N(n1871), .Y(top_core_KE_n2911) );
  OAI2BB2X1 U24387 ( .B0(n1423), .B1(n1878), .A0N(top_core_KE_key_mem_2__76_), 
        .A1N(n1889), .Y(top_core_KE_n3040) );
  OAI2BB2X1 U24388 ( .B0(n1423), .B1(n1898), .A0N(top_core_KE_key_mem_3__76_), 
        .A1N(n1908), .Y(top_core_KE_n3169) );
  OAI2BB2X1 U24389 ( .B0(n1423), .B1(n1918), .A0N(top_core_KE_key_mem_4__76_), 
        .A1N(n1929), .Y(top_core_KE_n3298) );
  OAI2BB2X1 U24390 ( .B0(n1423), .B1(n1951), .A0N(top_core_KE_key_mem_5__76_), 
        .A1N(n1948), .Y(top_core_KE_n3427) );
  OAI2BB2X1 U24391 ( .B0(n1423), .B1(n1958), .A0N(top_core_KE_key_mem_6__76_), 
        .A1N(n1968), .Y(top_core_KE_n3556) );
  OAI2BB2X1 U24392 ( .B0(n1423), .B1(n1977), .A0N(top_core_KE_key_mem_7__76_), 
        .A1N(n1988), .Y(top_core_KE_n3685) );
  OAI2BB2X1 U24393 ( .B0(n1423), .B1(n2038), .A0N(top_core_KE_key_mem_10__76_), 
        .A1N(n2045), .Y(top_core_KE_n4072) );
  OAI2BB2X1 U24394 ( .B0(n1423), .B1(n2057), .A0N(top_core_KE_key_mem_11__76_), 
        .A1N(n2068), .Y(top_core_KE_n4201) );
  OAI2BB2X1 U24395 ( .B0(n1423), .B1(n2091), .A0N(top_core_KE_key_mem_12__76_), 
        .A1N(n2088), .Y(top_core_KE_n4330) );
  OAI2BB2X1 U24396 ( .B0(n1423), .B1(n2097), .A0N(top_core_KE_key_mem_13__76_), 
        .A1N(n2108), .Y(top_core_KE_n4459) );
  OAI2BB2X1 U24397 ( .B0(n1423), .B1(n2117), .A0N(top_core_KE_key_mem_14__76_), 
        .A1N(n2128), .Y(top_core_KE_n4588) );
  OAI2BB2X1 U24398 ( .B0(n1431), .B1(n1860), .A0N(top_core_KE_key_mem_1__68_), 
        .A1N(n1872), .Y(top_core_KE_n2919) );
  OAI2BB2X1 U24399 ( .B0(n1431), .B1(n1879), .A0N(top_core_KE_key_mem_2__68_), 
        .A1N(n1889), .Y(top_core_KE_n3048) );
  OAI2BB2X1 U24400 ( .B0(n1431), .B1(n1906), .A0N(top_core_KE_key_mem_3__68_), 
        .A1N(n1908), .Y(top_core_KE_n3177) );
  OAI2BB2X1 U24401 ( .B0(n1431), .B1(n1919), .A0N(top_core_KE_key_mem_4__68_), 
        .A1N(n1929), .Y(top_core_KE_n3306) );
  OAI2BB2X1 U24402 ( .B0(n1431), .B1(n1938), .A0N(top_core_KE_key_mem_5__68_), 
        .A1N(n1948), .Y(top_core_KE_n3435) );
  OAI2BB2X1 U24403 ( .B0(n1431), .B1(n1959), .A0N(top_core_KE_key_mem_6__68_), 
        .A1N(n1968), .Y(top_core_KE_n3564) );
  OAI2BB2X1 U24404 ( .B0(n1431), .B1(n1978), .A0N(top_core_KE_key_mem_7__68_), 
        .A1N(n1988), .Y(top_core_KE_n3693) );
  OAI2BB2X1 U24405 ( .B0(n1431), .B1(n2039), .A0N(top_core_KE_key_mem_10__68_), 
        .A1N(n2042), .Y(top_core_KE_n4080) );
  OAI2BB2X1 U24406 ( .B0(n1431), .B1(n2058), .A0N(top_core_KE_key_mem_11__68_), 
        .A1N(n2068), .Y(top_core_KE_n4209) );
  OAI2BB2X1 U24407 ( .B0(n1431), .B1(n2078), .A0N(top_core_KE_key_mem_12__68_), 
        .A1N(n2088), .Y(top_core_KE_n4338) );
  OAI2BB2X1 U24408 ( .B0(n1431), .B1(n2098), .A0N(top_core_KE_key_mem_13__68_), 
        .A1N(n2108), .Y(top_core_KE_n4467) );
  OAI2BB2X1 U24409 ( .B0(n1431), .B1(n2118), .A0N(top_core_KE_key_mem_14__68_), 
        .A1N(n2128), .Y(top_core_KE_n4596) );
  OAI2BB2X1 U24410 ( .B0(n1422), .B1(n1859), .A0N(top_core_KE_key_mem_1__77_), 
        .A1N(n1871), .Y(top_core_KE_n2910) );
  OAI2BB2X1 U24411 ( .B0(n1422), .B1(n1878), .A0N(top_core_KE_key_mem_2__77_), 
        .A1N(n1889), .Y(top_core_KE_n3039) );
  OAI2BB2X1 U24412 ( .B0(n1422), .B1(n1898), .A0N(top_core_KE_key_mem_3__77_), 
        .A1N(n1908), .Y(top_core_KE_n3168) );
  OAI2BB2X1 U24413 ( .B0(n1422), .B1(n1918), .A0N(top_core_KE_key_mem_4__77_), 
        .A1N(n1929), .Y(top_core_KE_n3297) );
  OAI2BB2X1 U24414 ( .B0(n1422), .B1(n1944), .A0N(top_core_KE_key_mem_5__77_), 
        .A1N(n1948), .Y(top_core_KE_n3426) );
  OAI2BB2X1 U24415 ( .B0(n1422), .B1(n1958), .A0N(top_core_KE_key_mem_6__77_), 
        .A1N(n1968), .Y(top_core_KE_n3555) );
  OAI2BB2X1 U24416 ( .B0(n1422), .B1(n1977), .A0N(top_core_KE_key_mem_7__77_), 
        .A1N(n1988), .Y(top_core_KE_n3684) );
  OAI2BB2X1 U24417 ( .B0(n1422), .B1(n2038), .A0N(top_core_KE_key_mem_10__77_), 
        .A1N(n2043), .Y(top_core_KE_n4071) );
  OAI2BB2X1 U24418 ( .B0(n1422), .B1(n2057), .A0N(top_core_KE_key_mem_11__77_), 
        .A1N(n2068), .Y(top_core_KE_n4200) );
  OAI2BB2X1 U24419 ( .B0(n1422), .B1(n2084), .A0N(top_core_KE_key_mem_12__77_), 
        .A1N(n2088), .Y(top_core_KE_n4329) );
  OAI2BB2X1 U24420 ( .B0(n1422), .B1(n2097), .A0N(top_core_KE_key_mem_13__77_), 
        .A1N(n2108), .Y(top_core_KE_n4458) );
  OAI2BB2X1 U24421 ( .B0(n1422), .B1(n2117), .A0N(top_core_KE_key_mem_14__77_), 
        .A1N(n2128), .Y(top_core_KE_n4587) );
  OAI2BB2X1 U24422 ( .B0(n1430), .B1(n1860), .A0N(top_core_KE_key_mem_1__69_), 
        .A1N(n1872), .Y(top_core_KE_n2918) );
  OAI2BB2X1 U24423 ( .B0(n1430), .B1(n1879), .A0N(top_core_KE_key_mem_2__69_), 
        .A1N(n1889), .Y(top_core_KE_n3047) );
  OAI2BB2X1 U24424 ( .B0(n1430), .B1(n1907), .A0N(top_core_KE_key_mem_3__69_), 
        .A1N(n1908), .Y(top_core_KE_n3176) );
  OAI2BB2X1 U24425 ( .B0(n1430), .B1(n1919), .A0N(top_core_KE_key_mem_4__69_), 
        .A1N(n1929), .Y(top_core_KE_n3305) );
  OAI2BB2X1 U24426 ( .B0(n1430), .B1(n1938), .A0N(top_core_KE_key_mem_5__69_), 
        .A1N(n1948), .Y(top_core_KE_n3434) );
  OAI2BB2X1 U24427 ( .B0(n1430), .B1(n1959), .A0N(top_core_KE_key_mem_6__69_), 
        .A1N(n1968), .Y(top_core_KE_n3563) );
  OAI2BB2X1 U24428 ( .B0(n1430), .B1(n1978), .A0N(top_core_KE_key_mem_7__69_), 
        .A1N(n1988), .Y(top_core_KE_n3692) );
  OAI2BB2X1 U24429 ( .B0(n1430), .B1(n2039), .A0N(top_core_KE_key_mem_10__69_), 
        .A1N(n2041), .Y(top_core_KE_n4079) );
  OAI2BB2X1 U24430 ( .B0(n1430), .B1(n2058), .A0N(top_core_KE_key_mem_11__69_), 
        .A1N(n2068), .Y(top_core_KE_n4208) );
  OAI2BB2X1 U24431 ( .B0(n1430), .B1(n2078), .A0N(top_core_KE_key_mem_12__69_), 
        .A1N(n2088), .Y(top_core_KE_n4337) );
  OAI2BB2X1 U24432 ( .B0(n1430), .B1(n2098), .A0N(top_core_KE_key_mem_13__69_), 
        .A1N(n2108), .Y(top_core_KE_n4466) );
  OAI2BB2X1 U24433 ( .B0(n1430), .B1(n2118), .A0N(top_core_KE_key_mem_14__69_), 
        .A1N(n2128), .Y(top_core_KE_n4595) );
  OAI2BB2X1 U24434 ( .B0(n1419), .B1(n1859), .A0N(top_core_KE_key_mem_1__80_), 
        .A1N(n1870), .Y(top_core_KE_n2907) );
  OAI2BB2X1 U24435 ( .B0(n1419), .B1(n1877), .A0N(top_core_KE_key_mem_2__80_), 
        .A1N(n1889), .Y(top_core_KE_n3036) );
  OAI2BB2X1 U24436 ( .B0(n1419), .B1(n1897), .A0N(top_core_KE_key_mem_3__80_), 
        .A1N(n1908), .Y(top_core_KE_n3165) );
  OAI2BB2X1 U24437 ( .B0(n1419), .B1(n1917), .A0N(top_core_KE_key_mem_4__80_), 
        .A1N(n1929), .Y(top_core_KE_n3294) );
  OAI2BB2X1 U24438 ( .B0(n1419), .B1(n1937), .A0N(top_core_KE_key_mem_5__80_), 
        .A1N(n1948), .Y(top_core_KE_n3423) );
  OAI2BB2X1 U24439 ( .B0(n1419), .B1(n1957), .A0N(top_core_KE_key_mem_6__80_), 
        .A1N(n1968), .Y(top_core_KE_n3552) );
  OAI2BB2X1 U24440 ( .B0(n1419), .B1(n1992), .A0N(top_core_KE_key_mem_7__80_), 
        .A1N(n1988), .Y(top_core_KE_n3681) );
  OAI2BB2X1 U24441 ( .B0(n1419), .B1(n2037), .A0N(top_core_KE_key_mem_10__80_), 
        .A1N(n2038), .Y(top_core_KE_n4068) );
  OAI2BB2X1 U24442 ( .B0(n1419), .B1(n2072), .A0N(top_core_KE_key_mem_11__80_), 
        .A1N(n2068), .Y(top_core_KE_n4197) );
  OAI2BB2X1 U24443 ( .B0(n1419), .B1(n2077), .A0N(top_core_KE_key_mem_12__80_), 
        .A1N(n2088), .Y(top_core_KE_n4326) );
  OAI2BB2X1 U24444 ( .B0(n1419), .B1(n2112), .A0N(top_core_KE_key_mem_13__80_), 
        .A1N(n2108), .Y(top_core_KE_n4455) );
  OAI2BB2X1 U24445 ( .B0(n1419), .B1(n2132), .A0N(top_core_KE_key_mem_14__80_), 
        .A1N(n2128), .Y(top_core_KE_n4584) );
  OAI2BB2X1 U24446 ( .B0(n1387), .B1(n1857), .A0N(top_core_KE_key_mem_1__112_), 
        .A1N(n1867), .Y(top_core_KE_n2875) );
  OAI2BB2X1 U24447 ( .B0(n1387), .B1(n1882), .A0N(top_core_KE_key_mem_2__112_), 
        .A1N(n1885), .Y(top_core_KE_n3004) );
  OAI2BB2X1 U24448 ( .B0(n1387), .B1(n1901), .A0N(top_core_KE_key_mem_3__112_), 
        .A1N(n1904), .Y(top_core_KE_n3133) );
  OAI2BB2X1 U24449 ( .B0(n1387), .B1(n1922), .A0N(top_core_KE_key_mem_4__112_), 
        .A1N(n1925), .Y(top_core_KE_n3262) );
  OAI2BB2X1 U24450 ( .B0(n1387), .B1(n1941), .A0N(top_core_KE_key_mem_5__112_), 
        .A1N(n1944), .Y(top_core_KE_n3391) );
  OAI2BB2X1 U24451 ( .B0(n1387), .B1(n1962), .A0N(top_core_KE_key_mem_6__112_), 
        .A1N(n1965), .Y(top_core_KE_n3520) );
  OAI2BB2X1 U24452 ( .B0(n1387), .B1(n1981), .A0N(top_core_KE_key_mem_7__112_), 
        .A1N(n1984), .Y(top_core_KE_n3649) );
  OAI2BB2X1 U24453 ( .B0(n1387), .B1(n2042), .A0N(top_core_KE_key_mem_10__112_), .A1N(n2045), .Y(top_core_KE_n4036) );
  OAI2BB2X1 U24454 ( .B0(n1387), .B1(n2061), .A0N(top_core_KE_key_mem_11__112_), .A1N(n2064), .Y(top_core_KE_n4165) );
  OAI2BB2X1 U24455 ( .B0(n1387), .B1(n2081), .A0N(top_core_KE_key_mem_12__112_), .A1N(n2084), .Y(top_core_KE_n4294) );
  OAI2BB2X1 U24456 ( .B0(n1387), .B1(n2101), .A0N(top_core_KE_key_mem_13__112_), .A1N(n2104), .Y(top_core_KE_n4423) );
  OAI2BB2X1 U24457 ( .B0(n1387), .B1(n2121), .A0N(top_core_KE_key_mem_14__112_), .A1N(n2124), .Y(top_core_KE_n4552) );
  OAI2BB2X1 U24458 ( .B0(n1418), .B1(n1859), .A0N(top_core_KE_key_mem_1__81_), 
        .A1N(n1870), .Y(top_core_KE_n2906) );
  OAI2BB2X1 U24459 ( .B0(n1418), .B1(n1877), .A0N(top_core_KE_key_mem_2__81_), 
        .A1N(n1889), .Y(top_core_KE_n3035) );
  OAI2BB2X1 U24460 ( .B0(n1418), .B1(n1897), .A0N(top_core_KE_key_mem_3__81_), 
        .A1N(n1908), .Y(top_core_KE_n3164) );
  OAI2BB2X1 U24461 ( .B0(n1418), .B1(n1917), .A0N(top_core_KE_key_mem_4__81_), 
        .A1N(n1929), .Y(top_core_KE_n3293) );
  OAI2BB2X1 U24462 ( .B0(n1418), .B1(n1937), .A0N(top_core_KE_key_mem_5__81_), 
        .A1N(n1948), .Y(top_core_KE_n3422) );
  OAI2BB2X1 U24463 ( .B0(n1418), .B1(n1957), .A0N(top_core_KE_key_mem_6__81_), 
        .A1N(n1968), .Y(top_core_KE_n3551) );
  OAI2BB2X1 U24464 ( .B0(n1418), .B1(n1986), .A0N(top_core_KE_key_mem_7__81_), 
        .A1N(n1988), .Y(top_core_KE_n3680) );
  OAI2BB2X1 U24465 ( .B0(n1418), .B1(n2037), .A0N(top_core_KE_key_mem_10__81_), 
        .A1N(n2040), .Y(top_core_KE_n4067) );
  OAI2BB2X1 U24466 ( .B0(n1418), .B1(n2066), .A0N(top_core_KE_key_mem_11__81_), 
        .A1N(n2068), .Y(top_core_KE_n4196) );
  OAI2BB2X1 U24467 ( .B0(n1418), .B1(n2077), .A0N(top_core_KE_key_mem_12__81_), 
        .A1N(n2088), .Y(top_core_KE_n4325) );
  OAI2BB2X1 U24468 ( .B0(n1418), .B1(n2106), .A0N(top_core_KE_key_mem_13__81_), 
        .A1N(n2108), .Y(top_core_KE_n4454) );
  OAI2BB2X1 U24469 ( .B0(n1418), .B1(n2126), .A0N(top_core_KE_key_mem_14__81_), 
        .A1N(n2128), .Y(top_core_KE_n4583) );
  OAI2BB2X1 U24470 ( .B0(n1386), .B1(n1857), .A0N(top_core_KE_key_mem_1__113_), 
        .A1N(n1867), .Y(top_core_KE_n2874) );
  OAI2BB2X1 U24471 ( .B0(n1386), .B1(n1883), .A0N(top_core_KE_key_mem_2__113_), 
        .A1N(n1887), .Y(top_core_KE_n3003) );
  OAI2BB2X1 U24472 ( .B0(n1386), .B1(n1902), .A0N(top_core_KE_key_mem_3__113_), 
        .A1N(n1906), .Y(top_core_KE_n3132) );
  OAI2BB2X1 U24473 ( .B0(n1386), .B1(n1923), .A0N(top_core_KE_key_mem_4__113_), 
        .A1N(n1927), .Y(top_core_KE_n3261) );
  OAI2BB2X1 U24474 ( .B0(n1386), .B1(n1942), .A0N(top_core_KE_key_mem_5__113_), 
        .A1N(n1946), .Y(top_core_KE_n3390) );
  OAI2BB2X1 U24475 ( .B0(n1386), .B1(n1963), .A0N(top_core_KE_key_mem_6__113_), 
        .A1N(n1967), .Y(top_core_KE_n3519) );
  OAI2BB2X1 U24476 ( .B0(n1386), .B1(n1982), .A0N(top_core_KE_key_mem_7__113_), 
        .A1N(n1986), .Y(top_core_KE_n3648) );
  OAI2BB2X1 U24477 ( .B0(n1386), .B1(n2043), .A0N(top_core_KE_key_mem_10__113_), .A1N(n2047), .Y(top_core_KE_n4035) );
  OAI2BB2X1 U24478 ( .B0(n1386), .B1(n2062), .A0N(top_core_KE_key_mem_11__113_), .A1N(n2066), .Y(top_core_KE_n4164) );
  OAI2BB2X1 U24479 ( .B0(n1386), .B1(n2082), .A0N(top_core_KE_key_mem_12__113_), .A1N(n2086), .Y(top_core_KE_n4293) );
  OAI2BB2X1 U24480 ( .B0(n1386), .B1(n2102), .A0N(top_core_KE_key_mem_13__113_), .A1N(n2106), .Y(top_core_KE_n4422) );
  OAI2BB2X1 U24481 ( .B0(n1386), .B1(n2122), .A0N(top_core_KE_key_mem_14__113_), .A1N(n2126), .Y(top_core_KE_n4551) );
  OAI2BB2X1 U24482 ( .B0(n1417), .B1(n1859), .A0N(top_core_KE_key_mem_1__82_), 
        .A1N(n1870), .Y(top_core_KE_n2905) );
  OAI2BB2X1 U24483 ( .B0(n1417), .B1(n1877), .A0N(top_core_KE_key_mem_2__82_), 
        .A1N(n1888), .Y(top_core_KE_n3034) );
  OAI2BB2X1 U24484 ( .B0(n1417), .B1(n1897), .A0N(top_core_KE_key_mem_3__82_), 
        .A1N(n1907), .Y(top_core_KE_n3163) );
  OAI2BB2X1 U24485 ( .B0(n1417), .B1(n1917), .A0N(top_core_KE_key_mem_4__82_), 
        .A1N(n1928), .Y(top_core_KE_n3292) );
  OAI2BB2X1 U24486 ( .B0(n1417), .B1(n1937), .A0N(top_core_KE_key_mem_5__82_), 
        .A1N(n1947), .Y(top_core_KE_n3421) );
  OAI2BB2X1 U24487 ( .B0(n1417), .B1(n1957), .A0N(top_core_KE_key_mem_6__82_), 
        .A1N(n1966), .Y(top_core_KE_n3550) );
  OAI2BB2X1 U24488 ( .B0(n1417), .B1(n1991), .A0N(top_core_KE_key_mem_7__82_), 
        .A1N(n1987), .Y(top_core_KE_n3679) );
  OAI2BB2X1 U24489 ( .B0(n1417), .B1(n2037), .A0N(top_core_KE_key_mem_10__82_), 
        .A1N(n2048), .Y(top_core_KE_n4066) );
  OAI2BB2X1 U24490 ( .B0(n1417), .B1(n2071), .A0N(top_core_KE_key_mem_11__82_), 
        .A1N(n2067), .Y(top_core_KE_n4195) );
  OAI2BB2X1 U24491 ( .B0(n1417), .B1(n2077), .A0N(top_core_KE_key_mem_12__82_), 
        .A1N(n2087), .Y(top_core_KE_n4324) );
  OAI2BB2X1 U24492 ( .B0(n1417), .B1(n2111), .A0N(top_core_KE_key_mem_13__82_), 
        .A1N(n2107), .Y(top_core_KE_n4453) );
  OAI2BB2X1 U24493 ( .B0(n1417), .B1(n2131), .A0N(top_core_KE_key_mem_14__82_), 
        .A1N(n2127), .Y(top_core_KE_n4582) );
  OAI2BB2X1 U24494 ( .B0(n1385), .B1(n1857), .A0N(top_core_KE_key_mem_1__114_), 
        .A1N(n1867), .Y(top_core_KE_n2873) );
  OAI2BB2X1 U24495 ( .B0(n1385), .B1(n1883), .A0N(top_core_KE_key_mem_2__114_), 
        .A1N(n1886), .Y(top_core_KE_n3002) );
  OAI2BB2X1 U24496 ( .B0(n1385), .B1(n1902), .A0N(top_core_KE_key_mem_3__114_), 
        .A1N(n1905), .Y(top_core_KE_n3131) );
  OAI2BB2X1 U24497 ( .B0(n1385), .B1(n1923), .A0N(top_core_KE_key_mem_4__114_), 
        .A1N(n1926), .Y(top_core_KE_n3260) );
  OAI2BB2X1 U24498 ( .B0(n1385), .B1(n1942), .A0N(top_core_KE_key_mem_5__114_), 
        .A1N(n1945), .Y(top_core_KE_n3389) );
  OAI2BB2X1 U24499 ( .B0(n1385), .B1(n1963), .A0N(top_core_KE_key_mem_6__114_), 
        .A1N(n1966), .Y(top_core_KE_n3518) );
  OAI2BB2X1 U24500 ( .B0(n1385), .B1(n1982), .A0N(top_core_KE_key_mem_7__114_), 
        .A1N(n1985), .Y(top_core_KE_n3647) );
  OAI2BB2X1 U24501 ( .B0(n1385), .B1(n2043), .A0N(top_core_KE_key_mem_10__114_), .A1N(n2046), .Y(top_core_KE_n4034) );
  OAI2BB2X1 U24502 ( .B0(n1385), .B1(n2062), .A0N(top_core_KE_key_mem_11__114_), .A1N(n2065), .Y(top_core_KE_n4163) );
  OAI2BB2X1 U24503 ( .B0(n1385), .B1(n2082), .A0N(top_core_KE_key_mem_12__114_), .A1N(n2085), .Y(top_core_KE_n4292) );
  OAI2BB2X1 U24504 ( .B0(n1385), .B1(n2102), .A0N(top_core_KE_key_mem_13__114_), .A1N(n2105), .Y(top_core_KE_n4421) );
  OAI2BB2X1 U24505 ( .B0(n1385), .B1(n2122), .A0N(top_core_KE_key_mem_14__114_), .A1N(n2125), .Y(top_core_KE_n4550) );
  OAI2BB2X1 U24506 ( .B0(n1416), .B1(n1859), .A0N(top_core_KE_key_mem_1__83_), 
        .A1N(n1870), .Y(top_core_KE_n2904) );
  OAI2BB2X1 U24507 ( .B0(n1416), .B1(n1877), .A0N(top_core_KE_key_mem_2__83_), 
        .A1N(n1888), .Y(top_core_KE_n3033) );
  OAI2BB2X1 U24508 ( .B0(n1416), .B1(n1897), .A0N(top_core_KE_key_mem_3__83_), 
        .A1N(n1907), .Y(top_core_KE_n3162) );
  OAI2BB2X1 U24509 ( .B0(n1416), .B1(n1917), .A0N(top_core_KE_key_mem_4__83_), 
        .A1N(n1928), .Y(top_core_KE_n3291) );
  OAI2BB2X1 U24510 ( .B0(n1416), .B1(n1937), .A0N(top_core_KE_key_mem_5__83_), 
        .A1N(n1947), .Y(top_core_KE_n3420) );
  OAI2BB2X1 U24511 ( .B0(n1416), .B1(n1957), .A0N(top_core_KE_key_mem_6__83_), 
        .A1N(n1970), .Y(top_core_KE_n3549) );
  OAI2BB2X1 U24512 ( .B0(n1416), .B1(n1984), .A0N(top_core_KE_key_mem_7__83_), 
        .A1N(n1987), .Y(top_core_KE_n3678) );
  OAI2BB2X1 U24513 ( .B0(n1416), .B1(n2037), .A0N(top_core_KE_key_mem_10__83_), 
        .A1N(n2048), .Y(top_core_KE_n4065) );
  OAI2BB2X1 U24514 ( .B0(n1416), .B1(n2064), .A0N(top_core_KE_key_mem_11__83_), 
        .A1N(n2067), .Y(top_core_KE_n4194) );
  OAI2BB2X1 U24515 ( .B0(n1416), .B1(n2077), .A0N(top_core_KE_key_mem_12__83_), 
        .A1N(n2087), .Y(top_core_KE_n4323) );
  OAI2BB2X1 U24516 ( .B0(n1416), .B1(n2104), .A0N(top_core_KE_key_mem_13__83_), 
        .A1N(n2107), .Y(top_core_KE_n4452) );
  OAI2BB2X1 U24517 ( .B0(n1416), .B1(n2124), .A0N(top_core_KE_key_mem_14__83_), 
        .A1N(n2127), .Y(top_core_KE_n4581) );
  OAI2BB2X1 U24518 ( .B0(n1384), .B1(n1857), .A0N(top_core_KE_key_mem_1__115_), 
        .A1N(n1867), .Y(top_core_KE_n2872) );
  OAI2BB2X1 U24519 ( .B0(n1384), .B1(n1883), .A0N(top_core_KE_key_mem_2__115_), 
        .A1N(n1886), .Y(top_core_KE_n3001) );
  OAI2BB2X1 U24520 ( .B0(n1384), .B1(n1902), .A0N(top_core_KE_key_mem_3__115_), 
        .A1N(n1905), .Y(top_core_KE_n3130) );
  OAI2BB2X1 U24521 ( .B0(n1384), .B1(n1923), .A0N(top_core_KE_key_mem_4__115_), 
        .A1N(n1926), .Y(top_core_KE_n3259) );
  OAI2BB2X1 U24522 ( .B0(n1384), .B1(n1942), .A0N(top_core_KE_key_mem_5__115_), 
        .A1N(n1945), .Y(top_core_KE_n3388) );
  OAI2BB2X1 U24523 ( .B0(n1384), .B1(n1963), .A0N(top_core_KE_key_mem_6__115_), 
        .A1N(n1966), .Y(top_core_KE_n3517) );
  OAI2BB2X1 U24524 ( .B0(n1384), .B1(n1982), .A0N(top_core_KE_key_mem_7__115_), 
        .A1N(n1985), .Y(top_core_KE_n3646) );
  OAI2BB2X1 U24525 ( .B0(n1384), .B1(n2043), .A0N(top_core_KE_key_mem_10__115_), .A1N(n2046), .Y(top_core_KE_n4033) );
  OAI2BB2X1 U24526 ( .B0(n1384), .B1(n2062), .A0N(top_core_KE_key_mem_11__115_), .A1N(n2065), .Y(top_core_KE_n4162) );
  OAI2BB2X1 U24527 ( .B0(n1384), .B1(n2082), .A0N(top_core_KE_key_mem_12__115_), .A1N(n2085), .Y(top_core_KE_n4291) );
  OAI2BB2X1 U24528 ( .B0(n1384), .B1(n2102), .A0N(top_core_KE_key_mem_13__115_), .A1N(n2105), .Y(top_core_KE_n4420) );
  OAI2BB2X1 U24529 ( .B0(n1384), .B1(n2122), .A0N(top_core_KE_key_mem_14__115_), .A1N(n2125), .Y(top_core_KE_n4549) );
  OAI2BB2X1 U24530 ( .B0(n1415), .B1(n1859), .A0N(top_core_KE_key_mem_1__84_), 
        .A1N(n1870), .Y(top_core_KE_n2903) );
  OAI2BB2X1 U24531 ( .B0(n1415), .B1(n1877), .A0N(top_core_KE_key_mem_2__84_), 
        .A1N(n1888), .Y(top_core_KE_n3032) );
  OAI2BB2X1 U24532 ( .B0(n1415), .B1(n1897), .A0N(top_core_KE_key_mem_3__84_), 
        .A1N(n1907), .Y(top_core_KE_n3161) );
  OAI2BB2X1 U24533 ( .B0(n1415), .B1(n1917), .A0N(top_core_KE_key_mem_4__84_), 
        .A1N(n1928), .Y(top_core_KE_n3290) );
  OAI2BB2X1 U24534 ( .B0(n1415), .B1(n1937), .A0N(top_core_KE_key_mem_5__84_), 
        .A1N(n1947), .Y(top_core_KE_n3419) );
  OAI2BB2X1 U24535 ( .B0(n1415), .B1(n1957), .A0N(top_core_KE_key_mem_6__84_), 
        .A1N(n1971), .Y(top_core_KE_n3548) );
  OAI2BB2X1 U24536 ( .B0(n1415), .B1(n1981), .A0N(top_core_KE_key_mem_7__84_), 
        .A1N(n1987), .Y(top_core_KE_n3677) );
  OAI2BB2X1 U24537 ( .B0(n1415), .B1(n2037), .A0N(top_core_KE_key_mem_10__84_), 
        .A1N(n2048), .Y(top_core_KE_n4064) );
  OAI2BB2X1 U24538 ( .B0(n1415), .B1(n2061), .A0N(top_core_KE_key_mem_11__84_), 
        .A1N(n2067), .Y(top_core_KE_n4193) );
  OAI2BB2X1 U24539 ( .B0(n1415), .B1(n2077), .A0N(top_core_KE_key_mem_12__84_), 
        .A1N(n2087), .Y(top_core_KE_n4322) );
  OAI2BB2X1 U24540 ( .B0(n1415), .B1(n2101), .A0N(top_core_KE_key_mem_13__84_), 
        .A1N(n2107), .Y(top_core_KE_n4451) );
  OAI2BB2X1 U24541 ( .B0(n1415), .B1(n2121), .A0N(top_core_KE_key_mem_14__84_), 
        .A1N(n2127), .Y(top_core_KE_n4580) );
  OAI2BB2X1 U24542 ( .B0(n1383), .B1(n1863), .A0N(top_core_KE_key_mem_1__116_), 
        .A1N(n1867), .Y(top_core_KE_n2871) );
  OAI2BB2X1 U24543 ( .B0(n1383), .B1(n1883), .A0N(top_core_KE_key_mem_2__116_), 
        .A1N(n1887), .Y(top_core_KE_n3000) );
  OAI2BB2X1 U24544 ( .B0(n1383), .B1(n1902), .A0N(top_core_KE_key_mem_3__116_), 
        .A1N(n1906), .Y(top_core_KE_n3129) );
  OAI2BB2X1 U24545 ( .B0(n1383), .B1(n1923), .A0N(top_core_KE_key_mem_4__116_), 
        .A1N(n1927), .Y(top_core_KE_n3258) );
  OAI2BB2X1 U24546 ( .B0(n1383), .B1(n1942), .A0N(top_core_KE_key_mem_5__116_), 
        .A1N(n1946), .Y(top_core_KE_n3387) );
  OAI2BB2X1 U24547 ( .B0(n1383), .B1(n1963), .A0N(top_core_KE_key_mem_6__116_), 
        .A1N(n1967), .Y(top_core_KE_n3516) );
  OAI2BB2X1 U24548 ( .B0(n1383), .B1(n1982), .A0N(top_core_KE_key_mem_7__116_), 
        .A1N(n1986), .Y(top_core_KE_n3645) );
  OAI2BB2X1 U24549 ( .B0(n1383), .B1(n2043), .A0N(top_core_KE_key_mem_10__116_), .A1N(n2047), .Y(top_core_KE_n4032) );
  OAI2BB2X1 U24550 ( .B0(n1383), .B1(n2062), .A0N(top_core_KE_key_mem_11__116_), .A1N(n2066), .Y(top_core_KE_n4161) );
  OAI2BB2X1 U24551 ( .B0(n1383), .B1(n2082), .A0N(top_core_KE_key_mem_12__116_), .A1N(n2086), .Y(top_core_KE_n4290) );
  OAI2BB2X1 U24552 ( .B0(n1383), .B1(n2102), .A0N(top_core_KE_key_mem_13__116_), .A1N(n2106), .Y(top_core_KE_n4419) );
  OAI2BB2X1 U24553 ( .B0(n1383), .B1(n2122), .A0N(top_core_KE_key_mem_14__116_), .A1N(n2126), .Y(top_core_KE_n4548) );
  OAI2BB2X1 U24554 ( .B0(n1414), .B1(n1859), .A0N(top_core_KE_key_mem_1__85_), 
        .A1N(n1870), .Y(top_core_KE_n2902) );
  OAI2BB2X1 U24555 ( .B0(n1414), .B1(n1882), .A0N(top_core_KE_key_mem_2__85_), 
        .A1N(n1888), .Y(top_core_KE_n3031) );
  OAI2BB2X1 U24556 ( .B0(n1414), .B1(n1901), .A0N(top_core_KE_key_mem_3__85_), 
        .A1N(n1907), .Y(top_core_KE_n3160) );
  OAI2BB2X1 U24557 ( .B0(n1414), .B1(n1922), .A0N(top_core_KE_key_mem_4__85_), 
        .A1N(n1928), .Y(top_core_KE_n3289) );
  OAI2BB2X1 U24558 ( .B0(n1414), .B1(n1941), .A0N(top_core_KE_key_mem_5__85_), 
        .A1N(n1947), .Y(top_core_KE_n3418) );
  OAI2BB2X1 U24559 ( .B0(n1414), .B1(n1962), .A0N(top_core_KE_key_mem_6__85_), 
        .A1N(n1972), .Y(top_core_KE_n3547) );
  OAI2BB2X1 U24560 ( .B0(n1414), .B1(n1981), .A0N(top_core_KE_key_mem_7__85_), 
        .A1N(n1987), .Y(top_core_KE_n3676) );
  OAI2BB2X1 U24561 ( .B0(n1414), .B1(n2042), .A0N(top_core_KE_key_mem_10__85_), 
        .A1N(n2048), .Y(top_core_KE_n4063) );
  OAI2BB2X1 U24562 ( .B0(n1414), .B1(n2061), .A0N(top_core_KE_key_mem_11__85_), 
        .A1N(n2067), .Y(top_core_KE_n4192) );
  OAI2BB2X1 U24563 ( .B0(n1414), .B1(n2081), .A0N(top_core_KE_key_mem_12__85_), 
        .A1N(n2087), .Y(top_core_KE_n4321) );
  OAI2BB2X1 U24564 ( .B0(n1414), .B1(n2101), .A0N(top_core_KE_key_mem_13__85_), 
        .A1N(n2107), .Y(top_core_KE_n4450) );
  OAI2BB2X1 U24565 ( .B0(n1414), .B1(n2121), .A0N(top_core_KE_key_mem_14__85_), 
        .A1N(n2127), .Y(top_core_KE_n4579) );
  OAI2BB2X1 U24566 ( .B0(n1382), .B1(n1860), .A0N(top_core_KE_key_mem_1__117_), 
        .A1N(n1866), .Y(top_core_KE_n2870) );
  OAI2BB2X1 U24567 ( .B0(n1382), .B1(n1883), .A0N(top_core_KE_key_mem_2__117_), 
        .A1N(n1886), .Y(top_core_KE_n2999) );
  OAI2BB2X1 U24568 ( .B0(n1382), .B1(n1902), .A0N(top_core_KE_key_mem_3__117_), 
        .A1N(n1905), .Y(top_core_KE_n3128) );
  OAI2BB2X1 U24569 ( .B0(n1382), .B1(n1923), .A0N(top_core_KE_key_mem_4__117_), 
        .A1N(n1926), .Y(top_core_KE_n3257) );
  OAI2BB2X1 U24570 ( .B0(n1382), .B1(n1942), .A0N(top_core_KE_key_mem_5__117_), 
        .A1N(n1945), .Y(top_core_KE_n3386) );
  OAI2BB2X1 U24571 ( .B0(n1382), .B1(n1963), .A0N(top_core_KE_key_mem_6__117_), 
        .A1N(n1966), .Y(top_core_KE_n3515) );
  OAI2BB2X1 U24572 ( .B0(n1382), .B1(n1982), .A0N(top_core_KE_key_mem_7__117_), 
        .A1N(n1985), .Y(top_core_KE_n3644) );
  OAI2BB2X1 U24573 ( .B0(n1382), .B1(n2043), .A0N(top_core_KE_key_mem_10__117_), .A1N(n2046), .Y(top_core_KE_n4031) );
  OAI2BB2X1 U24574 ( .B0(n1382), .B1(n2062), .A0N(top_core_KE_key_mem_11__117_), .A1N(n2065), .Y(top_core_KE_n4160) );
  OAI2BB2X1 U24575 ( .B0(n1382), .B1(n2082), .A0N(top_core_KE_key_mem_12__117_), .A1N(n2085), .Y(top_core_KE_n4289) );
  OAI2BB2X1 U24576 ( .B0(n1382), .B1(n2102), .A0N(top_core_KE_key_mem_13__117_), .A1N(n2105), .Y(top_core_KE_n4418) );
  OAI2BB2X1 U24577 ( .B0(n1382), .B1(n2122), .A0N(top_core_KE_key_mem_14__117_), .A1N(n2125), .Y(top_core_KE_n4547) );
  OAI2BB2X1 U24578 ( .B0(n1413), .B1(n1859), .A0N(top_core_KE_key_mem_1__86_), 
        .A1N(n1870), .Y(top_core_KE_n2901) );
  OAI2BB2X1 U24579 ( .B0(n1413), .B1(n1877), .A0N(top_core_KE_key_mem_2__86_), 
        .A1N(n1888), .Y(top_core_KE_n3030) );
  OAI2BB2X1 U24580 ( .B0(n1413), .B1(n1897), .A0N(top_core_KE_key_mem_3__86_), 
        .A1N(n1907), .Y(top_core_KE_n3159) );
  OAI2BB2X1 U24581 ( .B0(n1413), .B1(n1917), .A0N(top_core_KE_key_mem_4__86_), 
        .A1N(n1928), .Y(top_core_KE_n3288) );
  OAI2BB2X1 U24582 ( .B0(n1413), .B1(n1937), .A0N(top_core_KE_key_mem_5__86_), 
        .A1N(n1947), .Y(top_core_KE_n3417) );
  OAI2BB2X1 U24583 ( .B0(n1413), .B1(n1957), .A0N(top_core_KE_key_mem_6__86_), 
        .A1N(n1967), .Y(top_core_KE_n3546) );
  OAI2BB2X1 U24584 ( .B0(n1413), .B1(n1982), .A0N(top_core_KE_key_mem_7__86_), 
        .A1N(n1987), .Y(top_core_KE_n3675) );
  OAI2BB2X1 U24585 ( .B0(n1413), .B1(n2037), .A0N(top_core_KE_key_mem_10__86_), 
        .A1N(n2048), .Y(top_core_KE_n4062) );
  OAI2BB2X1 U24586 ( .B0(n1413), .B1(n2062), .A0N(top_core_KE_key_mem_11__86_), 
        .A1N(n2067), .Y(top_core_KE_n4191) );
  OAI2BB2X1 U24587 ( .B0(n1413), .B1(n2077), .A0N(top_core_KE_key_mem_12__86_), 
        .A1N(n2087), .Y(top_core_KE_n4320) );
  OAI2BB2X1 U24588 ( .B0(n1413), .B1(n2102), .A0N(top_core_KE_key_mem_13__86_), 
        .A1N(n2107), .Y(top_core_KE_n4449) );
  OAI2BB2X1 U24589 ( .B0(n1413), .B1(n2122), .A0N(top_core_KE_key_mem_14__86_), 
        .A1N(n2127), .Y(top_core_KE_n4578) );
  OAI2BB2X1 U24590 ( .B0(n1381), .B1(n1859), .A0N(top_core_KE_key_mem_1__118_), 
        .A1N(n1866), .Y(top_core_KE_n2869) );
  OAI2BB2X1 U24591 ( .B0(n1381), .B1(n1884), .A0N(top_core_KE_key_mem_2__118_), 
        .A1N(n1886), .Y(top_core_KE_n2998) );
  OAI2BB2X1 U24592 ( .B0(n1381), .B1(n1903), .A0N(top_core_KE_key_mem_3__118_), 
        .A1N(n1905), .Y(top_core_KE_n3127) );
  OAI2BB2X1 U24593 ( .B0(n1381), .B1(n1924), .A0N(top_core_KE_key_mem_4__118_), 
        .A1N(n1926), .Y(top_core_KE_n3256) );
  OAI2BB2X1 U24594 ( .B0(n1381), .B1(n1943), .A0N(top_core_KE_key_mem_5__118_), 
        .A1N(n1945), .Y(top_core_KE_n3385) );
  OAI2BB2X1 U24595 ( .B0(n1381), .B1(n1964), .A0N(top_core_KE_key_mem_6__118_), 
        .A1N(n1966), .Y(top_core_KE_n3514) );
  OAI2BB2X1 U24596 ( .B0(n1381), .B1(n1983), .A0N(top_core_KE_key_mem_7__118_), 
        .A1N(n1985), .Y(top_core_KE_n3643) );
  OAI2BB2X1 U24597 ( .B0(n1381), .B1(n2044), .A0N(top_core_KE_key_mem_10__118_), .A1N(n2046), .Y(top_core_KE_n4030) );
  OAI2BB2X1 U24598 ( .B0(n1381), .B1(n2063), .A0N(top_core_KE_key_mem_11__118_), .A1N(n2065), .Y(top_core_KE_n4159) );
  OAI2BB2X1 U24599 ( .B0(n1381), .B1(n2083), .A0N(top_core_KE_key_mem_12__118_), .A1N(n2085), .Y(top_core_KE_n4288) );
  OAI2BB2X1 U24600 ( .B0(n1381), .B1(n2103), .A0N(top_core_KE_key_mem_13__118_), .A1N(n2105), .Y(top_core_KE_n4417) );
  OAI2BB2X1 U24601 ( .B0(n1381), .B1(n2123), .A0N(top_core_KE_key_mem_14__118_), .A1N(n2125), .Y(top_core_KE_n4546) );
  OAI2BB2X1 U24602 ( .B0(n1421), .B1(n1859), .A0N(top_core_KE_key_mem_1__78_), 
        .A1N(n1871), .Y(top_core_KE_n2909) );
  OAI2BB2X1 U24603 ( .B0(n1421), .B1(n1877), .A0N(top_core_KE_key_mem_2__78_), 
        .A1N(n1889), .Y(top_core_KE_n3038) );
  OAI2BB2X1 U24604 ( .B0(n1421), .B1(n1897), .A0N(top_core_KE_key_mem_3__78_), 
        .A1N(n1908), .Y(top_core_KE_n3167) );
  OAI2BB2X1 U24605 ( .B0(n1421), .B1(n1917), .A0N(top_core_KE_key_mem_4__78_), 
        .A1N(n1929), .Y(top_core_KE_n3296) );
  OAI2BB2X1 U24606 ( .B0(n1421), .B1(n1937), .A0N(top_core_KE_key_mem_5__78_), 
        .A1N(n1948), .Y(top_core_KE_n3425) );
  OAI2BB2X1 U24607 ( .B0(n1421), .B1(n1957), .A0N(top_core_KE_key_mem_6__78_), 
        .A1N(n1968), .Y(top_core_KE_n3554) );
  OAI2BB2X1 U24608 ( .B0(n1421), .B1(n1987), .A0N(top_core_KE_key_mem_7__78_), 
        .A1N(n1988), .Y(top_core_KE_n3683) );
  OAI2BB2X1 U24609 ( .B0(n1421), .B1(n2037), .A0N(top_core_KE_key_mem_10__78_), 
        .A1N(n2039), .Y(top_core_KE_n4070) );
  OAI2BB2X1 U24610 ( .B0(n1421), .B1(n2067), .A0N(top_core_KE_key_mem_11__78_), 
        .A1N(n2068), .Y(top_core_KE_n4199) );
  OAI2BB2X1 U24611 ( .B0(n1421), .B1(n2077), .A0N(top_core_KE_key_mem_12__78_), 
        .A1N(n2088), .Y(top_core_KE_n4328) );
  OAI2BB2X1 U24612 ( .B0(n1421), .B1(n2107), .A0N(top_core_KE_key_mem_13__78_), 
        .A1N(n2108), .Y(top_core_KE_n4457) );
  OAI2BB2X1 U24613 ( .B0(n1421), .B1(n2127), .A0N(top_core_KE_key_mem_14__78_), 
        .A1N(n2128), .Y(top_core_KE_n4586) );
  OAI2BB2X1 U24614 ( .B0(n1429), .B1(n1860), .A0N(top_core_KE_key_mem_1__70_), 
        .A1N(n1871), .Y(top_core_KE_n2917) );
  OAI2BB2X1 U24615 ( .B0(n1429), .B1(n1878), .A0N(top_core_KE_key_mem_2__70_), 
        .A1N(n1889), .Y(top_core_KE_n3046) );
  OAI2BB2X1 U24616 ( .B0(n1429), .B1(n1898), .A0N(top_core_KE_key_mem_3__70_), 
        .A1N(n1908), .Y(top_core_KE_n3175) );
  OAI2BB2X1 U24617 ( .B0(n1429), .B1(n1918), .A0N(top_core_KE_key_mem_4__70_), 
        .A1N(n1929), .Y(top_core_KE_n3304) );
  OAI2BB2X1 U24618 ( .B0(n1429), .B1(n1940), .A0N(top_core_KE_key_mem_5__70_), 
        .A1N(n1948), .Y(top_core_KE_n3433) );
  OAI2BB2X1 U24619 ( .B0(n1429), .B1(n1958), .A0N(top_core_KE_key_mem_6__70_), 
        .A1N(n1968), .Y(top_core_KE_n3562) );
  OAI2BB2X1 U24620 ( .B0(n1429), .B1(n1977), .A0N(top_core_KE_key_mem_7__70_), 
        .A1N(n1988), .Y(top_core_KE_n3691) );
  OAI2BB2X1 U24621 ( .B0(n1429), .B1(n2038), .A0N(top_core_KE_key_mem_10__70_), 
        .A1N(n2037), .Y(top_core_KE_n4078) );
  OAI2BB2X1 U24622 ( .B0(n1429), .B1(n2057), .A0N(top_core_KE_key_mem_11__70_), 
        .A1N(n2068), .Y(top_core_KE_n4207) );
  OAI2BB2X1 U24623 ( .B0(n1429), .B1(n2080), .A0N(top_core_KE_key_mem_12__70_), 
        .A1N(n2088), .Y(top_core_KE_n4336) );
  OAI2BB2X1 U24624 ( .B0(n1429), .B1(n2097), .A0N(top_core_KE_key_mem_13__70_), 
        .A1N(n2108), .Y(top_core_KE_n4465) );
  OAI2BB2X1 U24625 ( .B0(n1429), .B1(n2117), .A0N(top_core_KE_key_mem_14__70_), 
        .A1N(n2128), .Y(top_core_KE_n4594) );
  OAI2BB2X1 U24626 ( .B0(n1372), .B1(n1864), .A0N(top_core_KE_key_mem_1__127_), 
        .A1N(n1866), .Y(top_core_KE_n2860) );
  OAI2BB2X1 U24627 ( .B0(n1372), .B1(n1885), .A0N(top_core_KE_key_mem_2__127_), 
        .A1N(n1888), .Y(top_core_KE_n2989) );
  OAI2BB2X1 U24628 ( .B0(n1372), .B1(n1904), .A0N(top_core_KE_key_mem_3__127_), 
        .A1N(n1907), .Y(top_core_KE_n3118) );
  OAI2BB2X1 U24629 ( .B0(n1372), .B1(n1925), .A0N(top_core_KE_key_mem_4__127_), 
        .A1N(n1928), .Y(top_core_KE_n3247) );
  OAI2BB2X1 U24630 ( .B0(n1372), .B1(n1944), .A0N(top_core_KE_key_mem_5__127_), 
        .A1N(n1947), .Y(top_core_KE_n3376) );
  OAI2BB2X1 U24631 ( .B0(n1372), .B1(n1965), .A0N(top_core_KE_key_mem_6__127_), 
        .A1N(n1965), .Y(top_core_KE_n3505) );
  OAI2BB2X1 U24632 ( .B0(n1372), .B1(n1984), .A0N(top_core_KE_key_mem_7__127_), 
        .A1N(n1987), .Y(top_core_KE_n3634) );
  OAI2BB2X1 U24633 ( .B0(n1372), .B1(n2045), .A0N(top_core_KE_key_mem_10__127_), .A1N(n2048), .Y(top_core_KE_n4021) );
  OAI2BB2X1 U24634 ( .B0(n1372), .B1(n2064), .A0N(top_core_KE_key_mem_11__127_), .A1N(n2067), .Y(top_core_KE_n4150) );
  OAI2BB2X1 U24635 ( .B0(n1372), .B1(n2084), .A0N(top_core_KE_key_mem_12__127_), .A1N(n2087), .Y(top_core_KE_n4279) );
  OAI2BB2X1 U24636 ( .B0(n1372), .B1(n2104), .A0N(top_core_KE_key_mem_13__127_), .A1N(n2107), .Y(top_core_KE_n4408) );
  OAI2BB2X1 U24637 ( .B0(n1372), .B1(n2124), .A0N(top_core_KE_key_mem_14__127_), .A1N(n2127), .Y(top_core_KE_n4537) );
  OAI2BB2X1 U24638 ( .B0(n1412), .B1(n1859), .A0N(top_core_KE_key_mem_1__87_), 
        .A1N(n1870), .Y(top_core_KE_n2900) );
  OAI2BB2X1 U24639 ( .B0(n1412), .B1(n1877), .A0N(top_core_KE_key_mem_2__87_), 
        .A1N(n1888), .Y(top_core_KE_n3029) );
  OAI2BB2X1 U24640 ( .B0(n1412), .B1(n1897), .A0N(top_core_KE_key_mem_3__87_), 
        .A1N(n1907), .Y(top_core_KE_n3158) );
  OAI2BB2X1 U24641 ( .B0(n1412), .B1(n1917), .A0N(top_core_KE_key_mem_4__87_), 
        .A1N(n1928), .Y(top_core_KE_n3287) );
  OAI2BB2X1 U24642 ( .B0(n1412), .B1(n1937), .A0N(top_core_KE_key_mem_5__87_), 
        .A1N(n1947), .Y(top_core_KE_n3416) );
  OAI2BB2X1 U24643 ( .B0(n1412), .B1(n1957), .A0N(top_core_KE_key_mem_6__87_), 
        .A1N(n1962), .Y(top_core_KE_n3545) );
  OAI2BB2X1 U24644 ( .B0(n1412), .B1(n1980), .A0N(top_core_KE_key_mem_7__87_), 
        .A1N(n1987), .Y(top_core_KE_n3674) );
  OAI2BB2X1 U24645 ( .B0(n1412), .B1(n2037), .A0N(top_core_KE_key_mem_10__87_), 
        .A1N(n2048), .Y(top_core_KE_n4061) );
  OAI2BB2X1 U24646 ( .B0(n1412), .B1(n2060), .A0N(top_core_KE_key_mem_11__87_), 
        .A1N(n2067), .Y(top_core_KE_n4190) );
  OAI2BB2X1 U24647 ( .B0(n1412), .B1(n2077), .A0N(top_core_KE_key_mem_12__87_), 
        .A1N(n2087), .Y(top_core_KE_n4319) );
  OAI2BB2X1 U24648 ( .B0(n1412), .B1(n2100), .A0N(top_core_KE_key_mem_13__87_), 
        .A1N(n2107), .Y(top_core_KE_n4448) );
  OAI2BB2X1 U24649 ( .B0(n1412), .B1(n2120), .A0N(top_core_KE_key_mem_14__87_), 
        .A1N(n2127), .Y(top_core_KE_n4577) );
  OAI2BB2X1 U24650 ( .B0(n1380), .B1(n1862), .A0N(top_core_KE_key_mem_1__119_), 
        .A1N(n1867), .Y(top_core_KE_n2868) );
  OAI2BB2X1 U24651 ( .B0(n1380), .B1(n1884), .A0N(top_core_KE_key_mem_2__119_), 
        .A1N(n1888), .Y(top_core_KE_n2997) );
  OAI2BB2X1 U24652 ( .B0(n1380), .B1(n1903), .A0N(top_core_KE_key_mem_3__119_), 
        .A1N(n1907), .Y(top_core_KE_n3126) );
  OAI2BB2X1 U24653 ( .B0(n1380), .B1(n1924), .A0N(top_core_KE_key_mem_4__119_), 
        .A1N(n1928), .Y(top_core_KE_n3255) );
  OAI2BB2X1 U24654 ( .B0(n1380), .B1(n1943), .A0N(top_core_KE_key_mem_5__119_), 
        .A1N(n1947), .Y(top_core_KE_n3384) );
  OAI2BB2X1 U24655 ( .B0(n1380), .B1(n1964), .A0N(top_core_KE_key_mem_6__119_), 
        .A1N(n1963), .Y(top_core_KE_n3513) );
  OAI2BB2X1 U24656 ( .B0(n1380), .B1(n1983), .A0N(top_core_KE_key_mem_7__119_), 
        .A1N(n1987), .Y(top_core_KE_n3642) );
  OAI2BB2X1 U24657 ( .B0(n1380), .B1(n2044), .A0N(top_core_KE_key_mem_10__119_), .A1N(n2048), .Y(top_core_KE_n4029) );
  OAI2BB2X1 U24658 ( .B0(n1380), .B1(n2063), .A0N(top_core_KE_key_mem_11__119_), .A1N(n2067), .Y(top_core_KE_n4158) );
  OAI2BB2X1 U24659 ( .B0(n1380), .B1(n2083), .A0N(top_core_KE_key_mem_12__119_), .A1N(n2087), .Y(top_core_KE_n4287) );
  OAI2BB2X1 U24660 ( .B0(n1380), .B1(n2103), .A0N(top_core_KE_key_mem_13__119_), .A1N(n2107), .Y(top_core_KE_n4416) );
  OAI2BB2X1 U24661 ( .B0(n1380), .B1(n2123), .A0N(top_core_KE_key_mem_14__119_), .A1N(n2127), .Y(top_core_KE_n4545) );
  OAI2BB2X1 U24662 ( .B0(n1420), .B1(n1859), .A0N(top_core_KE_key_mem_1__79_), 
        .A1N(n1871), .Y(top_core_KE_n2908) );
  OAI2BB2X1 U24663 ( .B0(n1420), .B1(n1877), .A0N(top_core_KE_key_mem_2__79_), 
        .A1N(n1889), .Y(top_core_KE_n3037) );
  OAI2BB2X1 U24664 ( .B0(n1420), .B1(n1897), .A0N(top_core_KE_key_mem_3__79_), 
        .A1N(n1908), .Y(top_core_KE_n3166) );
  OAI2BB2X1 U24665 ( .B0(n1420), .B1(n1917), .A0N(top_core_KE_key_mem_4__79_), 
        .A1N(n1929), .Y(top_core_KE_n3295) );
  OAI2BB2X1 U24666 ( .B0(n1420), .B1(n1937), .A0N(top_core_KE_key_mem_5__79_), 
        .A1N(n1948), .Y(top_core_KE_n3424) );
  OAI2BB2X1 U24667 ( .B0(n1420), .B1(n1957), .A0N(top_core_KE_key_mem_6__79_), 
        .A1N(n1968), .Y(top_core_KE_n3553) );
  OAI2BB2X1 U24668 ( .B0(n1420), .B1(n1985), .A0N(top_core_KE_key_mem_7__79_), 
        .A1N(n1988), .Y(top_core_KE_n3682) );
  OAI2BB2X1 U24669 ( .B0(n1420), .B1(n2037), .A0N(top_core_KE_key_mem_10__79_), 
        .A1N(n2044), .Y(top_core_KE_n4069) );
  OAI2BB2X1 U24670 ( .B0(n1420), .B1(n2065), .A0N(top_core_KE_key_mem_11__79_), 
        .A1N(n2068), .Y(top_core_KE_n4198) );
  OAI2BB2X1 U24671 ( .B0(n1420), .B1(n2077), .A0N(top_core_KE_key_mem_12__79_), 
        .A1N(n2088), .Y(top_core_KE_n4327) );
  OAI2BB2X1 U24672 ( .B0(n1420), .B1(n2105), .A0N(top_core_KE_key_mem_13__79_), 
        .A1N(n2108), .Y(top_core_KE_n4456) );
  OAI2BB2X1 U24673 ( .B0(n1420), .B1(n2125), .A0N(top_core_KE_key_mem_14__79_), 
        .A1N(n2128), .Y(top_core_KE_n4585) );
  OAI2BB2X1 U24674 ( .B0(n1428), .B1(n1860), .A0N(top_core_KE_key_mem_1__71_), 
        .A1N(n1871), .Y(top_core_KE_n2916) );
  OAI2BB2X1 U24675 ( .B0(n1428), .B1(n1878), .A0N(top_core_KE_key_mem_2__71_), 
        .A1N(n1889), .Y(top_core_KE_n3045) );
  OAI2BB2X1 U24676 ( .B0(n1428), .B1(n1898), .A0N(top_core_KE_key_mem_3__71_), 
        .A1N(n1908), .Y(top_core_KE_n3174) );
  OAI2BB2X1 U24677 ( .B0(n1428), .B1(n1918), .A0N(top_core_KE_key_mem_4__71_), 
        .A1N(n1929), .Y(top_core_KE_n3303) );
  OAI2BB2X1 U24678 ( .B0(n1428), .B1(n1939), .A0N(top_core_KE_key_mem_5__71_), 
        .A1N(n1948), .Y(top_core_KE_n3432) );
  OAI2BB2X1 U24679 ( .B0(n1428), .B1(n1958), .A0N(top_core_KE_key_mem_6__71_), 
        .A1N(n1968), .Y(top_core_KE_n3561) );
  OAI2BB2X1 U24680 ( .B0(n1428), .B1(n1977), .A0N(top_core_KE_key_mem_7__71_), 
        .A1N(n1988), .Y(top_core_KE_n3690) );
  OAI2BB2X1 U24681 ( .B0(n1428), .B1(n2038), .A0N(top_core_KE_key_mem_10__71_), 
        .A1N(n2049), .Y(top_core_KE_n4077) );
  OAI2BB2X1 U24682 ( .B0(n1428), .B1(n2057), .A0N(top_core_KE_key_mem_11__71_), 
        .A1N(n2068), .Y(top_core_KE_n4206) );
  OAI2BB2X1 U24683 ( .B0(n1428), .B1(n2079), .A0N(top_core_KE_key_mem_12__71_), 
        .A1N(n2088), .Y(top_core_KE_n4335) );
  OAI2BB2X1 U24684 ( .B0(n1428), .B1(n2097), .A0N(top_core_KE_key_mem_13__71_), 
        .A1N(n2108), .Y(top_core_KE_n4464) );
  OAI2BB2X1 U24685 ( .B0(n1428), .B1(n2117), .A0N(top_core_KE_key_mem_14__71_), 
        .A1N(n2128), .Y(top_core_KE_n4593) );
  OAI2BB2X1 U24686 ( .B0(n1373), .B1(n1865), .A0N(top_core_KE_key_mem_1__126_), 
        .A1N(n1866), .Y(top_core_KE_n2861) );
  OAI2BB2X1 U24687 ( .B0(n1373), .B1(n1879), .A0N(top_core_KE_key_mem_2__126_), 
        .A1N(n1887), .Y(top_core_KE_n2990) );
  OAI2BB2X1 U24688 ( .B0(n1373), .B1(n1898), .A0N(top_core_KE_key_mem_3__126_), 
        .A1N(n1906), .Y(top_core_KE_n3119) );
  OAI2BB2X1 U24689 ( .B0(n1373), .B1(n1919), .A0N(top_core_KE_key_mem_4__126_), 
        .A1N(n1927), .Y(top_core_KE_n3248) );
  OAI2BB2X1 U24690 ( .B0(n1373), .B1(n1938), .A0N(top_core_KE_key_mem_5__126_), 
        .A1N(n1946), .Y(top_core_KE_n3377) );
  OAI2BB2X1 U24691 ( .B0(n1373), .B1(n1959), .A0N(top_core_KE_key_mem_6__126_), 
        .A1N(n1967), .Y(top_core_KE_n3506) );
  OAI2BB2X1 U24692 ( .B0(n1373), .B1(n1978), .A0N(top_core_KE_key_mem_7__126_), 
        .A1N(n1986), .Y(top_core_KE_n3635) );
  OAI2BB2X1 U24693 ( .B0(n1373), .B1(n2039), .A0N(top_core_KE_key_mem_10__126_), .A1N(n2047), .Y(top_core_KE_n4022) );
  OAI2BB2X1 U24694 ( .B0(n1373), .B1(n2058), .A0N(top_core_KE_key_mem_11__126_), .A1N(n2066), .Y(top_core_KE_n4151) );
  OAI2BB2X1 U24695 ( .B0(n1373), .B1(n2078), .A0N(top_core_KE_key_mem_12__126_), .A1N(n2086), .Y(top_core_KE_n4280) );
  OAI2BB2X1 U24696 ( .B0(n1373), .B1(n2098), .A0N(top_core_KE_key_mem_13__126_), .A1N(n2106), .Y(top_core_KE_n4409) );
  OAI2BB2X1 U24697 ( .B0(n1373), .B1(n2118), .A0N(top_core_KE_key_mem_14__126_), .A1N(n2126), .Y(top_core_KE_n4538) );
  OAI2BB2X1 U24698 ( .B0(n1374), .B1(n1861), .A0N(top_core_KE_key_mem_1__125_), 
        .A1N(n1868), .Y(top_core_KE_n2862) );
  OAI2BB2X1 U24699 ( .B0(n1374), .B1(n1885), .A0N(top_core_KE_key_mem_2__125_), 
        .A1N(n1888), .Y(top_core_KE_n2991) );
  OAI2BB2X1 U24700 ( .B0(n1374), .B1(n1904), .A0N(top_core_KE_key_mem_3__125_), 
        .A1N(n1907), .Y(top_core_KE_n3120) );
  OAI2BB2X1 U24701 ( .B0(n1374), .B1(n1925), .A0N(top_core_KE_key_mem_4__125_), 
        .A1N(n1928), .Y(top_core_KE_n3249) );
  OAI2BB2X1 U24702 ( .B0(n1374), .B1(n1944), .A0N(top_core_KE_key_mem_5__125_), 
        .A1N(n1947), .Y(top_core_KE_n3378) );
  OAI2BB2X1 U24703 ( .B0(n1374), .B1(n1965), .A0N(top_core_KE_key_mem_6__125_), 
        .A1N(n1961), .Y(top_core_KE_n3507) );
  OAI2BB2X1 U24704 ( .B0(n1374), .B1(n1984), .A0N(top_core_KE_key_mem_7__125_), 
        .A1N(n1987), .Y(top_core_KE_n3636) );
  OAI2BB2X1 U24705 ( .B0(n1374), .B1(n2045), .A0N(top_core_KE_key_mem_10__125_), .A1N(n2048), .Y(top_core_KE_n4023) );
  OAI2BB2X1 U24706 ( .B0(n1374), .B1(n2064), .A0N(top_core_KE_key_mem_11__125_), .A1N(n2067), .Y(top_core_KE_n4152) );
  OAI2BB2X1 U24707 ( .B0(n1374), .B1(n2084), .A0N(top_core_KE_key_mem_12__125_), .A1N(n2087), .Y(top_core_KE_n4281) );
  OAI2BB2X1 U24708 ( .B0(n1374), .B1(n2104), .A0N(top_core_KE_key_mem_13__125_), .A1N(n2107), .Y(top_core_KE_n4410) );
  OAI2BB2X1 U24709 ( .B0(n1374), .B1(n2124), .A0N(top_core_KE_key_mem_14__125_), .A1N(n2127), .Y(top_core_KE_n4539) );
  OAI2BB2X1 U24710 ( .B0(n1375), .B1(n1858), .A0N(top_core_KE_key_mem_1__124_), 
        .A1N(n1866), .Y(top_core_KE_n2863) );
  OAI2BB2X1 U24711 ( .B0(n1375), .B1(n1885), .A0N(top_core_KE_key_mem_2__124_), 
        .A1N(n1887), .Y(top_core_KE_n2992) );
  OAI2BB2X1 U24712 ( .B0(n1375), .B1(n1904), .A0N(top_core_KE_key_mem_3__124_), 
        .A1N(n1906), .Y(top_core_KE_n3121) );
  OAI2BB2X1 U24713 ( .B0(n1375), .B1(n1925), .A0N(top_core_KE_key_mem_4__124_), 
        .A1N(n1927), .Y(top_core_KE_n3250) );
  OAI2BB2X1 U24714 ( .B0(n1375), .B1(n1944), .A0N(top_core_KE_key_mem_5__124_), 
        .A1N(n1946), .Y(top_core_KE_n3379) );
  OAI2BB2X1 U24715 ( .B0(n1375), .B1(n1965), .A0N(top_core_KE_key_mem_6__124_), 
        .A1N(n1967), .Y(top_core_KE_n3508) );
  OAI2BB2X1 U24716 ( .B0(n1375), .B1(n1984), .A0N(top_core_KE_key_mem_7__124_), 
        .A1N(n1986), .Y(top_core_KE_n3637) );
  OAI2BB2X1 U24717 ( .B0(n1375), .B1(n2045), .A0N(top_core_KE_key_mem_10__124_), .A1N(n2047), .Y(top_core_KE_n4024) );
  OAI2BB2X1 U24718 ( .B0(n1375), .B1(n2064), .A0N(top_core_KE_key_mem_11__124_), .A1N(n2066), .Y(top_core_KE_n4153) );
  OAI2BB2X1 U24719 ( .B0(n1375), .B1(n2084), .A0N(top_core_KE_key_mem_12__124_), .A1N(n2086), .Y(top_core_KE_n4282) );
  OAI2BB2X1 U24720 ( .B0(n1375), .B1(n2104), .A0N(top_core_KE_key_mem_13__124_), .A1N(n2106), .Y(top_core_KE_n4411) );
  OAI2BB2X1 U24721 ( .B0(n1375), .B1(n2124), .A0N(top_core_KE_key_mem_14__124_), .A1N(n2126), .Y(top_core_KE_n4540) );
  OAI2BB2X1 U24722 ( .B0(n1376), .B1(n1867), .A0N(top_core_KE_key_mem_1__123_), 
        .A1N(n1866), .Y(top_core_KE_n2864) );
  OAI2BB2X1 U24723 ( .B0(n1376), .B1(n1877), .A0N(top_core_KE_key_mem_2__123_), 
        .A1N(n1887), .Y(top_core_KE_n2993) );
  OAI2BB2X1 U24724 ( .B0(n1376), .B1(n1897), .A0N(top_core_KE_key_mem_3__123_), 
        .A1N(n1906), .Y(top_core_KE_n3122) );
  OAI2BB2X1 U24725 ( .B0(n1376), .B1(n1917), .A0N(top_core_KE_key_mem_4__123_), 
        .A1N(n1927), .Y(top_core_KE_n3251) );
  OAI2BB2X1 U24726 ( .B0(n1376), .B1(n1937), .A0N(top_core_KE_key_mem_5__123_), 
        .A1N(n1946), .Y(top_core_KE_n3380) );
  OAI2BB2X1 U24727 ( .B0(n1376), .B1(n1957), .A0N(top_core_KE_key_mem_6__123_), 
        .A1N(n1967), .Y(top_core_KE_n3509) );
  OAI2BB2X1 U24728 ( .B0(n1376), .B1(n1990), .A0N(top_core_KE_key_mem_7__123_), 
        .A1N(n1986), .Y(top_core_KE_n3638) );
  OAI2BB2X1 U24729 ( .B0(n1376), .B1(n2037), .A0N(top_core_KE_key_mem_10__123_), .A1N(n2047), .Y(top_core_KE_n4025) );
  OAI2BB2X1 U24730 ( .B0(n1376), .B1(n2070), .A0N(top_core_KE_key_mem_11__123_), .A1N(n2066), .Y(top_core_KE_n4154) );
  OAI2BB2X1 U24731 ( .B0(n1376), .B1(n2077), .A0N(top_core_KE_key_mem_12__123_), .A1N(n2086), .Y(top_core_KE_n4283) );
  OAI2BB2X1 U24732 ( .B0(n1376), .B1(n2110), .A0N(top_core_KE_key_mem_13__123_), .A1N(n2106), .Y(top_core_KE_n4412) );
  OAI2BB2X1 U24733 ( .B0(n1376), .B1(n2130), .A0N(top_core_KE_key_mem_14__123_), .A1N(n2126), .Y(top_core_KE_n4541) );
  OAI2BB2X1 U24734 ( .B0(n1377), .B1(n1872), .A0N(top_core_KE_key_mem_1__122_), 
        .A1N(n1867), .Y(top_core_KE_n2865) );
  OAI2BB2X1 U24735 ( .B0(n1377), .B1(n1884), .A0N(top_core_KE_key_mem_2__122_), 
        .A1N(n1887), .Y(top_core_KE_n2994) );
  OAI2BB2X1 U24736 ( .B0(n1377), .B1(n1903), .A0N(top_core_KE_key_mem_3__122_), 
        .A1N(n1906), .Y(top_core_KE_n3123) );
  OAI2BB2X1 U24737 ( .B0(n1377), .B1(n1924), .A0N(top_core_KE_key_mem_4__122_), 
        .A1N(n1927), .Y(top_core_KE_n3252) );
  OAI2BB2X1 U24738 ( .B0(n1377), .B1(n1943), .A0N(top_core_KE_key_mem_5__122_), 
        .A1N(n1946), .Y(top_core_KE_n3381) );
  OAI2BB2X1 U24739 ( .B0(n1377), .B1(n1964), .A0N(top_core_KE_key_mem_6__122_), 
        .A1N(n1967), .Y(top_core_KE_n3510) );
  OAI2BB2X1 U24740 ( .B0(n1377), .B1(n1983), .A0N(top_core_KE_key_mem_7__122_), 
        .A1N(n1986), .Y(top_core_KE_n3639) );
  OAI2BB2X1 U24741 ( .B0(n1377), .B1(n2044), .A0N(top_core_KE_key_mem_10__122_), .A1N(n2047), .Y(top_core_KE_n4026) );
  OAI2BB2X1 U24742 ( .B0(n1377), .B1(n2063), .A0N(top_core_KE_key_mem_11__122_), .A1N(n2066), .Y(top_core_KE_n4155) );
  OAI2BB2X1 U24743 ( .B0(n1377), .B1(n2083), .A0N(top_core_KE_key_mem_12__122_), .A1N(n2086), .Y(top_core_KE_n4284) );
  OAI2BB2X1 U24744 ( .B0(n1377), .B1(n2103), .A0N(top_core_KE_key_mem_13__122_), .A1N(n2106), .Y(top_core_KE_n4413) );
  OAI2BB2X1 U24745 ( .B0(n1377), .B1(n2123), .A0N(top_core_KE_key_mem_14__122_), .A1N(n2126), .Y(top_core_KE_n4542) );
  OAI2BB2X1 U24746 ( .B0(n1378), .B1(n1871), .A0N(top_core_KE_key_mem_1__121_), 
        .A1N(n1866), .Y(top_core_KE_n2866) );
  OAI2BB2X1 U24747 ( .B0(n1378), .B1(n1882), .A0N(top_core_KE_key_mem_2__121_), 
        .A1N(n1887), .Y(top_core_KE_n2995) );
  OAI2BB2X1 U24748 ( .B0(n1378), .B1(n1901), .A0N(top_core_KE_key_mem_3__121_), 
        .A1N(n1906), .Y(top_core_KE_n3124) );
  OAI2BB2X1 U24749 ( .B0(n1378), .B1(n1922), .A0N(top_core_KE_key_mem_4__121_), 
        .A1N(n1927), .Y(top_core_KE_n3253) );
  OAI2BB2X1 U24750 ( .B0(n1378), .B1(n1941), .A0N(top_core_KE_key_mem_5__121_), 
        .A1N(n1946), .Y(top_core_KE_n3382) );
  OAI2BB2X1 U24751 ( .B0(n1378), .B1(n1962), .A0N(top_core_KE_key_mem_6__121_), 
        .A1N(n1967), .Y(top_core_KE_n3511) );
  OAI2BB2X1 U24752 ( .B0(n1378), .B1(n1981), .A0N(top_core_KE_key_mem_7__121_), 
        .A1N(n1986), .Y(top_core_KE_n3640) );
  OAI2BB2X1 U24753 ( .B0(n1378), .B1(n2042), .A0N(top_core_KE_key_mem_10__121_), .A1N(n2047), .Y(top_core_KE_n4027) );
  OAI2BB2X1 U24754 ( .B0(n1378), .B1(n2061), .A0N(top_core_KE_key_mem_11__121_), .A1N(n2066), .Y(top_core_KE_n4156) );
  OAI2BB2X1 U24755 ( .B0(n1378), .B1(n2081), .A0N(top_core_KE_key_mem_12__121_), .A1N(n2086), .Y(top_core_KE_n4285) );
  OAI2BB2X1 U24756 ( .B0(n1378), .B1(n2101), .A0N(top_core_KE_key_mem_13__121_), .A1N(n2106), .Y(top_core_KE_n4414) );
  OAI2BB2X1 U24757 ( .B0(n1378), .B1(n2121), .A0N(top_core_KE_key_mem_14__121_), .A1N(n2126), .Y(top_core_KE_n4543) );
  OAI2BB2X1 U24758 ( .B0(n1379), .B1(n1868), .A0N(top_core_KE_key_mem_1__120_), 
        .A1N(n1866), .Y(top_core_KE_n2867) );
  OAI2BB2X1 U24759 ( .B0(n1379), .B1(n1884), .A0N(top_core_KE_key_mem_2__120_), 
        .A1N(n1886), .Y(top_core_KE_n2996) );
  OAI2BB2X1 U24760 ( .B0(n1379), .B1(n1903), .A0N(top_core_KE_key_mem_3__120_), 
        .A1N(n1905), .Y(top_core_KE_n3125) );
  OAI2BB2X1 U24761 ( .B0(n1379), .B1(n1924), .A0N(top_core_KE_key_mem_4__120_), 
        .A1N(n1926), .Y(top_core_KE_n3254) );
  OAI2BB2X1 U24762 ( .B0(n1379), .B1(n1943), .A0N(top_core_KE_key_mem_5__120_), 
        .A1N(n1945), .Y(top_core_KE_n3383) );
  OAI2BB2X1 U24763 ( .B0(n1379), .B1(n1964), .A0N(top_core_KE_key_mem_6__120_), 
        .A1N(n1966), .Y(top_core_KE_n3512) );
  OAI2BB2X1 U24764 ( .B0(n1379), .B1(n1983), .A0N(top_core_KE_key_mem_7__120_), 
        .A1N(n1985), .Y(top_core_KE_n3641) );
  OAI2BB2X1 U24765 ( .B0(n1379), .B1(n2044), .A0N(top_core_KE_key_mem_10__120_), .A1N(n2046), .Y(top_core_KE_n4028) );
  OAI2BB2X1 U24766 ( .B0(n1379), .B1(n2063), .A0N(top_core_KE_key_mem_11__120_), .A1N(n2065), .Y(top_core_KE_n4157) );
  OAI2BB2X1 U24767 ( .B0(n1379), .B1(n2083), .A0N(top_core_KE_key_mem_12__120_), .A1N(n2085), .Y(top_core_KE_n4286) );
  OAI2BB2X1 U24768 ( .B0(n1379), .B1(n2103), .A0N(top_core_KE_key_mem_13__120_), .A1N(n2105), .Y(top_core_KE_n4415) );
  OAI2BB2X1 U24769 ( .B0(n1379), .B1(n2123), .A0N(top_core_KE_key_mem_14__120_), .A1N(n2125), .Y(top_core_KE_n4544) );
  OAI2BB2X1 U24770 ( .B0(n1388), .B1(n1857), .A0N(top_core_KE_key_mem_1__111_), 
        .A1N(n1867), .Y(top_core_KE_n2876) );
  OAI2BB2X1 U24771 ( .B0(n1388), .B1(n1882), .A0N(top_core_KE_key_mem_2__111_), 
        .A1N(n1885), .Y(top_core_KE_n3005) );
  OAI2BB2X1 U24772 ( .B0(n1388), .B1(n1901), .A0N(top_core_KE_key_mem_3__111_), 
        .A1N(n1904), .Y(top_core_KE_n3134) );
  OAI2BB2X1 U24773 ( .B0(n1388), .B1(n1922), .A0N(top_core_KE_key_mem_4__111_), 
        .A1N(n1925), .Y(top_core_KE_n3263) );
  OAI2BB2X1 U24774 ( .B0(n1388), .B1(n1941), .A0N(top_core_KE_key_mem_5__111_), 
        .A1N(n1944), .Y(top_core_KE_n3392) );
  OAI2BB2X1 U24775 ( .B0(n1388), .B1(n1962), .A0N(top_core_KE_key_mem_6__111_), 
        .A1N(n1965), .Y(top_core_KE_n3521) );
  OAI2BB2X1 U24776 ( .B0(n1388), .B1(n1981), .A0N(top_core_KE_key_mem_7__111_), 
        .A1N(n1984), .Y(top_core_KE_n3650) );
  OAI2BB2X1 U24777 ( .B0(n1388), .B1(n2042), .A0N(top_core_KE_key_mem_10__111_), .A1N(n2045), .Y(top_core_KE_n4037) );
  OAI2BB2X1 U24778 ( .B0(n1388), .B1(n2061), .A0N(top_core_KE_key_mem_11__111_), .A1N(n2064), .Y(top_core_KE_n4166) );
  OAI2BB2X1 U24779 ( .B0(n1388), .B1(n2081), .A0N(top_core_KE_key_mem_12__111_), .A1N(n2084), .Y(top_core_KE_n4295) );
  OAI2BB2X1 U24780 ( .B0(n1388), .B1(n2101), .A0N(top_core_KE_key_mem_13__111_), .A1N(n2104), .Y(top_core_KE_n4424) );
  OAI2BB2X1 U24781 ( .B0(n1388), .B1(n2121), .A0N(top_core_KE_key_mem_14__111_), .A1N(n2124), .Y(top_core_KE_n4553) );
  OAI2BB2X1 U24782 ( .B0(n1389), .B1(n1857), .A0N(top_core_KE_key_mem_1__110_), 
        .A1N(n1868), .Y(top_core_KE_n2877) );
  OAI2BB2X1 U24783 ( .B0(n1389), .B1(n1882), .A0N(top_core_KE_key_mem_2__110_), 
        .A1N(n1885), .Y(top_core_KE_n3006) );
  OAI2BB2X1 U24784 ( .B0(n1389), .B1(n1901), .A0N(top_core_KE_key_mem_3__110_), 
        .A1N(n1904), .Y(top_core_KE_n3135) );
  OAI2BB2X1 U24785 ( .B0(n1389), .B1(n1922), .A0N(top_core_KE_key_mem_4__110_), 
        .A1N(n1925), .Y(top_core_KE_n3264) );
  OAI2BB2X1 U24786 ( .B0(n1389), .B1(n1941), .A0N(top_core_KE_key_mem_5__110_), 
        .A1N(n1944), .Y(top_core_KE_n3393) );
  OAI2BB2X1 U24787 ( .B0(n1389), .B1(n1962), .A0N(top_core_KE_key_mem_6__110_), 
        .A1N(n1965), .Y(top_core_KE_n3522) );
  OAI2BB2X1 U24788 ( .B0(n1389), .B1(n1981), .A0N(top_core_KE_key_mem_7__110_), 
        .A1N(n1984), .Y(top_core_KE_n3651) );
  OAI2BB2X1 U24789 ( .B0(n1389), .B1(n2042), .A0N(top_core_KE_key_mem_10__110_), .A1N(n2045), .Y(top_core_KE_n4038) );
  OAI2BB2X1 U24790 ( .B0(n1389), .B1(n2061), .A0N(top_core_KE_key_mem_11__110_), .A1N(n2064), .Y(top_core_KE_n4167) );
  OAI2BB2X1 U24791 ( .B0(n1389), .B1(n2081), .A0N(top_core_KE_key_mem_12__110_), .A1N(n2084), .Y(top_core_KE_n4296) );
  OAI2BB2X1 U24792 ( .B0(n1389), .B1(n2101), .A0N(top_core_KE_key_mem_13__110_), .A1N(n2104), .Y(top_core_KE_n4425) );
  OAI2BB2X1 U24793 ( .B0(n1389), .B1(n2121), .A0N(top_core_KE_key_mem_14__110_), .A1N(n2124), .Y(top_core_KE_n4554) );
  OAI2BB2X1 U24794 ( .B0(n1390), .B1(n1857), .A0N(top_core_KE_key_mem_1__109_), 
        .A1N(n1868), .Y(top_core_KE_n2878) );
  OAI2BB2X1 U24795 ( .B0(n1390), .B1(n1881), .A0N(top_core_KE_key_mem_2__109_), 
        .A1N(n1885), .Y(top_core_KE_n3007) );
  OAI2BB2X1 U24796 ( .B0(n1390), .B1(n1900), .A0N(top_core_KE_key_mem_3__109_), 
        .A1N(n1904), .Y(top_core_KE_n3136) );
  OAI2BB2X1 U24797 ( .B0(n1390), .B1(n1921), .A0N(top_core_KE_key_mem_4__109_), 
        .A1N(n1925), .Y(top_core_KE_n3265) );
  OAI2BB2X1 U24798 ( .B0(n1390), .B1(n1940), .A0N(top_core_KE_key_mem_5__109_), 
        .A1N(n1944), .Y(top_core_KE_n3394) );
  OAI2BB2X1 U24799 ( .B0(n1390), .B1(n1961), .A0N(top_core_KE_key_mem_6__109_), 
        .A1N(n1965), .Y(top_core_KE_n3523) );
  OAI2BB2X1 U24800 ( .B0(n1390), .B1(n1980), .A0N(top_core_KE_key_mem_7__109_), 
        .A1N(n1984), .Y(top_core_KE_n3652) );
  OAI2BB2X1 U24801 ( .B0(n1390), .B1(n2041), .A0N(top_core_KE_key_mem_10__109_), .A1N(n2045), .Y(top_core_KE_n4039) );
  OAI2BB2X1 U24802 ( .B0(n1390), .B1(n2060), .A0N(top_core_KE_key_mem_11__109_), .A1N(n2064), .Y(top_core_KE_n4168) );
  OAI2BB2X1 U24803 ( .B0(n1390), .B1(n2080), .A0N(top_core_KE_key_mem_12__109_), .A1N(n2084), .Y(top_core_KE_n4297) );
  OAI2BB2X1 U24804 ( .B0(n1390), .B1(n2100), .A0N(top_core_KE_key_mem_13__109_), .A1N(n2104), .Y(top_core_KE_n4426) );
  OAI2BB2X1 U24805 ( .B0(n1390), .B1(n2120), .A0N(top_core_KE_key_mem_14__109_), .A1N(n2124), .Y(top_core_KE_n4555) );
  OAI2BB2X1 U24806 ( .B0(n1391), .B1(n1857), .A0N(top_core_KE_key_mem_1__108_), 
        .A1N(n1867), .Y(top_core_KE_n2879) );
  OAI2BB2X1 U24807 ( .B0(n1391), .B1(n1881), .A0N(top_core_KE_key_mem_2__108_), 
        .A1N(n1886), .Y(top_core_KE_n3008) );
  OAI2BB2X1 U24808 ( .B0(n1391), .B1(n1900), .A0N(top_core_KE_key_mem_3__108_), 
        .A1N(n1905), .Y(top_core_KE_n3137) );
  OAI2BB2X1 U24809 ( .B0(n1391), .B1(n1921), .A0N(top_core_KE_key_mem_4__108_), 
        .A1N(n1926), .Y(top_core_KE_n3266) );
  OAI2BB2X1 U24810 ( .B0(n1391), .B1(n1940), .A0N(top_core_KE_key_mem_5__108_), 
        .A1N(n1945), .Y(top_core_KE_n3395) );
  OAI2BB2X1 U24811 ( .B0(n1391), .B1(n1961), .A0N(top_core_KE_key_mem_6__108_), 
        .A1N(n1966), .Y(top_core_KE_n3524) );
  OAI2BB2X1 U24812 ( .B0(n1391), .B1(n1980), .A0N(top_core_KE_key_mem_7__108_), 
        .A1N(n1985), .Y(top_core_KE_n3653) );
  OAI2BB2X1 U24813 ( .B0(n1391), .B1(n2041), .A0N(top_core_KE_key_mem_10__108_), .A1N(n2046), .Y(top_core_KE_n4040) );
  OAI2BB2X1 U24814 ( .B0(n1391), .B1(n2060), .A0N(top_core_KE_key_mem_11__108_), .A1N(n2065), .Y(top_core_KE_n4169) );
  OAI2BB2X1 U24815 ( .B0(n1391), .B1(n2080), .A0N(top_core_KE_key_mem_12__108_), .A1N(n2085), .Y(top_core_KE_n4298) );
  OAI2BB2X1 U24816 ( .B0(n1391), .B1(n2100), .A0N(top_core_KE_key_mem_13__108_), .A1N(n2105), .Y(top_core_KE_n4427) );
  OAI2BB2X1 U24817 ( .B0(n1391), .B1(n2120), .A0N(top_core_KE_key_mem_14__108_), .A1N(n2125), .Y(top_core_KE_n4556) );
  OAI2BB2X1 U24818 ( .B0(n1392), .B1(n1857), .A0N(top_core_KE_key_mem_1__107_), 
        .A1N(n1868), .Y(top_core_KE_n2880) );
  OAI2BB2X1 U24819 ( .B0(n1392), .B1(n1881), .A0N(top_core_KE_key_mem_2__107_), 
        .A1N(n1886), .Y(top_core_KE_n3009) );
  OAI2BB2X1 U24820 ( .B0(n1392), .B1(n1900), .A0N(top_core_KE_key_mem_3__107_), 
        .A1N(n1905), .Y(top_core_KE_n3138) );
  OAI2BB2X1 U24821 ( .B0(n1392), .B1(n1921), .A0N(top_core_KE_key_mem_4__107_), 
        .A1N(n1926), .Y(top_core_KE_n3267) );
  OAI2BB2X1 U24822 ( .B0(n1392), .B1(n1940), .A0N(top_core_KE_key_mem_5__107_), 
        .A1N(n1945), .Y(top_core_KE_n3396) );
  OAI2BB2X1 U24823 ( .B0(n1392), .B1(n1961), .A0N(top_core_KE_key_mem_6__107_), 
        .A1N(n1966), .Y(top_core_KE_n3525) );
  OAI2BB2X1 U24824 ( .B0(n1392), .B1(n1980), .A0N(top_core_KE_key_mem_7__107_), 
        .A1N(n1985), .Y(top_core_KE_n3654) );
  OAI2BB2X1 U24825 ( .B0(n1392), .B1(n2041), .A0N(top_core_KE_key_mem_10__107_), .A1N(n2046), .Y(top_core_KE_n4041) );
  OAI2BB2X1 U24826 ( .B0(n1392), .B1(n2060), .A0N(top_core_KE_key_mem_11__107_), .A1N(n2065), .Y(top_core_KE_n4170) );
  OAI2BB2X1 U24827 ( .B0(n1392), .B1(n2080), .A0N(top_core_KE_key_mem_12__107_), .A1N(n2085), .Y(top_core_KE_n4299) );
  OAI2BB2X1 U24828 ( .B0(n1392), .B1(n2100), .A0N(top_core_KE_key_mem_13__107_), .A1N(n2105), .Y(top_core_KE_n4428) );
  OAI2BB2X1 U24829 ( .B0(n1392), .B1(n2120), .A0N(top_core_KE_key_mem_14__107_), .A1N(n2125), .Y(top_core_KE_n4557) );
  OAI2BB2X1 U24830 ( .B0(n1393), .B1(n1857), .A0N(top_core_KE_key_mem_1__106_), 
        .A1N(n1868), .Y(top_core_KE_n2881) );
  OAI2BB2X1 U24831 ( .B0(n1393), .B1(n1881), .A0N(top_core_KE_key_mem_2__106_), 
        .A1N(n1886), .Y(top_core_KE_n3010) );
  OAI2BB2X1 U24832 ( .B0(n1393), .B1(n1900), .A0N(top_core_KE_key_mem_3__106_), 
        .A1N(n1905), .Y(top_core_KE_n3139) );
  OAI2BB2X1 U24833 ( .B0(n1393), .B1(n1921), .A0N(top_core_KE_key_mem_4__106_), 
        .A1N(n1926), .Y(top_core_KE_n3268) );
  OAI2BB2X1 U24834 ( .B0(n1393), .B1(n1940), .A0N(top_core_KE_key_mem_5__106_), 
        .A1N(n1945), .Y(top_core_KE_n3397) );
  OAI2BB2X1 U24835 ( .B0(n1393), .B1(n1961), .A0N(top_core_KE_key_mem_6__106_), 
        .A1N(n1966), .Y(top_core_KE_n3526) );
  OAI2BB2X1 U24836 ( .B0(n1393), .B1(n1980), .A0N(top_core_KE_key_mem_7__106_), 
        .A1N(n1985), .Y(top_core_KE_n3655) );
  OAI2BB2X1 U24837 ( .B0(n1393), .B1(n2041), .A0N(top_core_KE_key_mem_10__106_), .A1N(n2046), .Y(top_core_KE_n4042) );
  OAI2BB2X1 U24838 ( .B0(n1393), .B1(n2060), .A0N(top_core_KE_key_mem_11__106_), .A1N(n2065), .Y(top_core_KE_n4171) );
  OAI2BB2X1 U24839 ( .B0(n1393), .B1(n2080), .A0N(top_core_KE_key_mem_12__106_), .A1N(n2085), .Y(top_core_KE_n4300) );
  OAI2BB2X1 U24840 ( .B0(n1393), .B1(n2100), .A0N(top_core_KE_key_mem_13__106_), .A1N(n2105), .Y(top_core_KE_n4429) );
  OAI2BB2X1 U24841 ( .B0(n1393), .B1(n2120), .A0N(top_core_KE_key_mem_14__106_), .A1N(n2125), .Y(top_core_KE_n4558) );
  OAI2BB2X1 U24842 ( .B0(n1394), .B1(n1857), .A0N(top_core_KE_key_mem_1__105_), 
        .A1N(n1868), .Y(top_core_KE_n2882) );
  OAI2BB2X1 U24843 ( .B0(n1394), .B1(n1880), .A0N(top_core_KE_key_mem_2__105_), 
        .A1N(n1886), .Y(top_core_KE_n3011) );
  OAI2BB2X1 U24844 ( .B0(n1394), .B1(n1899), .A0N(top_core_KE_key_mem_3__105_), 
        .A1N(n1905), .Y(top_core_KE_n3140) );
  OAI2BB2X1 U24845 ( .B0(n1394), .B1(n1920), .A0N(top_core_KE_key_mem_4__105_), 
        .A1N(n1926), .Y(top_core_KE_n3269) );
  OAI2BB2X1 U24846 ( .B0(n1394), .B1(n1939), .A0N(top_core_KE_key_mem_5__105_), 
        .A1N(n1945), .Y(top_core_KE_n3398) );
  OAI2BB2X1 U24847 ( .B0(n1394), .B1(n1960), .A0N(top_core_KE_key_mem_6__105_), 
        .A1N(n1966), .Y(top_core_KE_n3527) );
  OAI2BB2X1 U24848 ( .B0(n1394), .B1(n1979), .A0N(top_core_KE_key_mem_7__105_), 
        .A1N(n1985), .Y(top_core_KE_n3656) );
  OAI2BB2X1 U24849 ( .B0(n1394), .B1(n2040), .A0N(top_core_KE_key_mem_10__105_), .A1N(n2046), .Y(top_core_KE_n4043) );
  OAI2BB2X1 U24850 ( .B0(n1394), .B1(n2059), .A0N(top_core_KE_key_mem_11__105_), .A1N(n2065), .Y(top_core_KE_n4172) );
  OAI2BB2X1 U24851 ( .B0(n1394), .B1(n2079), .A0N(top_core_KE_key_mem_12__105_), .A1N(n2085), .Y(top_core_KE_n4301) );
  OAI2BB2X1 U24852 ( .B0(n1394), .B1(n2099), .A0N(top_core_KE_key_mem_13__105_), .A1N(n2105), .Y(top_core_KE_n4430) );
  OAI2BB2X1 U24853 ( .B0(n1394), .B1(n2119), .A0N(top_core_KE_key_mem_14__105_), .A1N(n2125), .Y(top_core_KE_n4559) );
  OAI2BB2X1 U24854 ( .B0(n1395), .B1(n1857), .A0N(top_core_KE_key_mem_1__104_), 
        .A1N(n1868), .Y(top_core_KE_n2883) );
  OAI2BB2X1 U24855 ( .B0(n1395), .B1(n1880), .A0N(top_core_KE_key_mem_2__104_), 
        .A1N(n1886), .Y(top_core_KE_n3012) );
  OAI2BB2X1 U24856 ( .B0(n1395), .B1(n1899), .A0N(top_core_KE_key_mem_3__104_), 
        .A1N(n1905), .Y(top_core_KE_n3141) );
  OAI2BB2X1 U24857 ( .B0(n1395), .B1(n1920), .A0N(top_core_KE_key_mem_4__104_), 
        .A1N(n1926), .Y(top_core_KE_n3270) );
  OAI2BB2X1 U24858 ( .B0(n1395), .B1(n1939), .A0N(top_core_KE_key_mem_5__104_), 
        .A1N(n1945), .Y(top_core_KE_n3399) );
  OAI2BB2X1 U24859 ( .B0(n1395), .B1(n1960), .A0N(top_core_KE_key_mem_6__104_), 
        .A1N(n1966), .Y(top_core_KE_n3528) );
  OAI2BB2X1 U24860 ( .B0(n1395), .B1(n1979), .A0N(top_core_KE_key_mem_7__104_), 
        .A1N(n1985), .Y(top_core_KE_n3657) );
  OAI2BB2X1 U24861 ( .B0(n1395), .B1(n2040), .A0N(top_core_KE_key_mem_10__104_), .A1N(n2046), .Y(top_core_KE_n4044) );
  OAI2BB2X1 U24862 ( .B0(n1395), .B1(n2059), .A0N(top_core_KE_key_mem_11__104_), .A1N(n2065), .Y(top_core_KE_n4173) );
  OAI2BB2X1 U24863 ( .B0(n1395), .B1(n2079), .A0N(top_core_KE_key_mem_12__104_), .A1N(n2085), .Y(top_core_KE_n4302) );
  OAI2BB2X1 U24864 ( .B0(n1395), .B1(n2099), .A0N(top_core_KE_key_mem_13__104_), .A1N(n2105), .Y(top_core_KE_n4431) );
  OAI2BB2X1 U24865 ( .B0(n1395), .B1(n2119), .A0N(top_core_KE_key_mem_14__104_), .A1N(n2125), .Y(top_core_KE_n4560) );
  OAI2BB2X1 U24866 ( .B0(n1396), .B1(n1857), .A0N(top_core_KE_key_mem_1__103_), 
        .A1N(n1868), .Y(top_core_KE_n2884) );
  OAI2BB2X1 U24867 ( .B0(n1396), .B1(n1880), .A0N(top_core_KE_key_mem_2__103_), 
        .A1N(n1886), .Y(top_core_KE_n3013) );
  OAI2BB2X1 U24868 ( .B0(n1396), .B1(n1899), .A0N(top_core_KE_key_mem_3__103_), 
        .A1N(n1905), .Y(top_core_KE_n3142) );
  OAI2BB2X1 U24869 ( .B0(n1396), .B1(n1920), .A0N(top_core_KE_key_mem_4__103_), 
        .A1N(n1926), .Y(top_core_KE_n3271) );
  OAI2BB2X1 U24870 ( .B0(n1396), .B1(n1939), .A0N(top_core_KE_key_mem_5__103_), 
        .A1N(n1945), .Y(top_core_KE_n3400) );
  OAI2BB2X1 U24871 ( .B0(n1396), .B1(n1960), .A0N(top_core_KE_key_mem_6__103_), 
        .A1N(n1966), .Y(top_core_KE_n3529) );
  OAI2BB2X1 U24872 ( .B0(n1396), .B1(n1979), .A0N(top_core_KE_key_mem_7__103_), 
        .A1N(n1985), .Y(top_core_KE_n3658) );
  OAI2BB2X1 U24873 ( .B0(n1396), .B1(n2040), .A0N(top_core_KE_key_mem_10__103_), .A1N(n2046), .Y(top_core_KE_n4045) );
  OAI2BB2X1 U24874 ( .B0(n1396), .B1(n2059), .A0N(top_core_KE_key_mem_11__103_), .A1N(n2065), .Y(top_core_KE_n4174) );
  OAI2BB2X1 U24875 ( .B0(n1396), .B1(n2079), .A0N(top_core_KE_key_mem_12__103_), .A1N(n2085), .Y(top_core_KE_n4303) );
  OAI2BB2X1 U24876 ( .B0(n1396), .B1(n2099), .A0N(top_core_KE_key_mem_13__103_), .A1N(n2105), .Y(top_core_KE_n4432) );
  OAI2BB2X1 U24877 ( .B0(n1396), .B1(n2119), .A0N(top_core_KE_key_mem_14__103_), .A1N(n2125), .Y(top_core_KE_n4561) );
  OAI2BB2X1 U24878 ( .B0(n1397), .B1(n1858), .A0N(top_core_KE_key_mem_1__102_), 
        .A1N(n1868), .Y(top_core_KE_n2885) );
  OAI2BB2X1 U24879 ( .B0(n1397), .B1(n1880), .A0N(top_core_KE_key_mem_2__102_), 
        .A1N(n1888), .Y(top_core_KE_n3014) );
  OAI2BB2X1 U24880 ( .B0(n1397), .B1(n1899), .A0N(top_core_KE_key_mem_3__102_), 
        .A1N(n1907), .Y(top_core_KE_n3143) );
  OAI2BB2X1 U24881 ( .B0(n1397), .B1(n1920), .A0N(top_core_KE_key_mem_4__102_), 
        .A1N(n1928), .Y(top_core_KE_n3272) );
  OAI2BB2X1 U24882 ( .B0(n1397), .B1(n1939), .A0N(top_core_KE_key_mem_5__102_), 
        .A1N(n1947), .Y(top_core_KE_n3401) );
  OAI2BB2X1 U24883 ( .B0(n1397), .B1(n1960), .A0N(top_core_KE_key_mem_6__102_), 
        .A1N(n1958), .Y(top_core_KE_n3530) );
  OAI2BB2X1 U24884 ( .B0(n1397), .B1(n1979), .A0N(top_core_KE_key_mem_7__102_), 
        .A1N(n1987), .Y(top_core_KE_n3659) );
  OAI2BB2X1 U24885 ( .B0(n1397), .B1(n2040), .A0N(top_core_KE_key_mem_10__102_), .A1N(n2048), .Y(top_core_KE_n4046) );
  OAI2BB2X1 U24886 ( .B0(n1397), .B1(n2059), .A0N(top_core_KE_key_mem_11__102_), .A1N(n2067), .Y(top_core_KE_n4175) );
  OAI2BB2X1 U24887 ( .B0(n1397), .B1(n2079), .A0N(top_core_KE_key_mem_12__102_), .A1N(n2087), .Y(top_core_KE_n4304) );
  OAI2BB2X1 U24888 ( .B0(n1397), .B1(n2099), .A0N(top_core_KE_key_mem_13__102_), .A1N(n2107), .Y(top_core_KE_n4433) );
  OAI2BB2X1 U24889 ( .B0(n1397), .B1(n2119), .A0N(top_core_KE_key_mem_14__102_), .A1N(n2127), .Y(top_core_KE_n4562) );
  OAI2BB2X1 U24890 ( .B0(n1398), .B1(n1858), .A0N(top_core_KE_key_mem_1__101_), 
        .A1N(n1868), .Y(top_core_KE_n2886) );
  OAI2BB2X1 U24891 ( .B0(n1398), .B1(top_core_KE_n874), .A0N(
        top_core_KE_key_mem_2__101_), .A1N(n1886), .Y(top_core_KE_n3015) );
  OAI2BB2X1 U24892 ( .B0(n1398), .B1(top_core_KE_n876), .A0N(
        top_core_KE_key_mem_3__101_), .A1N(n1905), .Y(top_core_KE_n3144) );
  OAI2BB2X1 U24893 ( .B0(n1398), .B1(top_core_KE_n877), .A0N(
        top_core_KE_key_mem_4__101_), .A1N(n1926), .Y(top_core_KE_n3273) );
  OAI2BB2X1 U24894 ( .B0(n1398), .B1(top_core_KE_n879), .A0N(
        top_core_KE_key_mem_5__101_), .A1N(n1945), .Y(top_core_KE_n3402) );
  OAI2BB2X1 U24895 ( .B0(n1398), .B1(top_core_KE_n880), .A0N(
        top_core_KE_key_mem_6__101_), .A1N(n1966), .Y(top_core_KE_n3531) );
  OAI2BB2X1 U24896 ( .B0(n1398), .B1(top_core_KE_n881), .A0N(
        top_core_KE_key_mem_7__101_), .A1N(n1985), .Y(top_core_KE_n3660) );
  OAI2BB2X1 U24897 ( .B0(n1398), .B1(top_core_KE_n886), .A0N(
        top_core_KE_key_mem_10__101_), .A1N(n2046), .Y(top_core_KE_n4047) );
  OAI2BB2X1 U24898 ( .B0(n1398), .B1(top_core_KE_n888), .A0N(
        top_core_KE_key_mem_11__101_), .A1N(n2065), .Y(top_core_KE_n4176) );
  OAI2BB2X1 U24899 ( .B0(n1398), .B1(top_core_KE_n889), .A0N(
        top_core_KE_key_mem_12__101_), .A1N(n2085), .Y(top_core_KE_n4305) );
  OAI2BB2X1 U24900 ( .B0(n1398), .B1(top_core_KE_n890), .A0N(
        top_core_KE_key_mem_13__101_), .A1N(n2105), .Y(top_core_KE_n4434) );
  OAI2BB2X1 U24901 ( .B0(n1398), .B1(top_core_KE_n891), .A0N(
        top_core_KE_key_mem_14__101_), .A1N(n2125), .Y(top_core_KE_n4563) );
  OAI2BB2X1 U24902 ( .B0(n1399), .B1(n1858), .A0N(top_core_KE_key_mem_1__100_), 
        .A1N(n1868), .Y(top_core_KE_n2887) );
  OAI2BB2X1 U24903 ( .B0(n1399), .B1(top_core_KE_n874), .A0N(
        top_core_KE_key_mem_2__100_), .A1N(n1886), .Y(top_core_KE_n3016) );
  OAI2BB2X1 U24904 ( .B0(n1399), .B1(top_core_KE_n876), .A0N(
        top_core_KE_key_mem_3__100_), .A1N(n1905), .Y(top_core_KE_n3145) );
  OAI2BB2X1 U24905 ( .B0(n1399), .B1(top_core_KE_n877), .A0N(
        top_core_KE_key_mem_4__100_), .A1N(n1926), .Y(top_core_KE_n3274) );
  OAI2BB2X1 U24906 ( .B0(n1399), .B1(top_core_KE_n879), .A0N(
        top_core_KE_key_mem_5__100_), .A1N(n1945), .Y(top_core_KE_n3403) );
  OAI2BB2X1 U24907 ( .B0(n1399), .B1(top_core_KE_n880), .A0N(
        top_core_KE_key_mem_6__100_), .A1N(n1966), .Y(top_core_KE_n3532) );
  OAI2BB2X1 U24908 ( .B0(n1399), .B1(top_core_KE_n881), .A0N(
        top_core_KE_key_mem_7__100_), .A1N(n1985), .Y(top_core_KE_n3661) );
  OAI2BB2X1 U24909 ( .B0(n1399), .B1(top_core_KE_n886), .A0N(
        top_core_KE_key_mem_10__100_), .A1N(n2046), .Y(top_core_KE_n4048) );
  OAI2BB2X1 U24910 ( .B0(n1399), .B1(top_core_KE_n888), .A0N(
        top_core_KE_key_mem_11__100_), .A1N(n2065), .Y(top_core_KE_n4177) );
  OAI2BB2X1 U24911 ( .B0(n1399), .B1(top_core_KE_n889), .A0N(
        top_core_KE_key_mem_12__100_), .A1N(n2085), .Y(top_core_KE_n4306) );
  OAI2BB2X1 U24912 ( .B0(n1399), .B1(top_core_KE_n890), .A0N(
        top_core_KE_key_mem_13__100_), .A1N(n2105), .Y(top_core_KE_n4435) );
  OAI2BB2X1 U24913 ( .B0(n1399), .B1(top_core_KE_n891), .A0N(
        top_core_KE_key_mem_14__100_), .A1N(n2125), .Y(top_core_KE_n4564) );
  OAI2BB2X1 U24914 ( .B0(n1400), .B1(n1858), .A0N(top_core_KE_key_mem_1__99_), 
        .A1N(n1868), .Y(top_core_KE_n2888) );
  OAI2BB2X1 U24915 ( .B0(n1400), .B1(n1877), .A0N(top_core_KE_key_mem_2__99_), 
        .A1N(n1886), .Y(top_core_KE_n3017) );
  OAI2BB2X1 U24916 ( .B0(n1400), .B1(n1897), .A0N(top_core_KE_key_mem_3__99_), 
        .A1N(n1905), .Y(top_core_KE_n3146) );
  OAI2BB2X1 U24917 ( .B0(n1400), .B1(n1917), .A0N(top_core_KE_key_mem_4__99_), 
        .A1N(n1926), .Y(top_core_KE_n3275) );
  OAI2BB2X1 U24918 ( .B0(n1400), .B1(n1937), .A0N(top_core_KE_key_mem_5__99_), 
        .A1N(n1945), .Y(top_core_KE_n3404) );
  OAI2BB2X1 U24919 ( .B0(n1400), .B1(n1957), .A0N(top_core_KE_key_mem_6__99_), 
        .A1N(n1966), .Y(top_core_KE_n3533) );
  OAI2BB2X1 U24920 ( .B0(n1400), .B1(n1988), .A0N(top_core_KE_key_mem_7__99_), 
        .A1N(n1985), .Y(top_core_KE_n3662) );
  OAI2BB2X1 U24921 ( .B0(n1400), .B1(n2037), .A0N(top_core_KE_key_mem_10__99_), 
        .A1N(n2046), .Y(top_core_KE_n4049) );
  OAI2BB2X1 U24922 ( .B0(n1400), .B1(n2068), .A0N(top_core_KE_key_mem_11__99_), 
        .A1N(n2065), .Y(top_core_KE_n4178) );
  OAI2BB2X1 U24923 ( .B0(n1400), .B1(n2077), .A0N(top_core_KE_key_mem_12__99_), 
        .A1N(n2085), .Y(top_core_KE_n4307) );
  OAI2BB2X1 U24924 ( .B0(n1400), .B1(n2108), .A0N(top_core_KE_key_mem_13__99_), 
        .A1N(n2105), .Y(top_core_KE_n4436) );
  OAI2BB2X1 U24925 ( .B0(n1400), .B1(n2128), .A0N(top_core_KE_key_mem_14__99_), 
        .A1N(n2125), .Y(top_core_KE_n4565) );
  OAI2BB2X1 U24926 ( .B0(n1401), .B1(n1858), .A0N(top_core_KE_key_mem_1__98_), 
        .A1N(n1869), .Y(top_core_KE_n2889) );
  OAI2BB2X1 U24927 ( .B0(n1401), .B1(n1884), .A0N(top_core_KE_key_mem_2__98_), 
        .A1N(n1886), .Y(top_core_KE_n3018) );
  OAI2BB2X1 U24928 ( .B0(n1401), .B1(n1903), .A0N(top_core_KE_key_mem_3__98_), 
        .A1N(n1905), .Y(top_core_KE_n3147) );
  OAI2BB2X1 U24929 ( .B0(n1401), .B1(n1924), .A0N(top_core_KE_key_mem_4__98_), 
        .A1N(n1926), .Y(top_core_KE_n3276) );
  OAI2BB2X1 U24930 ( .B0(n1401), .B1(n1943), .A0N(top_core_KE_key_mem_5__98_), 
        .A1N(n1945), .Y(top_core_KE_n3405) );
  OAI2BB2X1 U24931 ( .B0(n1401), .B1(n1964), .A0N(top_core_KE_key_mem_6__98_), 
        .A1N(n1966), .Y(top_core_KE_n3534) );
  OAI2BB2X1 U24932 ( .B0(n1401), .B1(n1983), .A0N(top_core_KE_key_mem_7__98_), 
        .A1N(n1985), .Y(top_core_KE_n3663) );
  OAI2BB2X1 U24933 ( .B0(n1401), .B1(n2044), .A0N(top_core_KE_key_mem_10__98_), 
        .A1N(n2046), .Y(top_core_KE_n4050) );
  OAI2BB2X1 U24934 ( .B0(n1401), .B1(n2063), .A0N(top_core_KE_key_mem_11__98_), 
        .A1N(n2065), .Y(top_core_KE_n4179) );
  OAI2BB2X1 U24935 ( .B0(n1401), .B1(n2083), .A0N(top_core_KE_key_mem_12__98_), 
        .A1N(n2085), .Y(top_core_KE_n4308) );
  OAI2BB2X1 U24936 ( .B0(n1401), .B1(n2103), .A0N(top_core_KE_key_mem_13__98_), 
        .A1N(n2105), .Y(top_core_KE_n4437) );
  OAI2BB2X1 U24937 ( .B0(n1401), .B1(n2123), .A0N(top_core_KE_key_mem_14__98_), 
        .A1N(n2125), .Y(top_core_KE_n4566) );
  OAI2BB2X1 U24938 ( .B0(n1402), .B1(n1858), .A0N(top_core_KE_key_mem_1__97_), 
        .A1N(n1869), .Y(top_core_KE_n2890) );
  OAI2BB2X1 U24939 ( .B0(n1402), .B1(n1879), .A0N(top_core_KE_key_mem_2__97_), 
        .A1N(n1887), .Y(top_core_KE_n3019) );
  OAI2BB2X1 U24940 ( .B0(n1402), .B1(n1899), .A0N(top_core_KE_key_mem_3__97_), 
        .A1N(n1906), .Y(top_core_KE_n3148) );
  OAI2BB2X1 U24941 ( .B0(n1402), .B1(n1919), .A0N(top_core_KE_key_mem_4__97_), 
        .A1N(n1927), .Y(top_core_KE_n3277) );
  OAI2BB2X1 U24942 ( .B0(n1402), .B1(n1938), .A0N(top_core_KE_key_mem_5__97_), 
        .A1N(n1946), .Y(top_core_KE_n3406) );
  OAI2BB2X1 U24943 ( .B0(n1402), .B1(n1959), .A0N(top_core_KE_key_mem_6__97_), 
        .A1N(n1967), .Y(top_core_KE_n3535) );
  OAI2BB2X1 U24944 ( .B0(n1402), .B1(n1978), .A0N(top_core_KE_key_mem_7__97_), 
        .A1N(n1986), .Y(top_core_KE_n3664) );
  OAI2BB2X1 U24945 ( .B0(n1402), .B1(n2039), .A0N(top_core_KE_key_mem_10__97_), 
        .A1N(n2047), .Y(top_core_KE_n4051) );
  OAI2BB2X1 U24946 ( .B0(n1402), .B1(n2058), .A0N(top_core_KE_key_mem_11__97_), 
        .A1N(n2066), .Y(top_core_KE_n4180) );
  OAI2BB2X1 U24947 ( .B0(n1402), .B1(n2078), .A0N(top_core_KE_key_mem_12__97_), 
        .A1N(n2086), .Y(top_core_KE_n4309) );
  OAI2BB2X1 U24948 ( .B0(n1402), .B1(n2098), .A0N(top_core_KE_key_mem_13__97_), 
        .A1N(n2106), .Y(top_core_KE_n4438) );
  OAI2BB2X1 U24949 ( .B0(n1402), .B1(n2118), .A0N(top_core_KE_key_mem_14__97_), 
        .A1N(n2126), .Y(top_core_KE_n4567) );
  OAI2BB2X1 U24950 ( .B0(n1403), .B1(n1858), .A0N(top_core_KE_key_mem_1__96_), 
        .A1N(n1869), .Y(top_core_KE_n2891) );
  OAI2BB2X1 U24951 ( .B0(n1403), .B1(n1879), .A0N(top_core_KE_key_mem_2__96_), 
        .A1N(n1887), .Y(top_core_KE_n3020) );
  OAI2BB2X1 U24952 ( .B0(n1403), .B1(n1897), .A0N(top_core_KE_key_mem_3__96_), 
        .A1N(n1906), .Y(top_core_KE_n3149) );
  OAI2BB2X1 U24953 ( .B0(n1403), .B1(n1919), .A0N(top_core_KE_key_mem_4__96_), 
        .A1N(n1927), .Y(top_core_KE_n3278) );
  OAI2BB2X1 U24954 ( .B0(n1403), .B1(n1938), .A0N(top_core_KE_key_mem_5__96_), 
        .A1N(n1946), .Y(top_core_KE_n3407) );
  OAI2BB2X1 U24955 ( .B0(n1403), .B1(n1959), .A0N(top_core_KE_key_mem_6__96_), 
        .A1N(n1967), .Y(top_core_KE_n3536) );
  OAI2BB2X1 U24956 ( .B0(n1403), .B1(n1978), .A0N(top_core_KE_key_mem_7__96_), 
        .A1N(n1986), .Y(top_core_KE_n3665) );
  OAI2BB2X1 U24957 ( .B0(n1403), .B1(n2039), .A0N(top_core_KE_key_mem_10__96_), 
        .A1N(n2047), .Y(top_core_KE_n4052) );
  OAI2BB2X1 U24958 ( .B0(n1403), .B1(n2058), .A0N(top_core_KE_key_mem_11__96_), 
        .A1N(n2066), .Y(top_core_KE_n4181) );
  OAI2BB2X1 U24959 ( .B0(n1403), .B1(n2078), .A0N(top_core_KE_key_mem_12__96_), 
        .A1N(n2086), .Y(top_core_KE_n4310) );
  OAI2BB2X1 U24960 ( .B0(n1403), .B1(n2098), .A0N(top_core_KE_key_mem_13__96_), 
        .A1N(n2106), .Y(top_core_KE_n4439) );
  OAI2BB2X1 U24961 ( .B0(n1403), .B1(n2118), .A0N(top_core_KE_key_mem_14__96_), 
        .A1N(n2126), .Y(top_core_KE_n4568) );
  OAI2BB2X1 U24962 ( .B0(n1404), .B1(n1858), .A0N(top_core_KE_key_mem_1__95_), 
        .A1N(n1869), .Y(top_core_KE_n2892) );
  OAI2BB2X1 U24963 ( .B0(n1404), .B1(n1879), .A0N(top_core_KE_key_mem_2__95_), 
        .A1N(n1887), .Y(top_core_KE_n3021) );
  OAI2BB2X1 U24964 ( .B0(n1404), .B1(n1903), .A0N(top_core_KE_key_mem_3__95_), 
        .A1N(n1906), .Y(top_core_KE_n3150) );
  OAI2BB2X1 U24965 ( .B0(n1404), .B1(n1919), .A0N(top_core_KE_key_mem_4__95_), 
        .A1N(n1927), .Y(top_core_KE_n3279) );
  OAI2BB2X1 U24966 ( .B0(n1404), .B1(n1938), .A0N(top_core_KE_key_mem_5__95_), 
        .A1N(n1946), .Y(top_core_KE_n3408) );
  OAI2BB2X1 U24967 ( .B0(n1404), .B1(n1959), .A0N(top_core_KE_key_mem_6__95_), 
        .A1N(n1967), .Y(top_core_KE_n3537) );
  OAI2BB2X1 U24968 ( .B0(n1404), .B1(n1978), .A0N(top_core_KE_key_mem_7__95_), 
        .A1N(n1986), .Y(top_core_KE_n3666) );
  OAI2BB2X1 U24969 ( .B0(n1404), .B1(n2039), .A0N(top_core_KE_key_mem_10__95_), 
        .A1N(n2047), .Y(top_core_KE_n4053) );
  OAI2BB2X1 U24970 ( .B0(n1404), .B1(n2058), .A0N(top_core_KE_key_mem_11__95_), 
        .A1N(n2066), .Y(top_core_KE_n4182) );
  OAI2BB2X1 U24971 ( .B0(n1404), .B1(n2078), .A0N(top_core_KE_key_mem_12__95_), 
        .A1N(n2086), .Y(top_core_KE_n4311) );
  OAI2BB2X1 U24972 ( .B0(n1404), .B1(n2098), .A0N(top_core_KE_key_mem_13__95_), 
        .A1N(n2106), .Y(top_core_KE_n4440) );
  OAI2BB2X1 U24973 ( .B0(n1404), .B1(n2118), .A0N(top_core_KE_key_mem_14__95_), 
        .A1N(n2126), .Y(top_core_KE_n4569) );
  OAI2BB2X1 U24974 ( .B0(n1405), .B1(n1858), .A0N(top_core_KE_key_mem_1__94_), 
        .A1N(n1869), .Y(top_core_KE_n2893) );
  OAI2BB2X1 U24975 ( .B0(n1405), .B1(n1879), .A0N(top_core_KE_key_mem_2__94_), 
        .A1N(n1887), .Y(top_core_KE_n3022) );
  OAI2BB2X1 U24976 ( .B0(n1405), .B1(n1908), .A0N(top_core_KE_key_mem_3__94_), 
        .A1N(n1906), .Y(top_core_KE_n3151) );
  OAI2BB2X1 U24977 ( .B0(n1405), .B1(n1919), .A0N(top_core_KE_key_mem_4__94_), 
        .A1N(n1927), .Y(top_core_KE_n3280) );
  OAI2BB2X1 U24978 ( .B0(n1405), .B1(n1938), .A0N(top_core_KE_key_mem_5__94_), 
        .A1N(n1946), .Y(top_core_KE_n3409) );
  OAI2BB2X1 U24979 ( .B0(n1405), .B1(n1959), .A0N(top_core_KE_key_mem_6__94_), 
        .A1N(n1967), .Y(top_core_KE_n3538) );
  OAI2BB2X1 U24980 ( .B0(n1405), .B1(n1978), .A0N(top_core_KE_key_mem_7__94_), 
        .A1N(n1986), .Y(top_core_KE_n3667) );
  OAI2BB2X1 U24981 ( .B0(n1405), .B1(n2039), .A0N(top_core_KE_key_mem_10__94_), 
        .A1N(n2047), .Y(top_core_KE_n4054) );
  OAI2BB2X1 U24982 ( .B0(n1405), .B1(n2058), .A0N(top_core_KE_key_mem_11__94_), 
        .A1N(n2066), .Y(top_core_KE_n4183) );
  OAI2BB2X1 U24983 ( .B0(n1405), .B1(n2078), .A0N(top_core_KE_key_mem_12__94_), 
        .A1N(n2086), .Y(top_core_KE_n4312) );
  OAI2BB2X1 U24984 ( .B0(n1405), .B1(n2098), .A0N(top_core_KE_key_mem_13__94_), 
        .A1N(n2106), .Y(top_core_KE_n4441) );
  OAI2BB2X1 U24985 ( .B0(n1405), .B1(n2118), .A0N(top_core_KE_key_mem_14__94_), 
        .A1N(n2126), .Y(top_core_KE_n4570) );
  OAI2BB2X1 U24986 ( .B0(n1406), .B1(n1858), .A0N(top_core_KE_key_mem_1__93_), 
        .A1N(n1869), .Y(top_core_KE_n2894) );
  OAI2BB2X1 U24987 ( .B0(n1406), .B1(n1878), .A0N(top_core_KE_key_mem_2__93_), 
        .A1N(n1887), .Y(top_core_KE_n3023) );
  OAI2BB2X1 U24988 ( .B0(n1406), .B1(n1898), .A0N(top_core_KE_key_mem_3__93_), 
        .A1N(n1906), .Y(top_core_KE_n3152) );
  OAI2BB2X1 U24989 ( .B0(n1406), .B1(n1918), .A0N(top_core_KE_key_mem_4__93_), 
        .A1N(n1927), .Y(top_core_KE_n3281) );
  OAI2BB2X1 U24990 ( .B0(n1406), .B1(n1948), .A0N(top_core_KE_key_mem_5__93_), 
        .A1N(n1946), .Y(top_core_KE_n3410) );
  OAI2BB2X1 U24991 ( .B0(n1406), .B1(n1958), .A0N(top_core_KE_key_mem_6__93_), 
        .A1N(n1967), .Y(top_core_KE_n3539) );
  OAI2BB2X1 U24992 ( .B0(n1406), .B1(n1977), .A0N(top_core_KE_key_mem_7__93_), 
        .A1N(n1986), .Y(top_core_KE_n3668) );
  OAI2BB2X1 U24993 ( .B0(n1406), .B1(n2038), .A0N(top_core_KE_key_mem_10__93_), 
        .A1N(n2047), .Y(top_core_KE_n4055) );
  OAI2BB2X1 U24994 ( .B0(n1406), .B1(n2057), .A0N(top_core_KE_key_mem_11__93_), 
        .A1N(n2066), .Y(top_core_KE_n4184) );
  OAI2BB2X1 U24995 ( .B0(n1406), .B1(n2088), .A0N(top_core_KE_key_mem_12__93_), 
        .A1N(n2086), .Y(top_core_KE_n4313) );
  OAI2BB2X1 U24996 ( .B0(n1406), .B1(n2097), .A0N(top_core_KE_key_mem_13__93_), 
        .A1N(n2106), .Y(top_core_KE_n4442) );
  OAI2BB2X1 U24997 ( .B0(n1406), .B1(n2117), .A0N(top_core_KE_key_mem_14__93_), 
        .A1N(n2126), .Y(top_core_KE_n4571) );
  OAI2BB2X1 U24998 ( .B0(n1407), .B1(n1858), .A0N(top_core_KE_key_mem_1__92_), 
        .A1N(n1869), .Y(top_core_KE_n2895) );
  OAI2BB2X1 U24999 ( .B0(n1407), .B1(n1878), .A0N(top_core_KE_key_mem_2__92_), 
        .A1N(n1887), .Y(top_core_KE_n3024) );
  OAI2BB2X1 U25000 ( .B0(n1407), .B1(n1898), .A0N(top_core_KE_key_mem_3__92_), 
        .A1N(n1906), .Y(top_core_KE_n3153) );
  OAI2BB2X1 U25001 ( .B0(n1407), .B1(n1918), .A0N(top_core_KE_key_mem_4__92_), 
        .A1N(n1927), .Y(top_core_KE_n3282) );
  OAI2BB2X1 U25002 ( .B0(n1407), .B1(n1949), .A0N(top_core_KE_key_mem_5__92_), 
        .A1N(n1946), .Y(top_core_KE_n3411) );
  OAI2BB2X1 U25003 ( .B0(n1407), .B1(n1958), .A0N(top_core_KE_key_mem_6__92_), 
        .A1N(n1967), .Y(top_core_KE_n3540) );
  OAI2BB2X1 U25004 ( .B0(n1407), .B1(n1977), .A0N(top_core_KE_key_mem_7__92_), 
        .A1N(n1986), .Y(top_core_KE_n3669) );
  OAI2BB2X1 U25005 ( .B0(n1407), .B1(n2038), .A0N(top_core_KE_key_mem_10__92_), 
        .A1N(n2047), .Y(top_core_KE_n4056) );
  OAI2BB2X1 U25006 ( .B0(n1407), .B1(n2057), .A0N(top_core_KE_key_mem_11__92_), 
        .A1N(n2066), .Y(top_core_KE_n4185) );
  OAI2BB2X1 U25007 ( .B0(n1407), .B1(n2089), .A0N(top_core_KE_key_mem_12__92_), 
        .A1N(n2086), .Y(top_core_KE_n4314) );
  OAI2BB2X1 U25008 ( .B0(n1407), .B1(n2097), .A0N(top_core_KE_key_mem_13__92_), 
        .A1N(n2106), .Y(top_core_KE_n4443) );
  OAI2BB2X1 U25009 ( .B0(n1407), .B1(n2117), .A0N(top_core_KE_key_mem_14__92_), 
        .A1N(n2126), .Y(top_core_KE_n4572) );
  OAI2BB2X1 U25010 ( .B0(n1408), .B1(n1858), .A0N(top_core_KE_key_mem_1__91_), 
        .A1N(n1869), .Y(top_core_KE_n2896) );
  OAI2BB2X1 U25011 ( .B0(n1408), .B1(n1878), .A0N(top_core_KE_key_mem_2__91_), 
        .A1N(n1887), .Y(top_core_KE_n3025) );
  OAI2BB2X1 U25012 ( .B0(n1408), .B1(n1898), .A0N(top_core_KE_key_mem_3__91_), 
        .A1N(n1906), .Y(top_core_KE_n3154) );
  OAI2BB2X1 U25013 ( .B0(n1408), .B1(n1918), .A0N(top_core_KE_key_mem_4__91_), 
        .A1N(n1927), .Y(top_core_KE_n3283) );
  OAI2BB2X1 U25014 ( .B0(n1408), .B1(n1952), .A0N(top_core_KE_key_mem_5__91_), 
        .A1N(n1946), .Y(top_core_KE_n3412) );
  OAI2BB2X1 U25015 ( .B0(n1408), .B1(n1958), .A0N(top_core_KE_key_mem_6__91_), 
        .A1N(n1967), .Y(top_core_KE_n3541) );
  OAI2BB2X1 U25016 ( .B0(n1408), .B1(n1977), .A0N(top_core_KE_key_mem_7__91_), 
        .A1N(n1986), .Y(top_core_KE_n3670) );
  OAI2BB2X1 U25017 ( .B0(n1408), .B1(n2038), .A0N(top_core_KE_key_mem_10__91_), 
        .A1N(n2047), .Y(top_core_KE_n4057) );
  OAI2BB2X1 U25018 ( .B0(n1408), .B1(n2057), .A0N(top_core_KE_key_mem_11__91_), 
        .A1N(n2066), .Y(top_core_KE_n4186) );
  OAI2BB2X1 U25019 ( .B0(n1408), .B1(n2092), .A0N(top_core_KE_key_mem_12__91_), 
        .A1N(n2086), .Y(top_core_KE_n4315) );
  OAI2BB2X1 U25020 ( .B0(n1408), .B1(n2097), .A0N(top_core_KE_key_mem_13__91_), 
        .A1N(n2106), .Y(top_core_KE_n4444) );
  OAI2BB2X1 U25021 ( .B0(n1408), .B1(n2117), .A0N(top_core_KE_key_mem_14__91_), 
        .A1N(n2126), .Y(top_core_KE_n4573) );
  OAI2BB2X1 U25022 ( .B0(n1409), .B1(n1858), .A0N(top_core_KE_key_mem_1__90_), 
        .A1N(n1869), .Y(top_core_KE_n2897) );
  OAI2BB2X1 U25023 ( .B0(n1409), .B1(n1878), .A0N(top_core_KE_key_mem_2__90_), 
        .A1N(n1887), .Y(top_core_KE_n3026) );
  OAI2BB2X1 U25024 ( .B0(n1409), .B1(n1898), .A0N(top_core_KE_key_mem_3__90_), 
        .A1N(n1906), .Y(top_core_KE_n3155) );
  OAI2BB2X1 U25025 ( .B0(n1409), .B1(n1918), .A0N(top_core_KE_key_mem_4__90_), 
        .A1N(n1927), .Y(top_core_KE_n3284) );
  OAI2BB2X1 U25026 ( .B0(n1409), .B1(n1946), .A0N(top_core_KE_key_mem_5__90_), 
        .A1N(n1946), .Y(top_core_KE_n3413) );
  OAI2BB2X1 U25027 ( .B0(n1409), .B1(n1958), .A0N(top_core_KE_key_mem_6__90_), 
        .A1N(n1967), .Y(top_core_KE_n3542) );
  OAI2BB2X1 U25028 ( .B0(n1409), .B1(n1977), .A0N(top_core_KE_key_mem_7__90_), 
        .A1N(n1986), .Y(top_core_KE_n3671) );
  OAI2BB2X1 U25029 ( .B0(n1409), .B1(n2038), .A0N(top_core_KE_key_mem_10__90_), 
        .A1N(n2047), .Y(top_core_KE_n4058) );
  OAI2BB2X1 U25030 ( .B0(n1409), .B1(n2057), .A0N(top_core_KE_key_mem_11__90_), 
        .A1N(n2066), .Y(top_core_KE_n4187) );
  OAI2BB2X1 U25031 ( .B0(n1409), .B1(n2086), .A0N(top_core_KE_key_mem_12__90_), 
        .A1N(n2086), .Y(top_core_KE_n4316) );
  OAI2BB2X1 U25032 ( .B0(n1409), .B1(n2097), .A0N(top_core_KE_key_mem_13__90_), 
        .A1N(n2106), .Y(top_core_KE_n4445) );
  OAI2BB2X1 U25033 ( .B0(n1409), .B1(n2117), .A0N(top_core_KE_key_mem_14__90_), 
        .A1N(n2126), .Y(top_core_KE_n4574) );
  OAI2BB2X1 U25034 ( .B0(n1410), .B1(n1859), .A0N(top_core_KE_key_mem_1__89_), 
        .A1N(n1870), .Y(top_core_KE_n2898) );
  OAI2BB2X1 U25035 ( .B0(n1410), .B1(n1877), .A0N(top_core_KE_key_mem_2__89_), 
        .A1N(n1888), .Y(top_core_KE_n3027) );
  OAI2BB2X1 U25036 ( .B0(n1410), .B1(n1897), .A0N(top_core_KE_key_mem_3__89_), 
        .A1N(n1907), .Y(top_core_KE_n3156) );
  OAI2BB2X1 U25037 ( .B0(n1410), .B1(n1917), .A0N(top_core_KE_key_mem_4__89_), 
        .A1N(n1928), .Y(top_core_KE_n3285) );
  OAI2BB2X1 U25038 ( .B0(n1410), .B1(n1937), .A0N(top_core_KE_key_mem_5__89_), 
        .A1N(n1947), .Y(top_core_KE_n3414) );
  OAI2BB2X1 U25039 ( .B0(n1410), .B1(n1957), .A0N(top_core_KE_key_mem_6__89_), 
        .A1N(n1960), .Y(top_core_KE_n3543) );
  OAI2BB2X1 U25040 ( .B0(n1410), .B1(n1977), .A0N(top_core_KE_key_mem_7__89_), 
        .A1N(n1987), .Y(top_core_KE_n3672) );
  OAI2BB2X1 U25041 ( .B0(n1410), .B1(n2037), .A0N(top_core_KE_key_mem_10__89_), 
        .A1N(n2048), .Y(top_core_KE_n4059) );
  OAI2BB2X1 U25042 ( .B0(n1410), .B1(n2057), .A0N(top_core_KE_key_mem_11__89_), 
        .A1N(n2067), .Y(top_core_KE_n4188) );
  OAI2BB2X1 U25043 ( .B0(n1410), .B1(n2077), .A0N(top_core_KE_key_mem_12__89_), 
        .A1N(n2087), .Y(top_core_KE_n4317) );
  OAI2BB2X1 U25044 ( .B0(n1410), .B1(n2097), .A0N(top_core_KE_key_mem_13__89_), 
        .A1N(n2107), .Y(top_core_KE_n4446) );
  OAI2BB2X1 U25045 ( .B0(n1410), .B1(n2117), .A0N(top_core_KE_key_mem_14__89_), 
        .A1N(n2127), .Y(top_core_KE_n4575) );
  OAI2BB2X1 U25046 ( .B0(n1411), .B1(n1859), .A0N(top_core_KE_key_mem_1__88_), 
        .A1N(n1870), .Y(top_core_KE_n2899) );
  OAI2BB2X1 U25047 ( .B0(n1411), .B1(n1877), .A0N(top_core_KE_key_mem_2__88_), 
        .A1N(n1888), .Y(top_core_KE_n3028) );
  OAI2BB2X1 U25048 ( .B0(n1411), .B1(n1897), .A0N(top_core_KE_key_mem_3__88_), 
        .A1N(n1907), .Y(top_core_KE_n3157) );
  OAI2BB2X1 U25049 ( .B0(n1411), .B1(n1917), .A0N(top_core_KE_key_mem_4__88_), 
        .A1N(n1928), .Y(top_core_KE_n3286) );
  OAI2BB2X1 U25050 ( .B0(n1411), .B1(n1937), .A0N(top_core_KE_key_mem_5__88_), 
        .A1N(n1947), .Y(top_core_KE_n3415) );
  OAI2BB2X1 U25051 ( .B0(n1411), .B1(n1957), .A0N(top_core_KE_key_mem_6__88_), 
        .A1N(n1959), .Y(top_core_KE_n3544) );
  OAI2BB2X1 U25052 ( .B0(n1411), .B1(n1979), .A0N(top_core_KE_key_mem_7__88_), 
        .A1N(n1987), .Y(top_core_KE_n3673) );
  OAI2BB2X1 U25053 ( .B0(n1411), .B1(n2037), .A0N(top_core_KE_key_mem_10__88_), 
        .A1N(n2048), .Y(top_core_KE_n4060) );
  OAI2BB2X1 U25054 ( .B0(n1411), .B1(n2059), .A0N(top_core_KE_key_mem_11__88_), 
        .A1N(n2067), .Y(top_core_KE_n4189) );
  OAI2BB2X1 U25055 ( .B0(n1411), .B1(n2077), .A0N(top_core_KE_key_mem_12__88_), 
        .A1N(n2087), .Y(top_core_KE_n4318) );
  OAI2BB2X1 U25056 ( .B0(n1411), .B1(n2099), .A0N(top_core_KE_key_mem_13__88_), 
        .A1N(n2107), .Y(top_core_KE_n4447) );
  OAI2BB2X1 U25057 ( .B0(n1411), .B1(n2119), .A0N(top_core_KE_key_mem_14__88_), 
        .A1N(n2127), .Y(top_core_KE_n4576) );
  OAI2BB2X1 U25058 ( .B0(n1436), .B1(n1862), .A0N(top_core_KE_key_mem_1__63_), 
        .A1N(n1872), .Y(top_core_KE_n2924) );
  OAI2BB2X1 U25059 ( .B0(n1436), .B1(n1879), .A0N(top_core_KE_key_mem_2__63_), 
        .A1N(n1890), .Y(top_core_KE_n3053) );
  OAI2BB2X1 U25060 ( .B0(n1436), .B1(n1904), .A0N(top_core_KE_key_mem_3__63_), 
        .A1N(n1909), .Y(top_core_KE_n3182) );
  OAI2BB2X1 U25061 ( .B0(n1436), .B1(n1919), .A0N(top_core_KE_key_mem_4__63_), 
        .A1N(n1930), .Y(top_core_KE_n3311) );
  OAI2BB2X1 U25062 ( .B0(n1436), .B1(n1938), .A0N(top_core_KE_key_mem_5__63_), 
        .A1N(n1949), .Y(top_core_KE_n3440) );
  OAI2BB2X1 U25063 ( .B0(n1436), .B1(n1959), .A0N(top_core_KE_key_mem_6__63_), 
        .A1N(n1969), .Y(top_core_KE_n3569) );
  OAI2BB2X1 U25064 ( .B0(n1436), .B1(n1978), .A0N(top_core_KE_key_mem_7__63_), 
        .A1N(n1989), .Y(top_core_KE_n3698) );
  OAI2BB2X1 U25065 ( .B0(n1436), .B1(n2039), .A0N(top_core_KE_key_mem_10__63_), 
        .A1N(n2049), .Y(top_core_KE_n4085) );
  OAI2BB2X1 U25066 ( .B0(n1436), .B1(n2058), .A0N(top_core_KE_key_mem_11__63_), 
        .A1N(n2069), .Y(top_core_KE_n4214) );
  OAI2BB2X1 U25067 ( .B0(n1436), .B1(n2078), .A0N(top_core_KE_key_mem_12__63_), 
        .A1N(n2089), .Y(top_core_KE_n4343) );
  OAI2BB2X1 U25068 ( .B0(n1436), .B1(n2098), .A0N(top_core_KE_key_mem_13__63_), 
        .A1N(n2109), .Y(top_core_KE_n4472) );
  OAI2BB2X1 U25069 ( .B0(n1436), .B1(n2118), .A0N(top_core_KE_key_mem_14__63_), 
        .A1N(n2129), .Y(top_core_KE_n4601) );
  OAI2BB2X1 U25070 ( .B0(n1437), .B1(n1861), .A0N(top_core_KE_key_mem_1__62_), 
        .A1N(n1872), .Y(top_core_KE_n2925) );
  OAI2BB2X1 U25071 ( .B0(n1437), .B1(n1879), .A0N(top_core_KE_key_mem_2__62_), 
        .A1N(n1890), .Y(top_core_KE_n3054) );
  OAI2BB2X1 U25072 ( .B0(n1437), .B1(n1901), .A0N(top_core_KE_key_mem_3__62_), 
        .A1N(n1909), .Y(top_core_KE_n3183) );
  OAI2BB2X1 U25073 ( .B0(n1437), .B1(n1919), .A0N(top_core_KE_key_mem_4__62_), 
        .A1N(n1931), .Y(top_core_KE_n3312) );
  OAI2BB2X1 U25074 ( .B0(n1437), .B1(n1938), .A0N(top_core_KE_key_mem_5__62_), 
        .A1N(n1949), .Y(top_core_KE_n3441) );
  OAI2BB2X1 U25075 ( .B0(n1437), .B1(n1959), .A0N(top_core_KE_key_mem_6__62_), 
        .A1N(n1969), .Y(top_core_KE_n3570) );
  OAI2BB2X1 U25076 ( .B0(n1437), .B1(n1978), .A0N(top_core_KE_key_mem_7__62_), 
        .A1N(n1989), .Y(top_core_KE_n3699) );
  OAI2BB2X1 U25077 ( .B0(n1437), .B1(n2039), .A0N(top_core_KE_key_mem_10__62_), 
        .A1N(n2049), .Y(top_core_KE_n4086) );
  OAI2BB2X1 U25078 ( .B0(n1437), .B1(n2058), .A0N(top_core_KE_key_mem_11__62_), 
        .A1N(n2069), .Y(top_core_KE_n4215) );
  OAI2BB2X1 U25079 ( .B0(n1437), .B1(n2078), .A0N(top_core_KE_key_mem_12__62_), 
        .A1N(n2089), .Y(top_core_KE_n4344) );
  OAI2BB2X1 U25080 ( .B0(n1437), .B1(n2098), .A0N(top_core_KE_key_mem_13__62_), 
        .A1N(n2109), .Y(top_core_KE_n4473) );
  OAI2BB2X1 U25081 ( .B0(n1437), .B1(n2118), .A0N(top_core_KE_key_mem_14__62_), 
        .A1N(n2129), .Y(top_core_KE_n4602) );
  OAI2BB2X1 U25082 ( .B0(n1438), .B1(n1861), .A0N(top_core_KE_key_mem_1__61_), 
        .A1N(n1872), .Y(top_core_KE_n2926) );
  OAI2BB2X1 U25083 ( .B0(n1438), .B1(n1882), .A0N(top_core_KE_key_mem_2__61_), 
        .A1N(n1890), .Y(top_core_KE_n3055) );
  OAI2BB2X1 U25084 ( .B0(n1438), .B1(n1901), .A0N(top_core_KE_key_mem_3__61_), 
        .A1N(n1909), .Y(top_core_KE_n3184) );
  OAI2BB2X1 U25085 ( .B0(n1438), .B1(n1922), .A0N(top_core_KE_key_mem_4__61_), 
        .A1N(n1925), .Y(top_core_KE_n3313) );
  OAI2BB2X1 U25086 ( .B0(n1438), .B1(n1941), .A0N(top_core_KE_key_mem_5__61_), 
        .A1N(n1949), .Y(top_core_KE_n3442) );
  OAI2BB2X1 U25087 ( .B0(n1438), .B1(n1962), .A0N(top_core_KE_key_mem_6__61_), 
        .A1N(n1969), .Y(top_core_KE_n3571) );
  OAI2BB2X1 U25088 ( .B0(n1438), .B1(n1981), .A0N(top_core_KE_key_mem_7__61_), 
        .A1N(n1989), .Y(top_core_KE_n3700) );
  OAI2BB2X1 U25089 ( .B0(n1438), .B1(n2042), .A0N(top_core_KE_key_mem_10__61_), 
        .A1N(n2049), .Y(top_core_KE_n4087) );
  OAI2BB2X1 U25090 ( .B0(n1438), .B1(n2061), .A0N(top_core_KE_key_mem_11__61_), 
        .A1N(n2069), .Y(top_core_KE_n4216) );
  OAI2BB2X1 U25091 ( .B0(n1438), .B1(n2081), .A0N(top_core_KE_key_mem_12__61_), 
        .A1N(n2089), .Y(top_core_KE_n4345) );
  OAI2BB2X1 U25092 ( .B0(n1438), .B1(n2101), .A0N(top_core_KE_key_mem_13__61_), 
        .A1N(n2109), .Y(top_core_KE_n4474) );
  OAI2BB2X1 U25093 ( .B0(n1438), .B1(n2121), .A0N(top_core_KE_key_mem_14__61_), 
        .A1N(n2129), .Y(top_core_KE_n4603) );
  OAI2BB2X1 U25094 ( .B0(n1439), .B1(n1861), .A0N(top_core_KE_key_mem_1__60_), 
        .A1N(n1872), .Y(top_core_KE_n2927) );
  OAI2BB2X1 U25095 ( .B0(n1439), .B1(n1883), .A0N(top_core_KE_key_mem_2__60_), 
        .A1N(n1890), .Y(top_core_KE_n3056) );
  OAI2BB2X1 U25096 ( .B0(n1439), .B1(n1902), .A0N(top_core_KE_key_mem_3__60_), 
        .A1N(n1909), .Y(top_core_KE_n3185) );
  OAI2BB2X1 U25097 ( .B0(n1439), .B1(n1923), .A0N(top_core_KE_key_mem_4__60_), 
        .A1N(n1922), .Y(top_core_KE_n3314) );
  OAI2BB2X1 U25098 ( .B0(n1439), .B1(n1942), .A0N(top_core_KE_key_mem_5__60_), 
        .A1N(n1949), .Y(top_core_KE_n3443) );
  OAI2BB2X1 U25099 ( .B0(n1439), .B1(n1963), .A0N(top_core_KE_key_mem_6__60_), 
        .A1N(n1969), .Y(top_core_KE_n3572) );
  OAI2BB2X1 U25100 ( .B0(n1439), .B1(n1982), .A0N(top_core_KE_key_mem_7__60_), 
        .A1N(n1989), .Y(top_core_KE_n3701) );
  OAI2BB2X1 U25101 ( .B0(n1439), .B1(n2043), .A0N(top_core_KE_key_mem_10__60_), 
        .A1N(n2049), .Y(top_core_KE_n4088) );
  OAI2BB2X1 U25102 ( .B0(n1439), .B1(n2062), .A0N(top_core_KE_key_mem_11__60_), 
        .A1N(n2069), .Y(top_core_KE_n4217) );
  OAI2BB2X1 U25103 ( .B0(n1439), .B1(n2082), .A0N(top_core_KE_key_mem_12__60_), 
        .A1N(n2089), .Y(top_core_KE_n4346) );
  OAI2BB2X1 U25104 ( .B0(n1439), .B1(n2102), .A0N(top_core_KE_key_mem_13__60_), 
        .A1N(n2109), .Y(top_core_KE_n4475) );
  OAI2BB2X1 U25105 ( .B0(n1439), .B1(n2122), .A0N(top_core_KE_key_mem_14__60_), 
        .A1N(n2129), .Y(top_core_KE_n4604) );
  OAI2BB2X1 U25106 ( .B0(n1440), .B1(n1861), .A0N(top_core_KE_key_mem_1__59_), 
        .A1N(n1870), .Y(top_core_KE_n2928) );
  OAI2BB2X1 U25107 ( .B0(n1440), .B1(top_core_KE_n874), .A0N(
        top_core_KE_key_mem_2__59_), .A1N(n1890), .Y(top_core_KE_n3057) );
  OAI2BB2X1 U25108 ( .B0(n1440), .B1(top_core_KE_n876), .A0N(
        top_core_KE_key_mem_3__59_), .A1N(n1909), .Y(top_core_KE_n3186) );
  OAI2BB2X1 U25109 ( .B0(n1440), .B1(top_core_KE_n877), .A0N(
        top_core_KE_key_mem_4__59_), .A1N(n1923), .Y(top_core_KE_n3315) );
  OAI2BB2X1 U25110 ( .B0(n1440), .B1(top_core_KE_n879), .A0N(
        top_core_KE_key_mem_5__59_), .A1N(n1949), .Y(top_core_KE_n3444) );
  OAI2BB2X1 U25111 ( .B0(n1440), .B1(top_core_KE_n880), .A0N(
        top_core_KE_key_mem_6__59_), .A1N(n1969), .Y(top_core_KE_n3573) );
  OAI2BB2X1 U25112 ( .B0(n1440), .B1(top_core_KE_n881), .A0N(
        top_core_KE_key_mem_7__59_), .A1N(n1989), .Y(top_core_KE_n3702) );
  OAI2BB2X1 U25113 ( .B0(n1440), .B1(top_core_KE_n886), .A0N(
        top_core_KE_key_mem_10__59_), .A1N(n2049), .Y(top_core_KE_n4089) );
  OAI2BB2X1 U25114 ( .B0(n1440), .B1(top_core_KE_n888), .A0N(
        top_core_KE_key_mem_11__59_), .A1N(n2069), .Y(top_core_KE_n4218) );
  OAI2BB2X1 U25115 ( .B0(n1440), .B1(top_core_KE_n889), .A0N(
        top_core_KE_key_mem_12__59_), .A1N(n2089), .Y(top_core_KE_n4347) );
  OAI2BB2X1 U25116 ( .B0(n1440), .B1(top_core_KE_n890), .A0N(
        top_core_KE_key_mem_13__59_), .A1N(n2109), .Y(top_core_KE_n4476) );
  OAI2BB2X1 U25117 ( .B0(n1440), .B1(top_core_KE_n891), .A0N(
        top_core_KE_key_mem_14__59_), .A1N(n2129), .Y(top_core_KE_n4605) );
  OAI2BB2X1 U25118 ( .B0(n1441), .B1(n1861), .A0N(top_core_KE_key_mem_1__58_), 
        .A1N(n1869), .Y(top_core_KE_n2929) );
  OAI2BB2X1 U25119 ( .B0(n1441), .B1(n1881), .A0N(top_core_KE_key_mem_2__58_), 
        .A1N(n1890), .Y(top_core_KE_n3058) );
  OAI2BB2X1 U25120 ( .B0(n1441), .B1(n1900), .A0N(top_core_KE_key_mem_3__58_), 
        .A1N(n1909), .Y(top_core_KE_n3187) );
  OAI2BB2X1 U25121 ( .B0(n1441), .B1(n1921), .A0N(top_core_KE_key_mem_4__58_), 
        .A1N(n1921), .Y(top_core_KE_n3316) );
  OAI2BB2X1 U25122 ( .B0(n1441), .B1(n1940), .A0N(top_core_KE_key_mem_5__58_), 
        .A1N(n1949), .Y(top_core_KE_n3445) );
  OAI2BB2X1 U25123 ( .B0(n1441), .B1(n1961), .A0N(top_core_KE_key_mem_6__58_), 
        .A1N(n1969), .Y(top_core_KE_n3574) );
  OAI2BB2X1 U25124 ( .B0(n1441), .B1(n1980), .A0N(top_core_KE_key_mem_7__58_), 
        .A1N(n1989), .Y(top_core_KE_n3703) );
  OAI2BB2X1 U25125 ( .B0(n1441), .B1(n2041), .A0N(top_core_KE_key_mem_10__58_), 
        .A1N(n2049), .Y(top_core_KE_n4090) );
  OAI2BB2X1 U25126 ( .B0(n1441), .B1(n2060), .A0N(top_core_KE_key_mem_11__58_), 
        .A1N(n2069), .Y(top_core_KE_n4219) );
  OAI2BB2X1 U25127 ( .B0(n1441), .B1(n2080), .A0N(top_core_KE_key_mem_12__58_), 
        .A1N(n2089), .Y(top_core_KE_n4348) );
  OAI2BB2X1 U25128 ( .B0(n1441), .B1(n2100), .A0N(top_core_KE_key_mem_13__58_), 
        .A1N(n2109), .Y(top_core_KE_n4477) );
  OAI2BB2X1 U25129 ( .B0(n1441), .B1(n2120), .A0N(top_core_KE_key_mem_14__58_), 
        .A1N(n2129), .Y(top_core_KE_n4606) );
  OAI2BB2X1 U25130 ( .B0(n1442), .B1(n1861), .A0N(top_core_KE_key_mem_1__57_), 
        .A1N(n1866), .Y(top_core_KE_n2930) );
  OAI2BB2X1 U25131 ( .B0(n1442), .B1(n1879), .A0N(top_core_KE_key_mem_2__57_), 
        .A1N(n1890), .Y(top_core_KE_n3059) );
  OAI2BB2X1 U25132 ( .B0(n1442), .B1(n1902), .A0N(top_core_KE_key_mem_3__57_), 
        .A1N(n1909), .Y(top_core_KE_n3188) );
  OAI2BB2X1 U25133 ( .B0(n1442), .B1(n1919), .A0N(top_core_KE_key_mem_4__57_), 
        .A1N(n1918), .Y(top_core_KE_n3317) );
  OAI2BB2X1 U25134 ( .B0(n1442), .B1(n1938), .A0N(top_core_KE_key_mem_5__57_), 
        .A1N(n1949), .Y(top_core_KE_n3446) );
  OAI2BB2X1 U25135 ( .B0(n1442), .B1(n1959), .A0N(top_core_KE_key_mem_6__57_), 
        .A1N(n1969), .Y(top_core_KE_n3575) );
  OAI2BB2X1 U25136 ( .B0(n1442), .B1(n1978), .A0N(top_core_KE_key_mem_7__57_), 
        .A1N(n1989), .Y(top_core_KE_n3704) );
  OAI2BB2X1 U25137 ( .B0(n1442), .B1(n2039), .A0N(top_core_KE_key_mem_10__57_), 
        .A1N(n2049), .Y(top_core_KE_n4091) );
  OAI2BB2X1 U25138 ( .B0(n1442), .B1(n2058), .A0N(top_core_KE_key_mem_11__57_), 
        .A1N(n2069), .Y(top_core_KE_n4220) );
  OAI2BB2X1 U25139 ( .B0(n1442), .B1(n2078), .A0N(top_core_KE_key_mem_12__57_), 
        .A1N(n2089), .Y(top_core_KE_n4349) );
  OAI2BB2X1 U25140 ( .B0(n1442), .B1(n2098), .A0N(top_core_KE_key_mem_13__57_), 
        .A1N(n2109), .Y(top_core_KE_n4478) );
  OAI2BB2X1 U25141 ( .B0(n1442), .B1(n2118), .A0N(top_core_KE_key_mem_14__57_), 
        .A1N(n2129), .Y(top_core_KE_n4607) );
  OAI2BB2X1 U25142 ( .B0(n1443), .B1(n1861), .A0N(top_core_KE_key_mem_1__56_), 
        .A1N(n1863), .Y(top_core_KE_n2931) );
  OAI2BB2X1 U25143 ( .B0(n1443), .B1(n1885), .A0N(top_core_KE_key_mem_2__56_), 
        .A1N(n1890), .Y(top_core_KE_n3060) );
  OAI2BB2X1 U25144 ( .B0(n1443), .B1(n1904), .A0N(top_core_KE_key_mem_3__56_), 
        .A1N(n1909), .Y(top_core_KE_n3189) );
  OAI2BB2X1 U25145 ( .B0(n1443), .B1(n1925), .A0N(top_core_KE_key_mem_4__56_), 
        .A1N(n1920), .Y(top_core_KE_n3318) );
  OAI2BB2X1 U25146 ( .B0(n1443), .B1(n1944), .A0N(top_core_KE_key_mem_5__56_), 
        .A1N(n1949), .Y(top_core_KE_n3447) );
  OAI2BB2X1 U25147 ( .B0(n1443), .B1(n1965), .A0N(top_core_KE_key_mem_6__56_), 
        .A1N(n1969), .Y(top_core_KE_n3576) );
  OAI2BB2X1 U25148 ( .B0(n1443), .B1(n1984), .A0N(top_core_KE_key_mem_7__56_), 
        .A1N(n1989), .Y(top_core_KE_n3705) );
  OAI2BB2X1 U25149 ( .B0(n1443), .B1(n2045), .A0N(top_core_KE_key_mem_10__56_), 
        .A1N(n2049), .Y(top_core_KE_n4092) );
  OAI2BB2X1 U25150 ( .B0(n1443), .B1(n2064), .A0N(top_core_KE_key_mem_11__56_), 
        .A1N(n2069), .Y(top_core_KE_n4221) );
  OAI2BB2X1 U25151 ( .B0(n1443), .B1(n2084), .A0N(top_core_KE_key_mem_12__56_), 
        .A1N(n2089), .Y(top_core_KE_n4350) );
  OAI2BB2X1 U25152 ( .B0(n1443), .B1(n2104), .A0N(top_core_KE_key_mem_13__56_), 
        .A1N(n2109), .Y(top_core_KE_n4479) );
  OAI2BB2X1 U25153 ( .B0(n1443), .B1(n2124), .A0N(top_core_KE_key_mem_14__56_), 
        .A1N(n2129), .Y(top_core_KE_n4608) );
  OAI2BB2X1 U25154 ( .B0(n1444), .B1(n1861), .A0N(top_core_KE_key_mem_1__55_), 
        .A1N(n1860), .Y(top_core_KE_n2932) );
  OAI2BB2X1 U25155 ( .B0(n1444), .B1(n1878), .A0N(top_core_KE_key_mem_2__55_), 
        .A1N(n1890), .Y(top_core_KE_n3061) );
  OAI2BB2X1 U25156 ( .B0(n1444), .B1(n1898), .A0N(top_core_KE_key_mem_3__55_), 
        .A1N(n1909), .Y(top_core_KE_n3190) );
  OAI2BB2X1 U25157 ( .B0(n1444), .B1(n1918), .A0N(top_core_KE_key_mem_4__55_), 
        .A1N(n1919), .Y(top_core_KE_n3319) );
  OAI2BB2X1 U25158 ( .B0(n1444), .B1(n1938), .A0N(top_core_KE_key_mem_5__55_), 
        .A1N(n1949), .Y(top_core_KE_n3448) );
  OAI2BB2X1 U25159 ( .B0(n1444), .B1(n1958), .A0N(top_core_KE_key_mem_6__55_), 
        .A1N(n1969), .Y(top_core_KE_n3577) );
  OAI2BB2X1 U25160 ( .B0(n1444), .B1(n1977), .A0N(top_core_KE_key_mem_7__55_), 
        .A1N(n1989), .Y(top_core_KE_n3706) );
  OAI2BB2X1 U25161 ( .B0(n1444), .B1(n2038), .A0N(top_core_KE_key_mem_10__55_), 
        .A1N(n2049), .Y(top_core_KE_n4093) );
  OAI2BB2X1 U25162 ( .B0(n1444), .B1(n2057), .A0N(top_core_KE_key_mem_11__55_), 
        .A1N(n2069), .Y(top_core_KE_n4222) );
  OAI2BB2X1 U25163 ( .B0(n1444), .B1(n2078), .A0N(top_core_KE_key_mem_12__55_), 
        .A1N(n2089), .Y(top_core_KE_n4351) );
  OAI2BB2X1 U25164 ( .B0(n1444), .B1(n2097), .A0N(top_core_KE_key_mem_13__55_), 
        .A1N(n2109), .Y(top_core_KE_n4480) );
  OAI2BB2X1 U25165 ( .B0(n1444), .B1(n2117), .A0N(top_core_KE_key_mem_14__55_), 
        .A1N(n2129), .Y(top_core_KE_n4609) );
  OAI2BB2X1 U25166 ( .B0(n1445), .B1(n1861), .A0N(top_core_KE_key_mem_1__54_), 
        .A1N(n1859), .Y(top_core_KE_n2933) );
  OAI2BB2X1 U25167 ( .B0(n1445), .B1(n1880), .A0N(top_core_KE_key_mem_2__54_), 
        .A1N(n1890), .Y(top_core_KE_n3062) );
  OAI2BB2X1 U25168 ( .B0(n1445), .B1(n1899), .A0N(top_core_KE_key_mem_3__54_), 
        .A1N(n1909), .Y(top_core_KE_n3191) );
  OAI2BB2X1 U25169 ( .B0(n1445), .B1(n1920), .A0N(top_core_KE_key_mem_4__54_), 
        .A1N(n1917), .Y(top_core_KE_n3320) );
  OAI2BB2X1 U25170 ( .B0(n1445), .B1(n1939), .A0N(top_core_KE_key_mem_5__54_), 
        .A1N(n1949), .Y(top_core_KE_n3449) );
  OAI2BB2X1 U25171 ( .B0(n1445), .B1(n1960), .A0N(top_core_KE_key_mem_6__54_), 
        .A1N(n1969), .Y(top_core_KE_n3578) );
  OAI2BB2X1 U25172 ( .B0(n1445), .B1(n1979), .A0N(top_core_KE_key_mem_7__54_), 
        .A1N(n1989), .Y(top_core_KE_n3707) );
  OAI2BB2X1 U25173 ( .B0(n1445), .B1(n2040), .A0N(top_core_KE_key_mem_10__54_), 
        .A1N(n2049), .Y(top_core_KE_n4094) );
  OAI2BB2X1 U25174 ( .B0(n1445), .B1(n2059), .A0N(top_core_KE_key_mem_11__54_), 
        .A1N(n2069), .Y(top_core_KE_n4223) );
  OAI2BB2X1 U25175 ( .B0(n1445), .B1(n2079), .A0N(top_core_KE_key_mem_12__54_), 
        .A1N(n2089), .Y(top_core_KE_n4352) );
  OAI2BB2X1 U25176 ( .B0(n1445), .B1(n2099), .A0N(top_core_KE_key_mem_13__54_), 
        .A1N(n2109), .Y(top_core_KE_n4481) );
  OAI2BB2X1 U25177 ( .B0(n1445), .B1(n2119), .A0N(top_core_KE_key_mem_14__54_), 
        .A1N(n2129), .Y(top_core_KE_n4610) );
  OAI2BB2X1 U25178 ( .B0(n1446), .B1(n1861), .A0N(top_core_KE_key_mem_1__53_), 
        .A1N(n1864), .Y(top_core_KE_n2934) );
  OAI2BB2X1 U25179 ( .B0(n1446), .B1(n1880), .A0N(top_core_KE_key_mem_2__53_), 
        .A1N(n1890), .Y(top_core_KE_n3063) );
  OAI2BB2X1 U25180 ( .B0(n1446), .B1(n1899), .A0N(top_core_KE_key_mem_3__53_), 
        .A1N(n1909), .Y(top_core_KE_n3192) );
  OAI2BB2X1 U25181 ( .B0(n1446), .B1(n1920), .A0N(top_core_KE_key_mem_4__53_), 
        .A1N(n1924), .Y(top_core_KE_n3321) );
  OAI2BB2X1 U25182 ( .B0(n1446), .B1(n1939), .A0N(top_core_KE_key_mem_5__53_), 
        .A1N(n1949), .Y(top_core_KE_n3450) );
  OAI2BB2X1 U25183 ( .B0(n1446), .B1(n1960), .A0N(top_core_KE_key_mem_6__53_), 
        .A1N(n1969), .Y(top_core_KE_n3579) );
  OAI2BB2X1 U25184 ( .B0(n1446), .B1(n1979), .A0N(top_core_KE_key_mem_7__53_), 
        .A1N(n1989), .Y(top_core_KE_n3708) );
  OAI2BB2X1 U25185 ( .B0(n1446), .B1(n2040), .A0N(top_core_KE_key_mem_10__53_), 
        .A1N(n2049), .Y(top_core_KE_n4095) );
  OAI2BB2X1 U25186 ( .B0(n1446), .B1(n2059), .A0N(top_core_KE_key_mem_11__53_), 
        .A1N(n2069), .Y(top_core_KE_n4224) );
  OAI2BB2X1 U25187 ( .B0(n1446), .B1(n2079), .A0N(top_core_KE_key_mem_12__53_), 
        .A1N(n2089), .Y(top_core_KE_n4353) );
  OAI2BB2X1 U25188 ( .B0(n1446), .B1(n2099), .A0N(top_core_KE_key_mem_13__53_), 
        .A1N(n2109), .Y(top_core_KE_n4482) );
  OAI2BB2X1 U25189 ( .B0(n1446), .B1(n2119), .A0N(top_core_KE_key_mem_14__53_), 
        .A1N(n2129), .Y(top_core_KE_n4611) );
  OAI2BB2X1 U25190 ( .B0(n1447), .B1(n1861), .A0N(top_core_KE_key_mem_1__52_), 
        .A1N(n1862), .Y(top_core_KE_n2935) );
  OAI2BB2X1 U25191 ( .B0(n1447), .B1(n1880), .A0N(top_core_KE_key_mem_2__52_), 
        .A1N(n1890), .Y(top_core_KE_n3064) );
  OAI2BB2X1 U25192 ( .B0(n1447), .B1(n1899), .A0N(top_core_KE_key_mem_3__52_), 
        .A1N(n1909), .Y(top_core_KE_n3193) );
  OAI2BB2X1 U25193 ( .B0(n1447), .B1(n1920), .A0N(top_core_KE_key_mem_4__52_), 
        .A1N(n1929), .Y(top_core_KE_n3322) );
  OAI2BB2X1 U25194 ( .B0(n1447), .B1(n1939), .A0N(top_core_KE_key_mem_5__52_), 
        .A1N(n1949), .Y(top_core_KE_n3451) );
  OAI2BB2X1 U25195 ( .B0(n1447), .B1(n1960), .A0N(top_core_KE_key_mem_6__52_), 
        .A1N(n1969), .Y(top_core_KE_n3580) );
  OAI2BB2X1 U25196 ( .B0(n1447), .B1(n1979), .A0N(top_core_KE_key_mem_7__52_), 
        .A1N(n1989), .Y(top_core_KE_n3709) );
  OAI2BB2X1 U25197 ( .B0(n1447), .B1(n2040), .A0N(top_core_KE_key_mem_10__52_), 
        .A1N(n2049), .Y(top_core_KE_n4096) );
  OAI2BB2X1 U25198 ( .B0(n1447), .B1(n2059), .A0N(top_core_KE_key_mem_11__52_), 
        .A1N(n2069), .Y(top_core_KE_n4225) );
  OAI2BB2X1 U25199 ( .B0(n1447), .B1(n2079), .A0N(top_core_KE_key_mem_12__52_), 
        .A1N(n2089), .Y(top_core_KE_n4354) );
  OAI2BB2X1 U25200 ( .B0(n1447), .B1(n2099), .A0N(top_core_KE_key_mem_13__52_), 
        .A1N(n2109), .Y(top_core_KE_n4483) );
  OAI2BB2X1 U25201 ( .B0(n1447), .B1(n2119), .A0N(top_core_KE_key_mem_14__52_), 
        .A1N(n2129), .Y(top_core_KE_n4612) );
  OAI2BB2X1 U25202 ( .B0(n1448), .B1(n1861), .A0N(top_core_KE_key_mem_1__51_), 
        .A1N(n1865), .Y(top_core_KE_n2936) );
  OAI2BB2X1 U25203 ( .B0(n1448), .B1(n1880), .A0N(top_core_KE_key_mem_2__51_), 
        .A1N(n1891), .Y(top_core_KE_n3065) );
  OAI2BB2X1 U25204 ( .B0(n1448), .B1(n1899), .A0N(top_core_KE_key_mem_3__51_), 
        .A1N(n1910), .Y(top_core_KE_n3194) );
  OAI2BB2X1 U25205 ( .B0(n1448), .B1(n1920), .A0N(top_core_KE_key_mem_4__51_), 
        .A1N(n1930), .Y(top_core_KE_n3323) );
  OAI2BB2X1 U25206 ( .B0(n1448), .B1(n1939), .A0N(top_core_KE_key_mem_5__51_), 
        .A1N(n1950), .Y(top_core_KE_n3452) );
  OAI2BB2X1 U25207 ( .B0(n1448), .B1(n1960), .A0N(top_core_KE_key_mem_6__51_), 
        .A1N(n1970), .Y(top_core_KE_n3581) );
  OAI2BB2X1 U25208 ( .B0(n1448), .B1(n1979), .A0N(top_core_KE_key_mem_7__51_), 
        .A1N(n1990), .Y(top_core_KE_n3710) );
  OAI2BB2X1 U25209 ( .B0(n1448), .B1(n2040), .A0N(top_core_KE_key_mem_10__51_), 
        .A1N(n2050), .Y(top_core_KE_n4097) );
  OAI2BB2X1 U25210 ( .B0(n1448), .B1(n2059), .A0N(top_core_KE_key_mem_11__51_), 
        .A1N(n2070), .Y(top_core_KE_n4226) );
  OAI2BB2X1 U25211 ( .B0(n1448), .B1(n2079), .A0N(top_core_KE_key_mem_12__51_), 
        .A1N(n2090), .Y(top_core_KE_n4355) );
  OAI2BB2X1 U25212 ( .B0(n1448), .B1(n2099), .A0N(top_core_KE_key_mem_13__51_), 
        .A1N(n2110), .Y(top_core_KE_n4484) );
  OAI2BB2X1 U25213 ( .B0(n1448), .B1(n2119), .A0N(top_core_KE_key_mem_14__51_), 
        .A1N(n2130), .Y(top_core_KE_n4613) );
  OAI2BB2X1 U25214 ( .B0(n1449), .B1(n1862), .A0N(top_core_KE_key_mem_1__50_), 
        .A1N(n1861), .Y(top_core_KE_n2937) );
  OAI2BB2X1 U25215 ( .B0(n1449), .B1(n1880), .A0N(top_core_KE_key_mem_2__50_), 
        .A1N(n1891), .Y(top_core_KE_n3066) );
  OAI2BB2X1 U25216 ( .B0(n1449), .B1(n1899), .A0N(top_core_KE_key_mem_3__50_), 
        .A1N(n1910), .Y(top_core_KE_n3195) );
  OAI2BB2X1 U25217 ( .B0(n1449), .B1(n1920), .A0N(top_core_KE_key_mem_4__50_), 
        .A1N(n1930), .Y(top_core_KE_n3324) );
  OAI2BB2X1 U25218 ( .B0(n1449), .B1(n1939), .A0N(top_core_KE_key_mem_5__50_), 
        .A1N(n1950), .Y(top_core_KE_n3453) );
  OAI2BB2X1 U25219 ( .B0(n1449), .B1(n1960), .A0N(top_core_KE_key_mem_6__50_), 
        .A1N(n1970), .Y(top_core_KE_n3582) );
  OAI2BB2X1 U25220 ( .B0(n1449), .B1(n1979), .A0N(top_core_KE_key_mem_7__50_), 
        .A1N(n1990), .Y(top_core_KE_n3711) );
  OAI2BB2X1 U25221 ( .B0(n1449), .B1(n2040), .A0N(top_core_KE_key_mem_10__50_), 
        .A1N(n2050), .Y(top_core_KE_n4098) );
  OAI2BB2X1 U25222 ( .B0(n1449), .B1(n2059), .A0N(top_core_KE_key_mem_11__50_), 
        .A1N(n2070), .Y(top_core_KE_n4227) );
  OAI2BB2X1 U25223 ( .B0(n1449), .B1(n2079), .A0N(top_core_KE_key_mem_12__50_), 
        .A1N(n2090), .Y(top_core_KE_n4356) );
  OAI2BB2X1 U25224 ( .B0(n1449), .B1(n2099), .A0N(top_core_KE_key_mem_13__50_), 
        .A1N(n2110), .Y(top_core_KE_n4485) );
  OAI2BB2X1 U25225 ( .B0(n1449), .B1(n2119), .A0N(top_core_KE_key_mem_14__50_), 
        .A1N(n2130), .Y(top_core_KE_n4614) );
  OAI2BB2X1 U25226 ( .B0(n1450), .B1(n1862), .A0N(top_core_KE_key_mem_1__49_), 
        .A1N(top_core_KE_n873), .Y(top_core_KE_n2938) );
  OAI2BB2X1 U25227 ( .B0(n1450), .B1(n1880), .A0N(top_core_KE_key_mem_2__49_), 
        .A1N(n1891), .Y(top_core_KE_n3067) );
  OAI2BB2X1 U25228 ( .B0(n1450), .B1(n1899), .A0N(top_core_KE_key_mem_3__49_), 
        .A1N(n1910), .Y(top_core_KE_n3196) );
  OAI2BB2X1 U25229 ( .B0(n1450), .B1(n1920), .A0N(top_core_KE_key_mem_4__49_), 
        .A1N(n1930), .Y(top_core_KE_n3325) );
  OAI2BB2X1 U25230 ( .B0(n1450), .B1(n1939), .A0N(top_core_KE_key_mem_5__49_), 
        .A1N(n1950), .Y(top_core_KE_n3454) );
  OAI2BB2X1 U25231 ( .B0(n1450), .B1(n1960), .A0N(top_core_KE_key_mem_6__49_), 
        .A1N(n1970), .Y(top_core_KE_n3583) );
  OAI2BB2X1 U25232 ( .B0(n1450), .B1(n1979), .A0N(top_core_KE_key_mem_7__49_), 
        .A1N(n1990), .Y(top_core_KE_n3712) );
  OAI2BB2X1 U25233 ( .B0(n1450), .B1(n2040), .A0N(top_core_KE_key_mem_10__49_), 
        .A1N(n2050), .Y(top_core_KE_n4099) );
  OAI2BB2X1 U25234 ( .B0(n1450), .B1(n2059), .A0N(top_core_KE_key_mem_11__49_), 
        .A1N(n2070), .Y(top_core_KE_n4228) );
  OAI2BB2X1 U25235 ( .B0(n1450), .B1(n2079), .A0N(top_core_KE_key_mem_12__49_), 
        .A1N(n2090), .Y(top_core_KE_n4357) );
  OAI2BB2X1 U25236 ( .B0(n1450), .B1(n2099), .A0N(top_core_KE_key_mem_13__49_), 
        .A1N(n2110), .Y(top_core_KE_n4486) );
  OAI2BB2X1 U25237 ( .B0(n1450), .B1(n2119), .A0N(top_core_KE_key_mem_14__49_), 
        .A1N(n2130), .Y(top_core_KE_n4615) );
  OAI2BB2X1 U25238 ( .B0(n1451), .B1(n1862), .A0N(top_core_KE_key_mem_1__48_), 
        .A1N(n1857), .Y(top_core_KE_n2939) );
  OAI2BB2X1 U25239 ( .B0(n1451), .B1(n1880), .A0N(top_core_KE_key_mem_2__48_), 
        .A1N(n1891), .Y(top_core_KE_n3068) );
  OAI2BB2X1 U25240 ( .B0(n1451), .B1(n1899), .A0N(top_core_KE_key_mem_3__48_), 
        .A1N(n1910), .Y(top_core_KE_n3197) );
  OAI2BB2X1 U25241 ( .B0(n1451), .B1(n1920), .A0N(top_core_KE_key_mem_4__48_), 
        .A1N(n1930), .Y(top_core_KE_n3326) );
  OAI2BB2X1 U25242 ( .B0(n1451), .B1(n1939), .A0N(top_core_KE_key_mem_5__48_), 
        .A1N(n1950), .Y(top_core_KE_n3455) );
  OAI2BB2X1 U25243 ( .B0(n1451), .B1(n1960), .A0N(top_core_KE_key_mem_6__48_), 
        .A1N(n1970), .Y(top_core_KE_n3584) );
  OAI2BB2X1 U25244 ( .B0(n1451), .B1(n1979), .A0N(top_core_KE_key_mem_7__48_), 
        .A1N(n1990), .Y(top_core_KE_n3713) );
  OAI2BB2X1 U25245 ( .B0(n1451), .B1(n2040), .A0N(top_core_KE_key_mem_10__48_), 
        .A1N(n2050), .Y(top_core_KE_n4100) );
  OAI2BB2X1 U25246 ( .B0(n1451), .B1(n2059), .A0N(top_core_KE_key_mem_11__48_), 
        .A1N(n2070), .Y(top_core_KE_n4229) );
  OAI2BB2X1 U25247 ( .B0(n1451), .B1(n2079), .A0N(top_core_KE_key_mem_12__48_), 
        .A1N(n2090), .Y(top_core_KE_n4358) );
  OAI2BB2X1 U25248 ( .B0(n1451), .B1(n2099), .A0N(top_core_KE_key_mem_13__48_), 
        .A1N(n2110), .Y(top_core_KE_n4487) );
  OAI2BB2X1 U25249 ( .B0(n1451), .B1(n2119), .A0N(top_core_KE_key_mem_14__48_), 
        .A1N(n2130), .Y(top_core_KE_n4616) );
  OAI2BB2X1 U25250 ( .B0(n1452), .B1(n1862), .A0N(top_core_KE_key_mem_1__47_), 
        .A1N(n1863), .Y(top_core_KE_n2940) );
  OAI2BB2X1 U25251 ( .B0(n1452), .B1(n1880), .A0N(top_core_KE_key_mem_2__47_), 
        .A1N(n1891), .Y(top_core_KE_n3069) );
  OAI2BB2X1 U25252 ( .B0(n1452), .B1(n1899), .A0N(top_core_KE_key_mem_3__47_), 
        .A1N(n1910), .Y(top_core_KE_n3198) );
  OAI2BB2X1 U25253 ( .B0(n1452), .B1(n1920), .A0N(top_core_KE_key_mem_4__47_), 
        .A1N(n1930), .Y(top_core_KE_n3327) );
  OAI2BB2X1 U25254 ( .B0(n1452), .B1(n1939), .A0N(top_core_KE_key_mem_5__47_), 
        .A1N(n1950), .Y(top_core_KE_n3456) );
  OAI2BB2X1 U25255 ( .B0(n1452), .B1(n1960), .A0N(top_core_KE_key_mem_6__47_), 
        .A1N(n1970), .Y(top_core_KE_n3585) );
  OAI2BB2X1 U25256 ( .B0(n1452), .B1(n1979), .A0N(top_core_KE_key_mem_7__47_), 
        .A1N(n1990), .Y(top_core_KE_n3714) );
  OAI2BB2X1 U25257 ( .B0(n1452), .B1(n2040), .A0N(top_core_KE_key_mem_10__47_), 
        .A1N(n2050), .Y(top_core_KE_n4101) );
  OAI2BB2X1 U25258 ( .B0(n1452), .B1(n2059), .A0N(top_core_KE_key_mem_11__47_), 
        .A1N(n2070), .Y(top_core_KE_n4230) );
  OAI2BB2X1 U25259 ( .B0(n1452), .B1(n2079), .A0N(top_core_KE_key_mem_12__47_), 
        .A1N(n2090), .Y(top_core_KE_n4359) );
  OAI2BB2X1 U25260 ( .B0(n1452), .B1(n2099), .A0N(top_core_KE_key_mem_13__47_), 
        .A1N(n2110), .Y(top_core_KE_n4488) );
  OAI2BB2X1 U25261 ( .B0(n1452), .B1(n2119), .A0N(top_core_KE_key_mem_14__47_), 
        .A1N(n2130), .Y(top_core_KE_n4617) );
  OAI2BB2X1 U25262 ( .B0(n1453), .B1(n1862), .A0N(top_core_KE_key_mem_1__46_), 
        .A1N(n1860), .Y(top_core_KE_n2941) );
  OAI2BB2X1 U25263 ( .B0(n1453), .B1(n1880), .A0N(top_core_KE_key_mem_2__46_), 
        .A1N(n1891), .Y(top_core_KE_n3070) );
  OAI2BB2X1 U25264 ( .B0(n1453), .B1(n1899), .A0N(top_core_KE_key_mem_3__46_), 
        .A1N(n1910), .Y(top_core_KE_n3199) );
  OAI2BB2X1 U25265 ( .B0(n1453), .B1(n1920), .A0N(top_core_KE_key_mem_4__46_), 
        .A1N(n1930), .Y(top_core_KE_n3328) );
  OAI2BB2X1 U25266 ( .B0(n1453), .B1(n1939), .A0N(top_core_KE_key_mem_5__46_), 
        .A1N(n1950), .Y(top_core_KE_n3457) );
  OAI2BB2X1 U25267 ( .B0(n1453), .B1(n1960), .A0N(top_core_KE_key_mem_6__46_), 
        .A1N(n1970), .Y(top_core_KE_n3586) );
  OAI2BB2X1 U25268 ( .B0(n1453), .B1(n1979), .A0N(top_core_KE_key_mem_7__46_), 
        .A1N(n1990), .Y(top_core_KE_n3715) );
  OAI2BB2X1 U25269 ( .B0(n1453), .B1(n2040), .A0N(top_core_KE_key_mem_10__46_), 
        .A1N(n2050), .Y(top_core_KE_n4102) );
  OAI2BB2X1 U25270 ( .B0(n1453), .B1(n2059), .A0N(top_core_KE_key_mem_11__46_), 
        .A1N(n2070), .Y(top_core_KE_n4231) );
  OAI2BB2X1 U25271 ( .B0(n1453), .B1(n2079), .A0N(top_core_KE_key_mem_12__46_), 
        .A1N(n2090), .Y(top_core_KE_n4360) );
  OAI2BB2X1 U25272 ( .B0(n1453), .B1(n2099), .A0N(top_core_KE_key_mem_13__46_), 
        .A1N(n2110), .Y(top_core_KE_n4489) );
  OAI2BB2X1 U25273 ( .B0(n1453), .B1(n2119), .A0N(top_core_KE_key_mem_14__46_), 
        .A1N(n2130), .Y(top_core_KE_n4618) );
  OAI2BB2X1 U25274 ( .B0(n1454), .B1(n1862), .A0N(top_core_KE_key_mem_1__45_), 
        .A1N(n1859), .Y(top_core_KE_n2942) );
  OAI2BB2X1 U25275 ( .B0(n1454), .B1(n1881), .A0N(top_core_KE_key_mem_2__45_), 
        .A1N(n1891), .Y(top_core_KE_n3071) );
  OAI2BB2X1 U25276 ( .B0(n1454), .B1(n1900), .A0N(top_core_KE_key_mem_3__45_), 
        .A1N(n1910), .Y(top_core_KE_n3200) );
  OAI2BB2X1 U25277 ( .B0(n1454), .B1(n1921), .A0N(top_core_KE_key_mem_4__45_), 
        .A1N(n1930), .Y(top_core_KE_n3329) );
  OAI2BB2X1 U25278 ( .B0(n1454), .B1(n1940), .A0N(top_core_KE_key_mem_5__45_), 
        .A1N(n1950), .Y(top_core_KE_n3458) );
  OAI2BB2X1 U25279 ( .B0(n1454), .B1(n1961), .A0N(top_core_KE_key_mem_6__45_), 
        .A1N(n1970), .Y(top_core_KE_n3587) );
  OAI2BB2X1 U25280 ( .B0(n1454), .B1(n1980), .A0N(top_core_KE_key_mem_7__45_), 
        .A1N(n1990), .Y(top_core_KE_n3716) );
  OAI2BB2X1 U25281 ( .B0(n1454), .B1(n2041), .A0N(top_core_KE_key_mem_10__45_), 
        .A1N(n2050), .Y(top_core_KE_n4103) );
  OAI2BB2X1 U25282 ( .B0(n1454), .B1(n2060), .A0N(top_core_KE_key_mem_11__45_), 
        .A1N(n2070), .Y(top_core_KE_n4232) );
  OAI2BB2X1 U25283 ( .B0(n1454), .B1(n2080), .A0N(top_core_KE_key_mem_12__45_), 
        .A1N(n2090), .Y(top_core_KE_n4361) );
  OAI2BB2X1 U25284 ( .B0(n1454), .B1(n2100), .A0N(top_core_KE_key_mem_13__45_), 
        .A1N(n2110), .Y(top_core_KE_n4490) );
  OAI2BB2X1 U25285 ( .B0(n1454), .B1(n2120), .A0N(top_core_KE_key_mem_14__45_), 
        .A1N(n2130), .Y(top_core_KE_n4619) );
  OAI2BB2X1 U25286 ( .B0(n1455), .B1(n1862), .A0N(top_core_KE_key_mem_1__44_), 
        .A1N(n1864), .Y(top_core_KE_n2943) );
  OAI2BB2X1 U25287 ( .B0(n1455), .B1(n1881), .A0N(top_core_KE_key_mem_2__44_), 
        .A1N(n1891), .Y(top_core_KE_n3072) );
  OAI2BB2X1 U25288 ( .B0(n1455), .B1(n1900), .A0N(top_core_KE_key_mem_3__44_), 
        .A1N(n1910), .Y(top_core_KE_n3201) );
  OAI2BB2X1 U25289 ( .B0(n1455), .B1(n1921), .A0N(top_core_KE_key_mem_4__44_), 
        .A1N(n1930), .Y(top_core_KE_n3330) );
  OAI2BB2X1 U25290 ( .B0(n1455), .B1(n1940), .A0N(top_core_KE_key_mem_5__44_), 
        .A1N(n1950), .Y(top_core_KE_n3459) );
  OAI2BB2X1 U25291 ( .B0(n1455), .B1(n1961), .A0N(top_core_KE_key_mem_6__44_), 
        .A1N(n1970), .Y(top_core_KE_n3588) );
  OAI2BB2X1 U25292 ( .B0(n1455), .B1(n1980), .A0N(top_core_KE_key_mem_7__44_), 
        .A1N(n1990), .Y(top_core_KE_n3717) );
  OAI2BB2X1 U25293 ( .B0(n1455), .B1(n2041), .A0N(top_core_KE_key_mem_10__44_), 
        .A1N(n2050), .Y(top_core_KE_n4104) );
  OAI2BB2X1 U25294 ( .B0(n1455), .B1(n2060), .A0N(top_core_KE_key_mem_11__44_), 
        .A1N(n2070), .Y(top_core_KE_n4233) );
  OAI2BB2X1 U25295 ( .B0(n1455), .B1(n2080), .A0N(top_core_KE_key_mem_12__44_), 
        .A1N(n2090), .Y(top_core_KE_n4362) );
  OAI2BB2X1 U25296 ( .B0(n1455), .B1(n2100), .A0N(top_core_KE_key_mem_13__44_), 
        .A1N(n2110), .Y(top_core_KE_n4491) );
  OAI2BB2X1 U25297 ( .B0(n1455), .B1(n2120), .A0N(top_core_KE_key_mem_14__44_), 
        .A1N(n2130), .Y(top_core_KE_n4620) );
  OAI2BB2X1 U25298 ( .B0(n1456), .B1(n1862), .A0N(top_core_KE_key_mem_1__43_), 
        .A1N(n1866), .Y(top_core_KE_n2944) );
  OAI2BB2X1 U25299 ( .B0(n1456), .B1(n1881), .A0N(top_core_KE_key_mem_2__43_), 
        .A1N(n1891), .Y(top_core_KE_n3073) );
  OAI2BB2X1 U25300 ( .B0(n1456), .B1(n1900), .A0N(top_core_KE_key_mem_3__43_), 
        .A1N(n1910), .Y(top_core_KE_n3202) );
  OAI2BB2X1 U25301 ( .B0(n1456), .B1(n1921), .A0N(top_core_KE_key_mem_4__43_), 
        .A1N(n1930), .Y(top_core_KE_n3331) );
  OAI2BB2X1 U25302 ( .B0(n1456), .B1(n1940), .A0N(top_core_KE_key_mem_5__43_), 
        .A1N(n1950), .Y(top_core_KE_n3460) );
  OAI2BB2X1 U25303 ( .B0(n1456), .B1(n1961), .A0N(top_core_KE_key_mem_6__43_), 
        .A1N(n1970), .Y(top_core_KE_n3589) );
  OAI2BB2X1 U25304 ( .B0(n1456), .B1(n1980), .A0N(top_core_KE_key_mem_7__43_), 
        .A1N(n1990), .Y(top_core_KE_n3718) );
  OAI2BB2X1 U25305 ( .B0(n1456), .B1(n2041), .A0N(top_core_KE_key_mem_10__43_), 
        .A1N(n2050), .Y(top_core_KE_n4105) );
  OAI2BB2X1 U25306 ( .B0(n1456), .B1(n2060), .A0N(top_core_KE_key_mem_11__43_), 
        .A1N(n2070), .Y(top_core_KE_n4234) );
  OAI2BB2X1 U25307 ( .B0(n1456), .B1(n2080), .A0N(top_core_KE_key_mem_12__43_), 
        .A1N(n2090), .Y(top_core_KE_n4363) );
  OAI2BB2X1 U25308 ( .B0(n1456), .B1(n2100), .A0N(top_core_KE_key_mem_13__43_), 
        .A1N(n2110), .Y(top_core_KE_n4492) );
  OAI2BB2X1 U25309 ( .B0(n1456), .B1(n2120), .A0N(top_core_KE_key_mem_14__43_), 
        .A1N(n2130), .Y(top_core_KE_n4621) );
  OAI2BB2X1 U25310 ( .B0(n1457), .B1(n1862), .A0N(top_core_KE_key_mem_1__42_), 
        .A1N(n1862), .Y(top_core_KE_n2945) );
  OAI2BB2X1 U25311 ( .B0(n1457), .B1(n1881), .A0N(top_core_KE_key_mem_2__42_), 
        .A1N(n1891), .Y(top_core_KE_n3074) );
  OAI2BB2X1 U25312 ( .B0(n1457), .B1(n1900), .A0N(top_core_KE_key_mem_3__42_), 
        .A1N(n1910), .Y(top_core_KE_n3203) );
  OAI2BB2X1 U25313 ( .B0(n1457), .B1(n1921), .A0N(top_core_KE_key_mem_4__42_), 
        .A1N(n1930), .Y(top_core_KE_n3332) );
  OAI2BB2X1 U25314 ( .B0(n1457), .B1(n1940), .A0N(top_core_KE_key_mem_5__42_), 
        .A1N(n1950), .Y(top_core_KE_n3461) );
  OAI2BB2X1 U25315 ( .B0(n1457), .B1(n1961), .A0N(top_core_KE_key_mem_6__42_), 
        .A1N(n1970), .Y(top_core_KE_n3590) );
  OAI2BB2X1 U25316 ( .B0(n1457), .B1(n1980), .A0N(top_core_KE_key_mem_7__42_), 
        .A1N(n1990), .Y(top_core_KE_n3719) );
  OAI2BB2X1 U25317 ( .B0(n1457), .B1(n2041), .A0N(top_core_KE_key_mem_10__42_), 
        .A1N(n2050), .Y(top_core_KE_n4106) );
  OAI2BB2X1 U25318 ( .B0(n1457), .B1(n2060), .A0N(top_core_KE_key_mem_11__42_), 
        .A1N(n2070), .Y(top_core_KE_n4235) );
  OAI2BB2X1 U25319 ( .B0(n1457), .B1(n2080), .A0N(top_core_KE_key_mem_12__42_), 
        .A1N(n2090), .Y(top_core_KE_n4364) );
  OAI2BB2X1 U25320 ( .B0(n1457), .B1(n2100), .A0N(top_core_KE_key_mem_13__42_), 
        .A1N(n2110), .Y(top_core_KE_n4493) );
  OAI2BB2X1 U25321 ( .B0(n1457), .B1(n2120), .A0N(top_core_KE_key_mem_14__42_), 
        .A1N(n2130), .Y(top_core_KE_n4622) );
  OAI2BB2X1 U25322 ( .B0(n1458), .B1(n1862), .A0N(top_core_KE_key_mem_1__41_), 
        .A1N(n1865), .Y(top_core_KE_n2946) );
  OAI2BB2X1 U25323 ( .B0(n1458), .B1(n1881), .A0N(top_core_KE_key_mem_2__41_), 
        .A1N(n1891), .Y(top_core_KE_n3075) );
  OAI2BB2X1 U25324 ( .B0(n1458), .B1(n1900), .A0N(top_core_KE_key_mem_3__41_), 
        .A1N(n1910), .Y(top_core_KE_n3204) );
  OAI2BB2X1 U25325 ( .B0(n1458), .B1(n1921), .A0N(top_core_KE_key_mem_4__41_), 
        .A1N(n1930), .Y(top_core_KE_n3333) );
  OAI2BB2X1 U25326 ( .B0(n1458), .B1(n1940), .A0N(top_core_KE_key_mem_5__41_), 
        .A1N(n1950), .Y(top_core_KE_n3462) );
  OAI2BB2X1 U25327 ( .B0(n1458), .B1(n1961), .A0N(top_core_KE_key_mem_6__41_), 
        .A1N(n1970), .Y(top_core_KE_n3591) );
  OAI2BB2X1 U25328 ( .B0(n1458), .B1(n1980), .A0N(top_core_KE_key_mem_7__41_), 
        .A1N(n1990), .Y(top_core_KE_n3720) );
  OAI2BB2X1 U25329 ( .B0(n1458), .B1(n2041), .A0N(top_core_KE_key_mem_10__41_), 
        .A1N(n2050), .Y(top_core_KE_n4107) );
  OAI2BB2X1 U25330 ( .B0(n1458), .B1(n2060), .A0N(top_core_KE_key_mem_11__41_), 
        .A1N(n2070), .Y(top_core_KE_n4236) );
  OAI2BB2X1 U25331 ( .B0(n1458), .B1(n2080), .A0N(top_core_KE_key_mem_12__41_), 
        .A1N(n2090), .Y(top_core_KE_n4365) );
  OAI2BB2X1 U25332 ( .B0(n1458), .B1(n2100), .A0N(top_core_KE_key_mem_13__41_), 
        .A1N(n2110), .Y(top_core_KE_n4494) );
  OAI2BB2X1 U25333 ( .B0(n1458), .B1(n2120), .A0N(top_core_KE_key_mem_14__41_), 
        .A1N(n2130), .Y(top_core_KE_n4623) );
  OAI2BB2X1 U25334 ( .B0(n1459), .B1(n1863), .A0N(top_core_KE_key_mem_1__40_), 
        .A1N(n1861), .Y(top_core_KE_n2947) );
  OAI2BB2X1 U25335 ( .B0(n1459), .B1(n1881), .A0N(top_core_KE_key_mem_2__40_), 
        .A1N(n1891), .Y(top_core_KE_n3076) );
  OAI2BB2X1 U25336 ( .B0(n1459), .B1(n1900), .A0N(top_core_KE_key_mem_3__40_), 
        .A1N(n1910), .Y(top_core_KE_n3205) );
  OAI2BB2X1 U25337 ( .B0(n1459), .B1(n1921), .A0N(top_core_KE_key_mem_4__40_), 
        .A1N(n1930), .Y(top_core_KE_n3334) );
  OAI2BB2X1 U25338 ( .B0(n1459), .B1(n1940), .A0N(top_core_KE_key_mem_5__40_), 
        .A1N(n1950), .Y(top_core_KE_n3463) );
  OAI2BB2X1 U25339 ( .B0(n1459), .B1(n1961), .A0N(top_core_KE_key_mem_6__40_), 
        .A1N(n1970), .Y(top_core_KE_n3592) );
  OAI2BB2X1 U25340 ( .B0(n1459), .B1(n1980), .A0N(top_core_KE_key_mem_7__40_), 
        .A1N(n1990), .Y(top_core_KE_n3721) );
  OAI2BB2X1 U25341 ( .B0(n1459), .B1(n2041), .A0N(top_core_KE_key_mem_10__40_), 
        .A1N(n2050), .Y(top_core_KE_n4108) );
  OAI2BB2X1 U25342 ( .B0(n1459), .B1(n2060), .A0N(top_core_KE_key_mem_11__40_), 
        .A1N(n2070), .Y(top_core_KE_n4237) );
  OAI2BB2X1 U25343 ( .B0(n1459), .B1(n2080), .A0N(top_core_KE_key_mem_12__40_), 
        .A1N(n2090), .Y(top_core_KE_n4366) );
  OAI2BB2X1 U25344 ( .B0(n1459), .B1(n2100), .A0N(top_core_KE_key_mem_13__40_), 
        .A1N(n2110), .Y(top_core_KE_n4495) );
  OAI2BB2X1 U25345 ( .B0(n1459), .B1(n2120), .A0N(top_core_KE_key_mem_14__40_), 
        .A1N(n2130), .Y(top_core_KE_n4624) );
  OAI2BB2X1 U25346 ( .B0(n1460), .B1(n1863), .A0N(top_core_KE_key_mem_1__39_), 
        .A1N(n1858), .Y(top_core_KE_n2948) );
  OAI2BB2X1 U25347 ( .B0(n1460), .B1(n1881), .A0N(top_core_KE_key_mem_2__39_), 
        .A1N(n1891), .Y(top_core_KE_n3077) );
  OAI2BB2X1 U25348 ( .B0(n1460), .B1(n1900), .A0N(top_core_KE_key_mem_3__39_), 
        .A1N(n1910), .Y(top_core_KE_n3206) );
  OAI2BB2X1 U25349 ( .B0(n1460), .B1(n1921), .A0N(top_core_KE_key_mem_4__39_), 
        .A1N(n1930), .Y(top_core_KE_n3335) );
  OAI2BB2X1 U25350 ( .B0(n1460), .B1(n1940), .A0N(top_core_KE_key_mem_5__39_), 
        .A1N(n1950), .Y(top_core_KE_n3464) );
  OAI2BB2X1 U25351 ( .B0(n1460), .B1(n1961), .A0N(top_core_KE_key_mem_6__39_), 
        .A1N(n1970), .Y(top_core_KE_n3593) );
  OAI2BB2X1 U25352 ( .B0(n1460), .B1(n1980), .A0N(top_core_KE_key_mem_7__39_), 
        .A1N(n1990), .Y(top_core_KE_n3722) );
  OAI2BB2X1 U25353 ( .B0(n1460), .B1(n2041), .A0N(top_core_KE_key_mem_10__39_), 
        .A1N(n2050), .Y(top_core_KE_n4109) );
  OAI2BB2X1 U25354 ( .B0(n1460), .B1(n2060), .A0N(top_core_KE_key_mem_11__39_), 
        .A1N(n2070), .Y(top_core_KE_n4238) );
  OAI2BB2X1 U25355 ( .B0(n1460), .B1(n2080), .A0N(top_core_KE_key_mem_12__39_), 
        .A1N(n2090), .Y(top_core_KE_n4367) );
  OAI2BB2X1 U25356 ( .B0(n1460), .B1(n2100), .A0N(top_core_KE_key_mem_13__39_), 
        .A1N(n2110), .Y(top_core_KE_n4496) );
  OAI2BB2X1 U25357 ( .B0(n1460), .B1(n2120), .A0N(top_core_KE_key_mem_14__39_), 
        .A1N(n2130), .Y(top_core_KE_n4625) );
  OAI2BB2X1 U25358 ( .B0(n1461), .B1(n1863), .A0N(top_core_KE_key_mem_1__38_), 
        .A1N(n1858), .Y(top_core_KE_n2949) );
  OAI2BB2X1 U25359 ( .B0(n1461), .B1(n1881), .A0N(top_core_KE_key_mem_2__38_), 
        .A1N(n1891), .Y(top_core_KE_n3078) );
  OAI2BB2X1 U25360 ( .B0(n1461), .B1(n1900), .A0N(top_core_KE_key_mem_3__38_), 
        .A1N(n1910), .Y(top_core_KE_n3207) );
  OAI2BB2X1 U25361 ( .B0(n1461), .B1(n1921), .A0N(top_core_KE_key_mem_4__38_), 
        .A1N(n1930), .Y(top_core_KE_n3336) );
  OAI2BB2X1 U25362 ( .B0(n1461), .B1(n1940), .A0N(top_core_KE_key_mem_5__38_), 
        .A1N(n1950), .Y(top_core_KE_n3465) );
  OAI2BB2X1 U25363 ( .B0(n1461), .B1(n1961), .A0N(top_core_KE_key_mem_6__38_), 
        .A1N(n1970), .Y(top_core_KE_n3594) );
  OAI2BB2X1 U25364 ( .B0(n1461), .B1(n1980), .A0N(top_core_KE_key_mem_7__38_), 
        .A1N(n1990), .Y(top_core_KE_n3723) );
  OAI2BB2X1 U25365 ( .B0(n1461), .B1(n2041), .A0N(top_core_KE_key_mem_10__38_), 
        .A1N(n2050), .Y(top_core_KE_n4110) );
  OAI2BB2X1 U25366 ( .B0(n1461), .B1(n2060), .A0N(top_core_KE_key_mem_11__38_), 
        .A1N(n2070), .Y(top_core_KE_n4239) );
  OAI2BB2X1 U25367 ( .B0(n1461), .B1(n2080), .A0N(top_core_KE_key_mem_12__38_), 
        .A1N(n2090), .Y(top_core_KE_n4368) );
  OAI2BB2X1 U25368 ( .B0(n1461), .B1(n2100), .A0N(top_core_KE_key_mem_13__38_), 
        .A1N(n2110), .Y(top_core_KE_n4497) );
  OAI2BB2X1 U25369 ( .B0(n1461), .B1(n2120), .A0N(top_core_KE_key_mem_14__38_), 
        .A1N(n2130), .Y(top_core_KE_n4626) );
  OAI2BB2X1 U25370 ( .B0(n1462), .B1(n1863), .A0N(top_core_KE_key_mem_1__37_), 
        .A1N(n1857), .Y(top_core_KE_n2950) );
  OAI2BB2X1 U25371 ( .B0(n1462), .B1(n1882), .A0N(top_core_KE_key_mem_2__37_), 
        .A1N(n1891), .Y(top_core_KE_n3079) );
  OAI2BB2X1 U25372 ( .B0(n1462), .B1(n1901), .A0N(top_core_KE_key_mem_3__37_), 
        .A1N(n1910), .Y(top_core_KE_n3208) );
  OAI2BB2X1 U25373 ( .B0(n1462), .B1(n1922), .A0N(top_core_KE_key_mem_4__37_), 
        .A1N(n1930), .Y(top_core_KE_n3337) );
  OAI2BB2X1 U25374 ( .B0(n1462), .B1(n1941), .A0N(top_core_KE_key_mem_5__37_), 
        .A1N(n1950), .Y(top_core_KE_n3466) );
  OAI2BB2X1 U25375 ( .B0(n1462), .B1(n1962), .A0N(top_core_KE_key_mem_6__37_), 
        .A1N(n1970), .Y(top_core_KE_n3595) );
  OAI2BB2X1 U25376 ( .B0(n1462), .B1(n1981), .A0N(top_core_KE_key_mem_7__37_), 
        .A1N(n1990), .Y(top_core_KE_n3724) );
  OAI2BB2X1 U25377 ( .B0(n1462), .B1(n2042), .A0N(top_core_KE_key_mem_10__37_), 
        .A1N(n2050), .Y(top_core_KE_n4111) );
  OAI2BB2X1 U25378 ( .B0(n1462), .B1(n2061), .A0N(top_core_KE_key_mem_11__37_), 
        .A1N(n2070), .Y(top_core_KE_n4240) );
  OAI2BB2X1 U25379 ( .B0(n1462), .B1(n2081), .A0N(top_core_KE_key_mem_12__37_), 
        .A1N(n2090), .Y(top_core_KE_n4369) );
  OAI2BB2X1 U25380 ( .B0(n1462), .B1(n2101), .A0N(top_core_KE_key_mem_13__37_), 
        .A1N(n2110), .Y(top_core_KE_n4498) );
  OAI2BB2X1 U25381 ( .B0(n1462), .B1(n2121), .A0N(top_core_KE_key_mem_14__37_), 
        .A1N(n2130), .Y(top_core_KE_n4627) );
  OAI2BB2X1 U25382 ( .B0(n1463), .B1(n1863), .A0N(top_core_KE_key_mem_1__36_), 
        .A1N(n1870), .Y(top_core_KE_n2951) );
  OAI2BB2X1 U25383 ( .B0(n1463), .B1(n1882), .A0N(top_core_KE_key_mem_2__36_), 
        .A1N(n1892), .Y(top_core_KE_n3080) );
  OAI2BB2X1 U25384 ( .B0(n1463), .B1(n1901), .A0N(top_core_KE_key_mem_3__36_), 
        .A1N(n1911), .Y(top_core_KE_n3209) );
  OAI2BB2X1 U25385 ( .B0(n1463), .B1(n1922), .A0N(top_core_KE_key_mem_4__36_), 
        .A1N(n1931), .Y(top_core_KE_n3338) );
  OAI2BB2X1 U25386 ( .B0(n1463), .B1(n1941), .A0N(top_core_KE_key_mem_5__36_), 
        .A1N(n1951), .Y(top_core_KE_n3467) );
  OAI2BB2X1 U25387 ( .B0(n1463), .B1(n1962), .A0N(top_core_KE_key_mem_6__36_), 
        .A1N(n1971), .Y(top_core_KE_n3596) );
  OAI2BB2X1 U25388 ( .B0(n1463), .B1(n1981), .A0N(top_core_KE_key_mem_7__36_), 
        .A1N(n1991), .Y(top_core_KE_n3725) );
  OAI2BB2X1 U25389 ( .B0(n1463), .B1(n2042), .A0N(top_core_KE_key_mem_10__36_), 
        .A1N(n2051), .Y(top_core_KE_n4112) );
  OAI2BB2X1 U25390 ( .B0(n1463), .B1(n2061), .A0N(top_core_KE_key_mem_11__36_), 
        .A1N(n2071), .Y(top_core_KE_n4241) );
  OAI2BB2X1 U25391 ( .B0(n1463), .B1(n2081), .A0N(top_core_KE_key_mem_12__36_), 
        .A1N(n2091), .Y(top_core_KE_n4370) );
  OAI2BB2X1 U25392 ( .B0(n1463), .B1(n2101), .A0N(top_core_KE_key_mem_13__36_), 
        .A1N(n2111), .Y(top_core_KE_n4499) );
  OAI2BB2X1 U25393 ( .B0(n1463), .B1(n2121), .A0N(top_core_KE_key_mem_14__36_), 
        .A1N(n2131), .Y(top_core_KE_n4628) );
  OAI2BB2X1 U25394 ( .B0(n1464), .B1(n1864), .A0N(top_core_KE_key_mem_1__35_), 
        .A1N(n1869), .Y(top_core_KE_n2952) );
  OAI2BB2X1 U25395 ( .B0(n1464), .B1(n1882), .A0N(top_core_KE_key_mem_2__35_), 
        .A1N(n1892), .Y(top_core_KE_n3081) );
  OAI2BB2X1 U25396 ( .B0(n1464), .B1(n1901), .A0N(top_core_KE_key_mem_3__35_), 
        .A1N(n1911), .Y(top_core_KE_n3210) );
  OAI2BB2X1 U25397 ( .B0(n1464), .B1(n1922), .A0N(top_core_KE_key_mem_4__35_), 
        .A1N(n1931), .Y(top_core_KE_n3339) );
  OAI2BB2X1 U25398 ( .B0(n1464), .B1(n1941), .A0N(top_core_KE_key_mem_5__35_), 
        .A1N(n1951), .Y(top_core_KE_n3468) );
  OAI2BB2X1 U25399 ( .B0(n1464), .B1(n1962), .A0N(top_core_KE_key_mem_6__35_), 
        .A1N(n1971), .Y(top_core_KE_n3597) );
  OAI2BB2X1 U25400 ( .B0(n1464), .B1(n1981), .A0N(top_core_KE_key_mem_7__35_), 
        .A1N(n1991), .Y(top_core_KE_n3726) );
  OAI2BB2X1 U25401 ( .B0(n1464), .B1(n2042), .A0N(top_core_KE_key_mem_10__35_), 
        .A1N(n2051), .Y(top_core_KE_n4113) );
  OAI2BB2X1 U25402 ( .B0(n1464), .B1(n2061), .A0N(top_core_KE_key_mem_11__35_), 
        .A1N(n2071), .Y(top_core_KE_n4242) );
  OAI2BB2X1 U25403 ( .B0(n1464), .B1(n2081), .A0N(top_core_KE_key_mem_12__35_), 
        .A1N(n2091), .Y(top_core_KE_n4371) );
  OAI2BB2X1 U25404 ( .B0(n1464), .B1(n2101), .A0N(top_core_KE_key_mem_13__35_), 
        .A1N(n2111), .Y(top_core_KE_n4500) );
  OAI2BB2X1 U25405 ( .B0(n1464), .B1(n2121), .A0N(top_core_KE_key_mem_14__35_), 
        .A1N(n2131), .Y(top_core_KE_n4629) );
  OAI2BB2X1 U25406 ( .B0(n1465), .B1(n1864), .A0N(top_core_KE_key_mem_1__34_), 
        .A1N(n1866), .Y(top_core_KE_n2953) );
  OAI2BB2X1 U25407 ( .B0(n1465), .B1(n1882), .A0N(top_core_KE_key_mem_2__34_), 
        .A1N(n1892), .Y(top_core_KE_n3082) );
  OAI2BB2X1 U25408 ( .B0(n1465), .B1(n1901), .A0N(top_core_KE_key_mem_3__34_), 
        .A1N(n1911), .Y(top_core_KE_n3211) );
  OAI2BB2X1 U25409 ( .B0(n1465), .B1(n1922), .A0N(top_core_KE_key_mem_4__34_), 
        .A1N(n1931), .Y(top_core_KE_n3340) );
  OAI2BB2X1 U25410 ( .B0(n1465), .B1(n1941), .A0N(top_core_KE_key_mem_5__34_), 
        .A1N(n1951), .Y(top_core_KE_n3469) );
  OAI2BB2X1 U25411 ( .B0(n1465), .B1(n1962), .A0N(top_core_KE_key_mem_6__34_), 
        .A1N(n1971), .Y(top_core_KE_n3598) );
  OAI2BB2X1 U25412 ( .B0(n1465), .B1(n1981), .A0N(top_core_KE_key_mem_7__34_), 
        .A1N(n1991), .Y(top_core_KE_n3727) );
  OAI2BB2X1 U25413 ( .B0(n1465), .B1(n2042), .A0N(top_core_KE_key_mem_10__34_), 
        .A1N(n2051), .Y(top_core_KE_n4114) );
  OAI2BB2X1 U25414 ( .B0(n1465), .B1(n2061), .A0N(top_core_KE_key_mem_11__34_), 
        .A1N(n2071), .Y(top_core_KE_n4243) );
  OAI2BB2X1 U25415 ( .B0(n1465), .B1(n2081), .A0N(top_core_KE_key_mem_12__34_), 
        .A1N(n2091), .Y(top_core_KE_n4372) );
  OAI2BB2X1 U25416 ( .B0(n1465), .B1(n2101), .A0N(top_core_KE_key_mem_13__34_), 
        .A1N(n2111), .Y(top_core_KE_n4501) );
  OAI2BB2X1 U25417 ( .B0(n1465), .B1(n2121), .A0N(top_core_KE_key_mem_14__34_), 
        .A1N(n2131), .Y(top_core_KE_n4630) );
  OAI2BB2X1 U25418 ( .B0(n1466), .B1(n1864), .A0N(top_core_KE_key_mem_1__33_), 
        .A1N(n1872), .Y(top_core_KE_n2954) );
  OAI2BB2X1 U25419 ( .B0(n1466), .B1(n1882), .A0N(top_core_KE_key_mem_2__33_), 
        .A1N(n1892), .Y(top_core_KE_n3083) );
  OAI2BB2X1 U25420 ( .B0(n1466), .B1(n1901), .A0N(top_core_KE_key_mem_3__33_), 
        .A1N(n1911), .Y(top_core_KE_n3212) );
  OAI2BB2X1 U25421 ( .B0(n1466), .B1(n1922), .A0N(top_core_KE_key_mem_4__33_), 
        .A1N(n1931), .Y(top_core_KE_n3341) );
  OAI2BB2X1 U25422 ( .B0(n1466), .B1(n1941), .A0N(top_core_KE_key_mem_5__33_), 
        .A1N(n1951), .Y(top_core_KE_n3470) );
  OAI2BB2X1 U25423 ( .B0(n1466), .B1(n1962), .A0N(top_core_KE_key_mem_6__33_), 
        .A1N(n1971), .Y(top_core_KE_n3599) );
  OAI2BB2X1 U25424 ( .B0(n1466), .B1(n1981), .A0N(top_core_KE_key_mem_7__33_), 
        .A1N(n1991), .Y(top_core_KE_n3728) );
  OAI2BB2X1 U25425 ( .B0(n1466), .B1(n2042), .A0N(top_core_KE_key_mem_10__33_), 
        .A1N(n2051), .Y(top_core_KE_n4115) );
  OAI2BB2X1 U25426 ( .B0(n1466), .B1(n2061), .A0N(top_core_KE_key_mem_11__33_), 
        .A1N(n2071), .Y(top_core_KE_n4244) );
  OAI2BB2X1 U25427 ( .B0(n1466), .B1(n2081), .A0N(top_core_KE_key_mem_12__33_), 
        .A1N(n2091), .Y(top_core_KE_n4373) );
  OAI2BB2X1 U25428 ( .B0(n1466), .B1(n2101), .A0N(top_core_KE_key_mem_13__33_), 
        .A1N(n2111), .Y(top_core_KE_n4502) );
  OAI2BB2X1 U25429 ( .B0(n1466), .B1(n2121), .A0N(top_core_KE_key_mem_14__33_), 
        .A1N(n2131), .Y(top_core_KE_n4631) );
  OAI2BB2X1 U25430 ( .B0(n1467), .B1(n1864), .A0N(top_core_KE_key_mem_1__32_), 
        .A1N(n1872), .Y(top_core_KE_n2955) );
  OAI2BB2X1 U25431 ( .B0(n1467), .B1(n1882), .A0N(top_core_KE_key_mem_2__32_), 
        .A1N(n1892), .Y(top_core_KE_n3084) );
  OAI2BB2X1 U25432 ( .B0(n1467), .B1(n1901), .A0N(top_core_KE_key_mem_3__32_), 
        .A1N(n1911), .Y(top_core_KE_n3213) );
  OAI2BB2X1 U25433 ( .B0(n1467), .B1(n1922), .A0N(top_core_KE_key_mem_4__32_), 
        .A1N(n1931), .Y(top_core_KE_n3342) );
  OAI2BB2X1 U25434 ( .B0(n1467), .B1(n1941), .A0N(top_core_KE_key_mem_5__32_), 
        .A1N(n1951), .Y(top_core_KE_n3471) );
  OAI2BB2X1 U25435 ( .B0(n1467), .B1(n1962), .A0N(top_core_KE_key_mem_6__32_), 
        .A1N(n1971), .Y(top_core_KE_n3600) );
  OAI2BB2X1 U25436 ( .B0(n1467), .B1(n1981), .A0N(top_core_KE_key_mem_7__32_), 
        .A1N(n1991), .Y(top_core_KE_n3729) );
  OAI2BB2X1 U25437 ( .B0(n1467), .B1(n2042), .A0N(top_core_KE_key_mem_10__32_), 
        .A1N(n2051), .Y(top_core_KE_n4116) );
  OAI2BB2X1 U25438 ( .B0(n1467), .B1(n2061), .A0N(top_core_KE_key_mem_11__32_), 
        .A1N(n2071), .Y(top_core_KE_n4245) );
  OAI2BB2X1 U25439 ( .B0(n1467), .B1(n2081), .A0N(top_core_KE_key_mem_12__32_), 
        .A1N(n2091), .Y(top_core_KE_n4374) );
  OAI2BB2X1 U25440 ( .B0(n1467), .B1(n2101), .A0N(top_core_KE_key_mem_13__32_), 
        .A1N(n2111), .Y(top_core_KE_n4503) );
  OAI2BB2X1 U25441 ( .B0(n1467), .B1(n2121), .A0N(top_core_KE_key_mem_14__32_), 
        .A1N(n2131), .Y(top_core_KE_n4632) );
  OAI2BB2X1 U25442 ( .B0(n1468), .B1(n1863), .A0N(top_core_KE_key_mem_1__31_), 
        .A1N(n1872), .Y(top_core_KE_n2956) );
  OAI2BB2X1 U25443 ( .B0(n1468), .B1(n1882), .A0N(top_core_KE_key_mem_2__31_), 
        .A1N(n1892), .Y(top_core_KE_n3085) );
  OAI2BB2X1 U25444 ( .B0(n1468), .B1(n1901), .A0N(top_core_KE_key_mem_3__31_), 
        .A1N(n1911), .Y(top_core_KE_n3214) );
  OAI2BB2X1 U25445 ( .B0(n1468), .B1(n1922), .A0N(top_core_KE_key_mem_4__31_), 
        .A1N(n1931), .Y(top_core_KE_n3343) );
  OAI2BB2X1 U25446 ( .B0(n1468), .B1(n1941), .A0N(top_core_KE_key_mem_5__31_), 
        .A1N(n1951), .Y(top_core_KE_n3472) );
  OAI2BB2X1 U25447 ( .B0(n1468), .B1(n1962), .A0N(top_core_KE_key_mem_6__31_), 
        .A1N(n1971), .Y(top_core_KE_n3601) );
  OAI2BB2X1 U25448 ( .B0(n1468), .B1(n1981), .A0N(top_core_KE_key_mem_7__31_), 
        .A1N(n1991), .Y(top_core_KE_n3730) );
  OAI2BB2X1 U25449 ( .B0(n1468), .B1(n2042), .A0N(top_core_KE_key_mem_10__31_), 
        .A1N(n2051), .Y(top_core_KE_n4117) );
  OAI2BB2X1 U25450 ( .B0(n1468), .B1(n2061), .A0N(top_core_KE_key_mem_11__31_), 
        .A1N(n2071), .Y(top_core_KE_n4246) );
  OAI2BB2X1 U25451 ( .B0(n1468), .B1(n2081), .A0N(top_core_KE_key_mem_12__31_), 
        .A1N(n2091), .Y(top_core_KE_n4375) );
  OAI2BB2X1 U25452 ( .B0(n1468), .B1(n2101), .A0N(top_core_KE_key_mem_13__31_), 
        .A1N(n2111), .Y(top_core_KE_n4504) );
  OAI2BB2X1 U25453 ( .B0(n1468), .B1(n2121), .A0N(top_core_KE_key_mem_14__31_), 
        .A1N(n2131), .Y(top_core_KE_n4633) );
  OAI2BB2X1 U25454 ( .B0(n1469), .B1(n1864), .A0N(top_core_KE_key_mem_1__30_), 
        .A1N(n1872), .Y(top_core_KE_n2957) );
  OAI2BB2X1 U25455 ( .B0(n1469), .B1(n1882), .A0N(top_core_KE_key_mem_2__30_), 
        .A1N(n1892), .Y(top_core_KE_n3086) );
  OAI2BB2X1 U25456 ( .B0(n1469), .B1(n1901), .A0N(top_core_KE_key_mem_3__30_), 
        .A1N(n1911), .Y(top_core_KE_n3215) );
  OAI2BB2X1 U25457 ( .B0(n1469), .B1(n1922), .A0N(top_core_KE_key_mem_4__30_), 
        .A1N(n1931), .Y(top_core_KE_n3344) );
  OAI2BB2X1 U25458 ( .B0(n1469), .B1(n1941), .A0N(top_core_KE_key_mem_5__30_), 
        .A1N(n1951), .Y(top_core_KE_n3473) );
  OAI2BB2X1 U25459 ( .B0(n1469), .B1(n1962), .A0N(top_core_KE_key_mem_6__30_), 
        .A1N(n1971), .Y(top_core_KE_n3602) );
  OAI2BB2X1 U25460 ( .B0(n1469), .B1(n1981), .A0N(top_core_KE_key_mem_7__30_), 
        .A1N(n1991), .Y(top_core_KE_n3731) );
  OAI2BB2X1 U25461 ( .B0(n1469), .B1(n2042), .A0N(top_core_KE_key_mem_10__30_), 
        .A1N(n2051), .Y(top_core_KE_n4118) );
  OAI2BB2X1 U25462 ( .B0(n1469), .B1(n2061), .A0N(top_core_KE_key_mem_11__30_), 
        .A1N(n2071), .Y(top_core_KE_n4247) );
  OAI2BB2X1 U25463 ( .B0(n1469), .B1(n2081), .A0N(top_core_KE_key_mem_12__30_), 
        .A1N(n2091), .Y(top_core_KE_n4376) );
  OAI2BB2X1 U25464 ( .B0(n1469), .B1(n2101), .A0N(top_core_KE_key_mem_13__30_), 
        .A1N(n2111), .Y(top_core_KE_n4505) );
  OAI2BB2X1 U25465 ( .B0(n1469), .B1(n2121), .A0N(top_core_KE_key_mem_14__30_), 
        .A1N(n2131), .Y(top_core_KE_n4634) );
  OAI2BB2X1 U25466 ( .B0(n1470), .B1(n1864), .A0N(top_core_KE_key_mem_1__29_), 
        .A1N(n1872), .Y(top_core_KE_n2958) );
  OAI2BB2X1 U25467 ( .B0(n1470), .B1(n1883), .A0N(top_core_KE_key_mem_2__29_), 
        .A1N(n1892), .Y(top_core_KE_n3087) );
  OAI2BB2X1 U25468 ( .B0(n1470), .B1(n1902), .A0N(top_core_KE_key_mem_3__29_), 
        .A1N(n1911), .Y(top_core_KE_n3216) );
  OAI2BB2X1 U25469 ( .B0(n1470), .B1(n1923), .A0N(top_core_KE_key_mem_4__29_), 
        .A1N(n1931), .Y(top_core_KE_n3345) );
  OAI2BB2X1 U25470 ( .B0(n1470), .B1(n1942), .A0N(top_core_KE_key_mem_5__29_), 
        .A1N(n1951), .Y(top_core_KE_n3474) );
  OAI2BB2X1 U25471 ( .B0(n1470), .B1(n1963), .A0N(top_core_KE_key_mem_6__29_), 
        .A1N(n1971), .Y(top_core_KE_n3603) );
  OAI2BB2X1 U25472 ( .B0(n1470), .B1(n1982), .A0N(top_core_KE_key_mem_7__29_), 
        .A1N(n1991), .Y(top_core_KE_n3732) );
  OAI2BB2X1 U25473 ( .B0(n1470), .B1(n2043), .A0N(top_core_KE_key_mem_10__29_), 
        .A1N(n2051), .Y(top_core_KE_n4119) );
  OAI2BB2X1 U25474 ( .B0(n1470), .B1(n2062), .A0N(top_core_KE_key_mem_11__29_), 
        .A1N(n2071), .Y(top_core_KE_n4248) );
  OAI2BB2X1 U25475 ( .B0(n1470), .B1(n2082), .A0N(top_core_KE_key_mem_12__29_), 
        .A1N(n2091), .Y(top_core_KE_n4377) );
  OAI2BB2X1 U25476 ( .B0(n1470), .B1(n2102), .A0N(top_core_KE_key_mem_13__29_), 
        .A1N(n2111), .Y(top_core_KE_n4506) );
  OAI2BB2X1 U25477 ( .B0(n1470), .B1(n2122), .A0N(top_core_KE_key_mem_14__29_), 
        .A1N(n2131), .Y(top_core_KE_n4635) );
  OAI2BB2X1 U25478 ( .B0(n1471), .B1(n1864), .A0N(top_core_KE_key_mem_1__28_), 
        .A1N(n1871), .Y(top_core_KE_n2959) );
  OAI2BB2X1 U25479 ( .B0(n1471), .B1(n1883), .A0N(top_core_KE_key_mem_2__28_), 
        .A1N(n1892), .Y(top_core_KE_n3088) );
  OAI2BB2X1 U25480 ( .B0(n1471), .B1(n1902), .A0N(top_core_KE_key_mem_3__28_), 
        .A1N(n1911), .Y(top_core_KE_n3217) );
  OAI2BB2X1 U25481 ( .B0(n1471), .B1(n1923), .A0N(top_core_KE_key_mem_4__28_), 
        .A1N(n1931), .Y(top_core_KE_n3346) );
  OAI2BB2X1 U25482 ( .B0(n1471), .B1(n1942), .A0N(top_core_KE_key_mem_5__28_), 
        .A1N(n1951), .Y(top_core_KE_n3475) );
  OAI2BB2X1 U25483 ( .B0(n1471), .B1(n1963), .A0N(top_core_KE_key_mem_6__28_), 
        .A1N(n1971), .Y(top_core_KE_n3604) );
  OAI2BB2X1 U25484 ( .B0(n1471), .B1(n1982), .A0N(top_core_KE_key_mem_7__28_), 
        .A1N(n1991), .Y(top_core_KE_n3733) );
  OAI2BB2X1 U25485 ( .B0(n1471), .B1(n2043), .A0N(top_core_KE_key_mem_10__28_), 
        .A1N(n2051), .Y(top_core_KE_n4120) );
  OAI2BB2X1 U25486 ( .B0(n1471), .B1(n2062), .A0N(top_core_KE_key_mem_11__28_), 
        .A1N(n2071), .Y(top_core_KE_n4249) );
  OAI2BB2X1 U25487 ( .B0(n1471), .B1(n2082), .A0N(top_core_KE_key_mem_12__28_), 
        .A1N(n2091), .Y(top_core_KE_n4378) );
  OAI2BB2X1 U25488 ( .B0(n1471), .B1(n2102), .A0N(top_core_KE_key_mem_13__28_), 
        .A1N(n2111), .Y(top_core_KE_n4507) );
  OAI2BB2X1 U25489 ( .B0(n1471), .B1(n2122), .A0N(top_core_KE_key_mem_14__28_), 
        .A1N(n2131), .Y(top_core_KE_n4636) );
  OAI2BB2X1 U25490 ( .B0(n1472), .B1(n1864), .A0N(top_core_KE_key_mem_1__27_), 
        .A1N(n1871), .Y(top_core_KE_n2960) );
  OAI2BB2X1 U25491 ( .B0(n1472), .B1(n1883), .A0N(top_core_KE_key_mem_2__27_), 
        .A1N(n1892), .Y(top_core_KE_n3089) );
  OAI2BB2X1 U25492 ( .B0(n1472), .B1(n1902), .A0N(top_core_KE_key_mem_3__27_), 
        .A1N(n1911), .Y(top_core_KE_n3218) );
  OAI2BB2X1 U25493 ( .B0(n1472), .B1(n1923), .A0N(top_core_KE_key_mem_4__27_), 
        .A1N(n1931), .Y(top_core_KE_n3347) );
  OAI2BB2X1 U25494 ( .B0(n1472), .B1(n1942), .A0N(top_core_KE_key_mem_5__27_), 
        .A1N(n1951), .Y(top_core_KE_n3476) );
  OAI2BB2X1 U25495 ( .B0(n1472), .B1(n1963), .A0N(top_core_KE_key_mem_6__27_), 
        .A1N(n1971), .Y(top_core_KE_n3605) );
  OAI2BB2X1 U25496 ( .B0(n1472), .B1(n1982), .A0N(top_core_KE_key_mem_7__27_), 
        .A1N(n1991), .Y(top_core_KE_n3734) );
  OAI2BB2X1 U25497 ( .B0(n1472), .B1(n2043), .A0N(top_core_KE_key_mem_10__27_), 
        .A1N(n2051), .Y(top_core_KE_n4121) );
  OAI2BB2X1 U25498 ( .B0(n1472), .B1(n2062), .A0N(top_core_KE_key_mem_11__27_), 
        .A1N(n2071), .Y(top_core_KE_n4250) );
  OAI2BB2X1 U25499 ( .B0(n1472), .B1(n2082), .A0N(top_core_KE_key_mem_12__27_), 
        .A1N(n2091), .Y(top_core_KE_n4379) );
  OAI2BB2X1 U25500 ( .B0(n1472), .B1(n2102), .A0N(top_core_KE_key_mem_13__27_), 
        .A1N(n2111), .Y(top_core_KE_n4508) );
  OAI2BB2X1 U25501 ( .B0(n1472), .B1(n2122), .A0N(top_core_KE_key_mem_14__27_), 
        .A1N(n2131), .Y(top_core_KE_n4637) );
  OAI2BB2X1 U25502 ( .B0(n1473), .B1(n1865), .A0N(top_core_KE_key_mem_1__26_), 
        .A1N(n1871), .Y(top_core_KE_n2961) );
  OAI2BB2X1 U25503 ( .B0(n1473), .B1(n1883), .A0N(top_core_KE_key_mem_2__26_), 
        .A1N(n1892), .Y(top_core_KE_n3090) );
  OAI2BB2X1 U25504 ( .B0(n1473), .B1(n1902), .A0N(top_core_KE_key_mem_3__26_), 
        .A1N(n1911), .Y(top_core_KE_n3219) );
  OAI2BB2X1 U25505 ( .B0(n1473), .B1(n1923), .A0N(top_core_KE_key_mem_4__26_), 
        .A1N(n1931), .Y(top_core_KE_n3348) );
  OAI2BB2X1 U25506 ( .B0(n1473), .B1(n1942), .A0N(top_core_KE_key_mem_5__26_), 
        .A1N(n1951), .Y(top_core_KE_n3477) );
  OAI2BB2X1 U25507 ( .B0(n1473), .B1(n1963), .A0N(top_core_KE_key_mem_6__26_), 
        .A1N(n1971), .Y(top_core_KE_n3606) );
  OAI2BB2X1 U25508 ( .B0(n1473), .B1(n1982), .A0N(top_core_KE_key_mem_7__26_), 
        .A1N(n1991), .Y(top_core_KE_n3735) );
  OAI2BB2X1 U25509 ( .B0(n1473), .B1(n2043), .A0N(top_core_KE_key_mem_10__26_), 
        .A1N(n2051), .Y(top_core_KE_n4122) );
  OAI2BB2X1 U25510 ( .B0(n1473), .B1(n2062), .A0N(top_core_KE_key_mem_11__26_), 
        .A1N(n2071), .Y(top_core_KE_n4251) );
  OAI2BB2X1 U25511 ( .B0(n1473), .B1(n2082), .A0N(top_core_KE_key_mem_12__26_), 
        .A1N(n2091), .Y(top_core_KE_n4380) );
  OAI2BB2X1 U25512 ( .B0(n1473), .B1(n2102), .A0N(top_core_KE_key_mem_13__26_), 
        .A1N(n2111), .Y(top_core_KE_n4509) );
  OAI2BB2X1 U25513 ( .B0(n1473), .B1(n2122), .A0N(top_core_KE_key_mem_14__26_), 
        .A1N(n2131), .Y(top_core_KE_n4638) );
  OAI2BB2X1 U25514 ( .B0(n1474), .B1(n1865), .A0N(top_core_KE_key_mem_1__25_), 
        .A1N(n1871), .Y(top_core_KE_n2962) );
  OAI2BB2X1 U25515 ( .B0(n1474), .B1(n1883), .A0N(top_core_KE_key_mem_2__25_), 
        .A1N(n1892), .Y(top_core_KE_n3091) );
  OAI2BB2X1 U25516 ( .B0(n1474), .B1(n1902), .A0N(top_core_KE_key_mem_3__25_), 
        .A1N(n1911), .Y(top_core_KE_n3220) );
  OAI2BB2X1 U25517 ( .B0(n1474), .B1(n1923), .A0N(top_core_KE_key_mem_4__25_), 
        .A1N(n1931), .Y(top_core_KE_n3349) );
  OAI2BB2X1 U25518 ( .B0(n1474), .B1(n1942), .A0N(top_core_KE_key_mem_5__25_), 
        .A1N(n1951), .Y(top_core_KE_n3478) );
  OAI2BB2X1 U25519 ( .B0(n1474), .B1(n1963), .A0N(top_core_KE_key_mem_6__25_), 
        .A1N(n1971), .Y(top_core_KE_n3607) );
  OAI2BB2X1 U25520 ( .B0(n1474), .B1(n1982), .A0N(top_core_KE_key_mem_7__25_), 
        .A1N(n1991), .Y(top_core_KE_n3736) );
  OAI2BB2X1 U25521 ( .B0(n1474), .B1(n2043), .A0N(top_core_KE_key_mem_10__25_), 
        .A1N(n2051), .Y(top_core_KE_n4123) );
  OAI2BB2X1 U25522 ( .B0(n1474), .B1(n2062), .A0N(top_core_KE_key_mem_11__25_), 
        .A1N(n2071), .Y(top_core_KE_n4252) );
  OAI2BB2X1 U25523 ( .B0(n1474), .B1(n2082), .A0N(top_core_KE_key_mem_12__25_), 
        .A1N(n2091), .Y(top_core_KE_n4381) );
  OAI2BB2X1 U25524 ( .B0(n1474), .B1(n2102), .A0N(top_core_KE_key_mem_13__25_), 
        .A1N(n2111), .Y(top_core_KE_n4510) );
  OAI2BB2X1 U25525 ( .B0(n1474), .B1(n2122), .A0N(top_core_KE_key_mem_14__25_), 
        .A1N(n2131), .Y(top_core_KE_n4639) );
  OAI2BB2X1 U25526 ( .B0(n1475), .B1(n1865), .A0N(top_core_KE_key_mem_1__24_), 
        .A1N(n1871), .Y(top_core_KE_n2963) );
  OAI2BB2X1 U25527 ( .B0(n1475), .B1(n1883), .A0N(top_core_KE_key_mem_2__24_), 
        .A1N(n1892), .Y(top_core_KE_n3092) );
  OAI2BB2X1 U25528 ( .B0(n1475), .B1(n1902), .A0N(top_core_KE_key_mem_3__24_), 
        .A1N(n1911), .Y(top_core_KE_n3221) );
  OAI2BB2X1 U25529 ( .B0(n1475), .B1(n1923), .A0N(top_core_KE_key_mem_4__24_), 
        .A1N(n1931), .Y(top_core_KE_n3350) );
  OAI2BB2X1 U25530 ( .B0(n1475), .B1(n1942), .A0N(top_core_KE_key_mem_5__24_), 
        .A1N(n1951), .Y(top_core_KE_n3479) );
  OAI2BB2X1 U25531 ( .B0(n1475), .B1(n1963), .A0N(top_core_KE_key_mem_6__24_), 
        .A1N(n1971), .Y(top_core_KE_n3608) );
  OAI2BB2X1 U25532 ( .B0(n1475), .B1(n1982), .A0N(top_core_KE_key_mem_7__24_), 
        .A1N(n1991), .Y(top_core_KE_n3737) );
  OAI2BB2X1 U25533 ( .B0(n1475), .B1(n2043), .A0N(top_core_KE_key_mem_10__24_), 
        .A1N(n2051), .Y(top_core_KE_n4124) );
  OAI2BB2X1 U25534 ( .B0(n1475), .B1(n2062), .A0N(top_core_KE_key_mem_11__24_), 
        .A1N(n2071), .Y(top_core_KE_n4253) );
  OAI2BB2X1 U25535 ( .B0(n1475), .B1(n2082), .A0N(top_core_KE_key_mem_12__24_), 
        .A1N(n2091), .Y(top_core_KE_n4382) );
  OAI2BB2X1 U25536 ( .B0(n1475), .B1(n2102), .A0N(top_core_KE_key_mem_13__24_), 
        .A1N(n2111), .Y(top_core_KE_n4511) );
  OAI2BB2X1 U25537 ( .B0(n1475), .B1(n2122), .A0N(top_core_KE_key_mem_14__24_), 
        .A1N(n2131), .Y(top_core_KE_n4640) );
  OAI2BB2X1 U25538 ( .B0(n1476), .B1(n1865), .A0N(top_core_KE_key_mem_1__23_), 
        .A1N(n1870), .Y(top_core_KE_n2964) );
  OAI2BB2X1 U25539 ( .B0(n1476), .B1(n1884), .A0N(top_core_KE_key_mem_2__23_), 
        .A1N(n1892), .Y(top_core_KE_n3093) );
  OAI2BB2X1 U25540 ( .B0(n1476), .B1(n1903), .A0N(top_core_KE_key_mem_3__23_), 
        .A1N(n1911), .Y(top_core_KE_n3222) );
  OAI2BB2X1 U25541 ( .B0(n1476), .B1(n1924), .A0N(top_core_KE_key_mem_4__23_), 
        .A1N(n1931), .Y(top_core_KE_n3351) );
  OAI2BB2X1 U25542 ( .B0(n1476), .B1(n1943), .A0N(top_core_KE_key_mem_5__23_), 
        .A1N(n1951), .Y(top_core_KE_n3480) );
  OAI2BB2X1 U25543 ( .B0(n1476), .B1(n1964), .A0N(top_core_KE_key_mem_6__23_), 
        .A1N(n1971), .Y(top_core_KE_n3609) );
  OAI2BB2X1 U25544 ( .B0(n1476), .B1(n1983), .A0N(top_core_KE_key_mem_7__23_), 
        .A1N(n1991), .Y(top_core_KE_n3738) );
  OAI2BB2X1 U25545 ( .B0(n1476), .B1(n2044), .A0N(top_core_KE_key_mem_10__23_), 
        .A1N(n2051), .Y(top_core_KE_n4125) );
  OAI2BB2X1 U25546 ( .B0(n1476), .B1(n2063), .A0N(top_core_KE_key_mem_11__23_), 
        .A1N(n2071), .Y(top_core_KE_n4254) );
  OAI2BB2X1 U25547 ( .B0(n1476), .B1(n2083), .A0N(top_core_KE_key_mem_12__23_), 
        .A1N(n2091), .Y(top_core_KE_n4383) );
  OAI2BB2X1 U25548 ( .B0(n1476), .B1(n2103), .A0N(top_core_KE_key_mem_13__23_), 
        .A1N(n2111), .Y(top_core_KE_n4512) );
  OAI2BB2X1 U25549 ( .B0(n1476), .B1(n2123), .A0N(top_core_KE_key_mem_14__23_), 
        .A1N(n2131), .Y(top_core_KE_n4641) );
  OAI2BB2X1 U25550 ( .B0(n1477), .B1(n1864), .A0N(top_core_KE_key_mem_1__22_), 
        .A1N(n1870), .Y(top_core_KE_n2965) );
  OAI2BB2X1 U25551 ( .B0(n1477), .B1(n1884), .A0N(top_core_KE_key_mem_2__22_), 
        .A1N(n1892), .Y(top_core_KE_n3094) );
  OAI2BB2X1 U25552 ( .B0(n1477), .B1(n1903), .A0N(top_core_KE_key_mem_3__22_), 
        .A1N(n1911), .Y(top_core_KE_n3223) );
  OAI2BB2X1 U25553 ( .B0(n1477), .B1(n1924), .A0N(top_core_KE_key_mem_4__22_), 
        .A1N(n1931), .Y(top_core_KE_n3352) );
  OAI2BB2X1 U25554 ( .B0(n1477), .B1(n1943), .A0N(top_core_KE_key_mem_5__22_), 
        .A1N(n1951), .Y(top_core_KE_n3481) );
  OAI2BB2X1 U25555 ( .B0(n1477), .B1(n1964), .A0N(top_core_KE_key_mem_6__22_), 
        .A1N(n1971), .Y(top_core_KE_n3610) );
  OAI2BB2X1 U25556 ( .B0(n1477), .B1(n1983), .A0N(top_core_KE_key_mem_7__22_), 
        .A1N(n1991), .Y(top_core_KE_n3739) );
  OAI2BB2X1 U25557 ( .B0(n1477), .B1(n2044), .A0N(top_core_KE_key_mem_10__22_), 
        .A1N(n2051), .Y(top_core_KE_n4126) );
  OAI2BB2X1 U25558 ( .B0(n1477), .B1(n2063), .A0N(top_core_KE_key_mem_11__22_), 
        .A1N(n2071), .Y(top_core_KE_n4255) );
  OAI2BB2X1 U25559 ( .B0(n1477), .B1(n2083), .A0N(top_core_KE_key_mem_12__22_), 
        .A1N(n2091), .Y(top_core_KE_n4384) );
  OAI2BB2X1 U25560 ( .B0(n1477), .B1(n2103), .A0N(top_core_KE_key_mem_13__22_), 
        .A1N(n2111), .Y(top_core_KE_n4513) );
  OAI2BB2X1 U25561 ( .B0(n1477), .B1(n2123), .A0N(top_core_KE_key_mem_14__22_), 
        .A1N(n2131), .Y(top_core_KE_n4642) );
  OAI2BB2X1 U25562 ( .B0(n1478), .B1(n1865), .A0N(top_core_KE_key_mem_1__21_), 
        .A1N(n1870), .Y(top_core_KE_n2966) );
  OAI2BB2X1 U25563 ( .B0(n1478), .B1(n1883), .A0N(top_core_KE_key_mem_2__21_), 
        .A1N(n1887), .Y(top_core_KE_n3095) );
  OAI2BB2X1 U25564 ( .B0(n1478), .B1(n1902), .A0N(top_core_KE_key_mem_3__21_), 
        .A1N(n1912), .Y(top_core_KE_n3224) );
  OAI2BB2X1 U25565 ( .B0(n1478), .B1(n1923), .A0N(top_core_KE_key_mem_4__21_), 
        .A1N(n1932), .Y(top_core_KE_n3353) );
  OAI2BB2X1 U25566 ( .B0(n1478), .B1(n1942), .A0N(top_core_KE_key_mem_5__21_), 
        .A1N(n1952), .Y(top_core_KE_n3482) );
  OAI2BB2X1 U25567 ( .B0(n1478), .B1(n1963), .A0N(top_core_KE_key_mem_6__21_), 
        .A1N(n1972), .Y(top_core_KE_n3611) );
  OAI2BB2X1 U25568 ( .B0(n1478), .B1(n1982), .A0N(top_core_KE_key_mem_7__21_), 
        .A1N(n1992), .Y(top_core_KE_n3740) );
  OAI2BB2X1 U25569 ( .B0(n1478), .B1(n2043), .A0N(top_core_KE_key_mem_10__21_), 
        .A1N(n2052), .Y(top_core_KE_n4127) );
  OAI2BB2X1 U25570 ( .B0(n1478), .B1(n2062), .A0N(top_core_KE_key_mem_11__21_), 
        .A1N(n2072), .Y(top_core_KE_n4256) );
  OAI2BB2X1 U25571 ( .B0(n1478), .B1(n2082), .A0N(top_core_KE_key_mem_12__21_), 
        .A1N(n2092), .Y(top_core_KE_n4385) );
  OAI2BB2X1 U25572 ( .B0(n1478), .B1(n2102), .A0N(top_core_KE_key_mem_13__21_), 
        .A1N(n2112), .Y(top_core_KE_n4514) );
  OAI2BB2X1 U25573 ( .B0(n1478), .B1(n2122), .A0N(top_core_KE_key_mem_14__21_), 
        .A1N(n2132), .Y(top_core_KE_n4643) );
  OAI2BB2X1 U25574 ( .B0(n1479), .B1(n1865), .A0N(top_core_KE_key_mem_1__20_), 
        .A1N(n1870), .Y(top_core_KE_n2967) );
  OAI2BB2X1 U25575 ( .B0(n1479), .B1(n1884), .A0N(top_core_KE_key_mem_2__20_), 
        .A1N(n1888), .Y(top_core_KE_n3096) );
  OAI2BB2X1 U25576 ( .B0(n1479), .B1(n1903), .A0N(top_core_KE_key_mem_3__20_), 
        .A1N(n1912), .Y(top_core_KE_n3225) );
  OAI2BB2X1 U25577 ( .B0(n1479), .B1(n1924), .A0N(top_core_KE_key_mem_4__20_), 
        .A1N(n1932), .Y(top_core_KE_n3354) );
  OAI2BB2X1 U25578 ( .B0(n1479), .B1(n1943), .A0N(top_core_KE_key_mem_5__20_), 
        .A1N(n1952), .Y(top_core_KE_n3483) );
  OAI2BB2X1 U25579 ( .B0(n1479), .B1(n1964), .A0N(top_core_KE_key_mem_6__20_), 
        .A1N(n1972), .Y(top_core_KE_n3612) );
  OAI2BB2X1 U25580 ( .B0(n1479), .B1(n1983), .A0N(top_core_KE_key_mem_7__20_), 
        .A1N(n1992), .Y(top_core_KE_n3741) );
  OAI2BB2X1 U25581 ( .B0(n1479), .B1(n2044), .A0N(top_core_KE_key_mem_10__20_), 
        .A1N(n2052), .Y(top_core_KE_n4128) );
  OAI2BB2X1 U25582 ( .B0(n1479), .B1(n2063), .A0N(top_core_KE_key_mem_11__20_), 
        .A1N(n2072), .Y(top_core_KE_n4257) );
  OAI2BB2X1 U25583 ( .B0(n1479), .B1(n2083), .A0N(top_core_KE_key_mem_12__20_), 
        .A1N(n2092), .Y(top_core_KE_n4386) );
  OAI2BB2X1 U25584 ( .B0(n1479), .B1(n2103), .A0N(top_core_KE_key_mem_13__20_), 
        .A1N(n2112), .Y(top_core_KE_n4515) );
  OAI2BB2X1 U25585 ( .B0(n1479), .B1(n2123), .A0N(top_core_KE_key_mem_14__20_), 
        .A1N(n2132), .Y(top_core_KE_n4644) );
  OAI2BB2X1 U25586 ( .B0(n1480), .B1(n1865), .A0N(top_core_KE_key_mem_1__19_), 
        .A1N(n1870), .Y(top_core_KE_n2968) );
  OAI2BB2X1 U25587 ( .B0(n1480), .B1(n1884), .A0N(top_core_KE_key_mem_2__19_), 
        .A1N(n1886), .Y(top_core_KE_n3097) );
  OAI2BB2X1 U25588 ( .B0(n1480), .B1(n1903), .A0N(top_core_KE_key_mem_3__19_), 
        .A1N(n1912), .Y(top_core_KE_n3226) );
  OAI2BB2X1 U25589 ( .B0(n1480), .B1(n1924), .A0N(top_core_KE_key_mem_4__19_), 
        .A1N(n1932), .Y(top_core_KE_n3355) );
  OAI2BB2X1 U25590 ( .B0(n1480), .B1(n1943), .A0N(top_core_KE_key_mem_5__19_), 
        .A1N(n1952), .Y(top_core_KE_n3484) );
  OAI2BB2X1 U25591 ( .B0(n1480), .B1(n1964), .A0N(top_core_KE_key_mem_6__19_), 
        .A1N(n1972), .Y(top_core_KE_n3613) );
  OAI2BB2X1 U25592 ( .B0(n1480), .B1(n1983), .A0N(top_core_KE_key_mem_7__19_), 
        .A1N(n1992), .Y(top_core_KE_n3742) );
  OAI2BB2X1 U25593 ( .B0(n1480), .B1(n2044), .A0N(top_core_KE_key_mem_10__19_), 
        .A1N(n2052), .Y(top_core_KE_n4129) );
  OAI2BB2X1 U25594 ( .B0(n1480), .B1(n2063), .A0N(top_core_KE_key_mem_11__19_), 
        .A1N(n2072), .Y(top_core_KE_n4258) );
  OAI2BB2X1 U25595 ( .B0(n1480), .B1(n2083), .A0N(top_core_KE_key_mem_12__19_), 
        .A1N(n2092), .Y(top_core_KE_n4387) );
  OAI2BB2X1 U25596 ( .B0(n1480), .B1(n2103), .A0N(top_core_KE_key_mem_13__19_), 
        .A1N(n2112), .Y(top_core_KE_n4516) );
  OAI2BB2X1 U25597 ( .B0(n1480), .B1(n2123), .A0N(top_core_KE_key_mem_14__19_), 
        .A1N(n2132), .Y(top_core_KE_n4645) );
  OAI2BB2X1 U25598 ( .B0(n1481), .B1(n1865), .A0N(top_core_KE_key_mem_1__18_), 
        .A1N(n1869), .Y(top_core_KE_n2969) );
  OAI2BB2X1 U25599 ( .B0(n1481), .B1(n1884), .A0N(top_core_KE_key_mem_2__18_), 
        .A1N(n1891), .Y(top_core_KE_n3098) );
  OAI2BB2X1 U25600 ( .B0(n1481), .B1(n1903), .A0N(top_core_KE_key_mem_3__18_), 
        .A1N(n1912), .Y(top_core_KE_n3227) );
  OAI2BB2X1 U25601 ( .B0(n1481), .B1(n1924), .A0N(top_core_KE_key_mem_4__18_), 
        .A1N(n1932), .Y(top_core_KE_n3356) );
  OAI2BB2X1 U25602 ( .B0(n1481), .B1(n1943), .A0N(top_core_KE_key_mem_5__18_), 
        .A1N(n1952), .Y(top_core_KE_n3485) );
  OAI2BB2X1 U25603 ( .B0(n1481), .B1(n1964), .A0N(top_core_KE_key_mem_6__18_), 
        .A1N(n1972), .Y(top_core_KE_n3614) );
  OAI2BB2X1 U25604 ( .B0(n1481), .B1(n1983), .A0N(top_core_KE_key_mem_7__18_), 
        .A1N(n1992), .Y(top_core_KE_n3743) );
  OAI2BB2X1 U25605 ( .B0(n1481), .B1(n2044), .A0N(top_core_KE_key_mem_10__18_), 
        .A1N(n2052), .Y(top_core_KE_n4130) );
  OAI2BB2X1 U25606 ( .B0(n1481), .B1(n2063), .A0N(top_core_KE_key_mem_11__18_), 
        .A1N(n2072), .Y(top_core_KE_n4259) );
  OAI2BB2X1 U25607 ( .B0(n1481), .B1(n2083), .A0N(top_core_KE_key_mem_12__18_), 
        .A1N(n2092), .Y(top_core_KE_n4388) );
  OAI2BB2X1 U25608 ( .B0(n1481), .B1(n2103), .A0N(top_core_KE_key_mem_13__18_), 
        .A1N(n2112), .Y(top_core_KE_n4517) );
  OAI2BB2X1 U25609 ( .B0(n1481), .B1(n2123), .A0N(top_core_KE_key_mem_14__18_), 
        .A1N(n2132), .Y(top_core_KE_n4646) );
  OAI2BB2X1 U25610 ( .B0(n1482), .B1(n1865), .A0N(top_core_KE_key_mem_1__17_), 
        .A1N(n1869), .Y(top_core_KE_n2970) );
  OAI2BB2X1 U25611 ( .B0(n1482), .B1(n1884), .A0N(top_core_KE_key_mem_2__17_), 
        .A1N(n1892), .Y(top_core_KE_n3099) );
  OAI2BB2X1 U25612 ( .B0(n1482), .B1(n1903), .A0N(top_core_KE_key_mem_3__17_), 
        .A1N(n1912), .Y(top_core_KE_n3228) );
  OAI2BB2X1 U25613 ( .B0(n1482), .B1(n1924), .A0N(top_core_KE_key_mem_4__17_), 
        .A1N(n1932), .Y(top_core_KE_n3357) );
  OAI2BB2X1 U25614 ( .B0(n1482), .B1(n1943), .A0N(top_core_KE_key_mem_5__17_), 
        .A1N(n1952), .Y(top_core_KE_n3486) );
  OAI2BB2X1 U25615 ( .B0(n1482), .B1(n1964), .A0N(top_core_KE_key_mem_6__17_), 
        .A1N(n1972), .Y(top_core_KE_n3615) );
  OAI2BB2X1 U25616 ( .B0(n1482), .B1(n1983), .A0N(top_core_KE_key_mem_7__17_), 
        .A1N(n1992), .Y(top_core_KE_n3744) );
  OAI2BB2X1 U25617 ( .B0(n1482), .B1(n2044), .A0N(top_core_KE_key_mem_10__17_), 
        .A1N(n2052), .Y(top_core_KE_n4131) );
  OAI2BB2X1 U25618 ( .B0(n1482), .B1(n2063), .A0N(top_core_KE_key_mem_11__17_), 
        .A1N(n2072), .Y(top_core_KE_n4260) );
  OAI2BB2X1 U25619 ( .B0(n1482), .B1(n2083), .A0N(top_core_KE_key_mem_12__17_), 
        .A1N(n2092), .Y(top_core_KE_n4389) );
  OAI2BB2X1 U25620 ( .B0(n1482), .B1(n2103), .A0N(top_core_KE_key_mem_13__17_), 
        .A1N(n2112), .Y(top_core_KE_n4518) );
  OAI2BB2X1 U25621 ( .B0(n1482), .B1(n2123), .A0N(top_core_KE_key_mem_14__17_), 
        .A1N(n2132), .Y(top_core_KE_n4647) );
  OAI2BB2X1 U25622 ( .B0(n1483), .B1(n1865), .A0N(top_core_KE_key_mem_1__16_), 
        .A1N(n1869), .Y(top_core_KE_n2971) );
  OAI2BB2X1 U25623 ( .B0(n1483), .B1(n1883), .A0N(top_core_KE_key_mem_2__16_), 
        .A1N(n1885), .Y(top_core_KE_n3100) );
  OAI2BB2X1 U25624 ( .B0(n1483), .B1(n1902), .A0N(top_core_KE_key_mem_3__16_), 
        .A1N(n1912), .Y(top_core_KE_n3229) );
  OAI2BB2X1 U25625 ( .B0(n1483), .B1(n1923), .A0N(top_core_KE_key_mem_4__16_), 
        .A1N(n1932), .Y(top_core_KE_n3358) );
  OAI2BB2X1 U25626 ( .B0(n1483), .B1(n1942), .A0N(top_core_KE_key_mem_5__16_), 
        .A1N(n1952), .Y(top_core_KE_n3487) );
  OAI2BB2X1 U25627 ( .B0(n1483), .B1(n1963), .A0N(top_core_KE_key_mem_6__16_), 
        .A1N(n1972), .Y(top_core_KE_n3616) );
  OAI2BB2X1 U25628 ( .B0(n1483), .B1(n1982), .A0N(top_core_KE_key_mem_7__16_), 
        .A1N(n1992), .Y(top_core_KE_n3745) );
  OAI2BB2X1 U25629 ( .B0(n1483), .B1(n2043), .A0N(top_core_KE_key_mem_10__16_), 
        .A1N(n2052), .Y(top_core_KE_n4132) );
  OAI2BB2X1 U25630 ( .B0(n1483), .B1(n2062), .A0N(top_core_KE_key_mem_11__16_), 
        .A1N(n2072), .Y(top_core_KE_n4261) );
  OAI2BB2X1 U25631 ( .B0(n1483), .B1(n2082), .A0N(top_core_KE_key_mem_12__16_), 
        .A1N(n2092), .Y(top_core_KE_n4390) );
  OAI2BB2X1 U25632 ( .B0(n1483), .B1(n2102), .A0N(top_core_KE_key_mem_13__16_), 
        .A1N(n2112), .Y(top_core_KE_n4519) );
  OAI2BB2X1 U25633 ( .B0(n1483), .B1(n2122), .A0N(top_core_KE_key_mem_14__16_), 
        .A1N(n2132), .Y(top_core_KE_n4648) );
  OAI2BB2X1 U25634 ( .B0(n1484), .B1(n1863), .A0N(top_core_KE_key_mem_1__15_), 
        .A1N(n1869), .Y(top_core_KE_n2972) );
  OAI2BB2X1 U25635 ( .B0(n1484), .B1(n1884), .A0N(top_core_KE_key_mem_2__15_), 
        .A1N(n1882), .Y(top_core_KE_n3101) );
  OAI2BB2X1 U25636 ( .B0(n1484), .B1(n1903), .A0N(top_core_KE_key_mem_3__15_), 
        .A1N(n1912), .Y(top_core_KE_n3230) );
  OAI2BB2X1 U25637 ( .B0(n1484), .B1(n1924), .A0N(top_core_KE_key_mem_4__15_), 
        .A1N(n1932), .Y(top_core_KE_n3359) );
  OAI2BB2X1 U25638 ( .B0(n1484), .B1(n1943), .A0N(top_core_KE_key_mem_5__15_), 
        .A1N(n1952), .Y(top_core_KE_n3488) );
  OAI2BB2X1 U25639 ( .B0(n1484), .B1(n1964), .A0N(top_core_KE_key_mem_6__15_), 
        .A1N(n1972), .Y(top_core_KE_n3617) );
  OAI2BB2X1 U25640 ( .B0(n1484), .B1(n1983), .A0N(top_core_KE_key_mem_7__15_), 
        .A1N(n1992), .Y(top_core_KE_n3746) );
  OAI2BB2X1 U25641 ( .B0(n1484), .B1(n2044), .A0N(top_core_KE_key_mem_10__15_), 
        .A1N(n2052), .Y(top_core_KE_n4133) );
  OAI2BB2X1 U25642 ( .B0(n1484), .B1(n2063), .A0N(top_core_KE_key_mem_11__15_), 
        .A1N(n2072), .Y(top_core_KE_n4262) );
  OAI2BB2X1 U25643 ( .B0(n1484), .B1(n2083), .A0N(top_core_KE_key_mem_12__15_), 
        .A1N(n2092), .Y(top_core_KE_n4391) );
  OAI2BB2X1 U25644 ( .B0(n1484), .B1(n2103), .A0N(top_core_KE_key_mem_13__15_), 
        .A1N(n2112), .Y(top_core_KE_n4520) );
  OAI2BB2X1 U25645 ( .B0(n1484), .B1(n2123), .A0N(top_core_KE_key_mem_14__15_), 
        .A1N(n2132), .Y(top_core_KE_n4649) );
  OAI2BB2X1 U25646 ( .B0(n1485), .B1(n1865), .A0N(top_core_KE_key_mem_1__14_), 
        .A1N(n1869), .Y(top_core_KE_n2973) );
  OAI2BB2X1 U25647 ( .B0(n1485), .B1(n1881), .A0N(top_core_KE_key_mem_2__14_), 
        .A1N(n1883), .Y(top_core_KE_n3102) );
  OAI2BB2X1 U25648 ( .B0(n1485), .B1(n1900), .A0N(top_core_KE_key_mem_3__14_), 
        .A1N(n1912), .Y(top_core_KE_n3231) );
  OAI2BB2X1 U25649 ( .B0(n1485), .B1(n1921), .A0N(top_core_KE_key_mem_4__14_), 
        .A1N(n1932), .Y(top_core_KE_n3360) );
  OAI2BB2X1 U25650 ( .B0(n1485), .B1(n1940), .A0N(top_core_KE_key_mem_5__14_), 
        .A1N(n1952), .Y(top_core_KE_n3489) );
  OAI2BB2X1 U25651 ( .B0(n1485), .B1(n1961), .A0N(top_core_KE_key_mem_6__14_), 
        .A1N(n1972), .Y(top_core_KE_n3618) );
  OAI2BB2X1 U25652 ( .B0(n1485), .B1(n1980), .A0N(top_core_KE_key_mem_7__14_), 
        .A1N(n1992), .Y(top_core_KE_n3747) );
  OAI2BB2X1 U25653 ( .B0(n1485), .B1(n2041), .A0N(top_core_KE_key_mem_10__14_), 
        .A1N(n2052), .Y(top_core_KE_n4134) );
  OAI2BB2X1 U25654 ( .B0(n1485), .B1(n2060), .A0N(top_core_KE_key_mem_11__14_), 
        .A1N(n2072), .Y(top_core_KE_n4263) );
  OAI2BB2X1 U25655 ( .B0(n1485), .B1(n2080), .A0N(top_core_KE_key_mem_12__14_), 
        .A1N(n2092), .Y(top_core_KE_n4392) );
  OAI2BB2X1 U25656 ( .B0(n1485), .B1(n2100), .A0N(top_core_KE_key_mem_13__14_), 
        .A1N(n2112), .Y(top_core_KE_n4521) );
  OAI2BB2X1 U25657 ( .B0(n1485), .B1(n2120), .A0N(top_core_KE_key_mem_14__14_), 
        .A1N(n2132), .Y(top_core_KE_n4650) );
  OAI2BB2X1 U25658 ( .B0(n1486), .B1(n1865), .A0N(top_core_KE_key_mem_1__13_), 
        .A1N(n1868), .Y(top_core_KE_n2974) );
  OAI2BB2X1 U25659 ( .B0(n1486), .B1(n1885), .A0N(top_core_KE_key_mem_2__13_), 
        .A1N(n1881), .Y(top_core_KE_n3103) );
  OAI2BB2X1 U25660 ( .B0(n1486), .B1(n1904), .A0N(top_core_KE_key_mem_3__13_), 
        .A1N(n1912), .Y(top_core_KE_n3232) );
  OAI2BB2X1 U25661 ( .B0(n1486), .B1(n1925), .A0N(top_core_KE_key_mem_4__13_), 
        .A1N(n1932), .Y(top_core_KE_n3361) );
  OAI2BB2X1 U25662 ( .B0(n1486), .B1(n1944), .A0N(top_core_KE_key_mem_5__13_), 
        .A1N(n1952), .Y(top_core_KE_n3490) );
  OAI2BB2X1 U25663 ( .B0(n1486), .B1(n1965), .A0N(top_core_KE_key_mem_6__13_), 
        .A1N(n1972), .Y(top_core_KE_n3619) );
  OAI2BB2X1 U25664 ( .B0(n1486), .B1(n1984), .A0N(top_core_KE_key_mem_7__13_), 
        .A1N(n1992), .Y(top_core_KE_n3748) );
  OAI2BB2X1 U25665 ( .B0(n1486), .B1(n2045), .A0N(top_core_KE_key_mem_10__13_), 
        .A1N(n2052), .Y(top_core_KE_n4135) );
  OAI2BB2X1 U25666 ( .B0(n1486), .B1(n2064), .A0N(top_core_KE_key_mem_11__13_), 
        .A1N(n2072), .Y(top_core_KE_n4264) );
  OAI2BB2X1 U25667 ( .B0(n1486), .B1(n2084), .A0N(top_core_KE_key_mem_12__13_), 
        .A1N(n2092), .Y(top_core_KE_n4393) );
  OAI2BB2X1 U25668 ( .B0(n1486), .B1(n2104), .A0N(top_core_KE_key_mem_13__13_), 
        .A1N(n2112), .Y(top_core_KE_n4522) );
  OAI2BB2X1 U25669 ( .B0(n1486), .B1(n2124), .A0N(top_core_KE_key_mem_14__13_), 
        .A1N(n2132), .Y(top_core_KE_n4651) );
  OAI2BB2X1 U25670 ( .B0(n1487), .B1(n1863), .A0N(top_core_KE_key_mem_1__12_), 
        .A1N(n1868), .Y(top_core_KE_n2975) );
  OAI2BB2X1 U25671 ( .B0(n1487), .B1(n1884), .A0N(top_core_KE_key_mem_2__12_), 
        .A1N(n1878), .Y(top_core_KE_n3104) );
  OAI2BB2X1 U25672 ( .B0(n1487), .B1(n1903), .A0N(top_core_KE_key_mem_3__12_), 
        .A1N(n1912), .Y(top_core_KE_n3233) );
  OAI2BB2X1 U25673 ( .B0(n1487), .B1(n1924), .A0N(top_core_KE_key_mem_4__12_), 
        .A1N(n1932), .Y(top_core_KE_n3362) );
  OAI2BB2X1 U25674 ( .B0(n1487), .B1(n1943), .A0N(top_core_KE_key_mem_5__12_), 
        .A1N(n1952), .Y(top_core_KE_n3491) );
  OAI2BB2X1 U25675 ( .B0(n1487), .B1(n1964), .A0N(top_core_KE_key_mem_6__12_), 
        .A1N(n1972), .Y(top_core_KE_n3620) );
  OAI2BB2X1 U25676 ( .B0(n1487), .B1(n1983), .A0N(top_core_KE_key_mem_7__12_), 
        .A1N(n1992), .Y(top_core_KE_n3749) );
  OAI2BB2X1 U25677 ( .B0(n1487), .B1(n2044), .A0N(top_core_KE_key_mem_10__12_), 
        .A1N(n2052), .Y(top_core_KE_n4136) );
  OAI2BB2X1 U25678 ( .B0(n1487), .B1(n2063), .A0N(top_core_KE_key_mem_11__12_), 
        .A1N(n2072), .Y(top_core_KE_n4265) );
  OAI2BB2X1 U25679 ( .B0(n1487), .B1(n2083), .A0N(top_core_KE_key_mem_12__12_), 
        .A1N(n2092), .Y(top_core_KE_n4394) );
  OAI2BB2X1 U25680 ( .B0(n1487), .B1(n2103), .A0N(top_core_KE_key_mem_13__12_), 
        .A1N(n2112), .Y(top_core_KE_n4523) );
  OAI2BB2X1 U25681 ( .B0(n1487), .B1(n2123), .A0N(top_core_KE_key_mem_14__12_), 
        .A1N(n2132), .Y(top_core_KE_n4652) );
  OAI2BB2X1 U25682 ( .B0(n1488), .B1(n1865), .A0N(top_core_KE_key_mem_1__11_), 
        .A1N(n1868), .Y(top_core_KE_n2976) );
  OAI2BB2X1 U25683 ( .B0(n1488), .B1(n1880), .A0N(top_core_KE_key_mem_2__11_), 
        .A1N(n1880), .Y(top_core_KE_n3105) );
  OAI2BB2X1 U25684 ( .B0(n1488), .B1(n1899), .A0N(top_core_KE_key_mem_3__11_), 
        .A1N(n1912), .Y(top_core_KE_n3234) );
  OAI2BB2X1 U25685 ( .B0(n1488), .B1(n1920), .A0N(top_core_KE_key_mem_4__11_), 
        .A1N(n1932), .Y(top_core_KE_n3363) );
  OAI2BB2X1 U25686 ( .B0(n1488), .B1(n1939), .A0N(top_core_KE_key_mem_5__11_), 
        .A1N(n1952), .Y(top_core_KE_n3492) );
  OAI2BB2X1 U25687 ( .B0(n1488), .B1(n1960), .A0N(top_core_KE_key_mem_6__11_), 
        .A1N(n1972), .Y(top_core_KE_n3621) );
  OAI2BB2X1 U25688 ( .B0(n1488), .B1(n1979), .A0N(top_core_KE_key_mem_7__11_), 
        .A1N(n1992), .Y(top_core_KE_n3750) );
  OAI2BB2X1 U25689 ( .B0(n1488), .B1(n2040), .A0N(top_core_KE_key_mem_10__11_), 
        .A1N(n2052), .Y(top_core_KE_n4137) );
  OAI2BB2X1 U25690 ( .B0(n1488), .B1(n2059), .A0N(top_core_KE_key_mem_11__11_), 
        .A1N(n2072), .Y(top_core_KE_n4266) );
  OAI2BB2X1 U25691 ( .B0(n1488), .B1(n2079), .A0N(top_core_KE_key_mem_12__11_), 
        .A1N(n2092), .Y(top_core_KE_n4395) );
  OAI2BB2X1 U25692 ( .B0(n1488), .B1(n2099), .A0N(top_core_KE_key_mem_13__11_), 
        .A1N(n2112), .Y(top_core_KE_n4524) );
  OAI2BB2X1 U25693 ( .B0(n1488), .B1(n2119), .A0N(top_core_KE_key_mem_14__11_), 
        .A1N(n2132), .Y(top_core_KE_n4653) );
  OAI2BB2X1 U25694 ( .B0(n1489), .B1(n1864), .A0N(top_core_KE_key_mem_1__10_), 
        .A1N(n1869), .Y(top_core_KE_n2977) );
  OAI2BB2X1 U25695 ( .B0(n1489), .B1(n1878), .A0N(top_core_KE_key_mem_2__10_), 
        .A1N(n1879), .Y(top_core_KE_n3106) );
  OAI2BB2X1 U25696 ( .B0(n1489), .B1(n1898), .A0N(top_core_KE_key_mem_3__10_), 
        .A1N(n1912), .Y(top_core_KE_n3235) );
  OAI2BB2X1 U25697 ( .B0(n1489), .B1(n1918), .A0N(top_core_KE_key_mem_4__10_), 
        .A1N(n1932), .Y(top_core_KE_n3364) );
  OAI2BB2X1 U25698 ( .B0(n1489), .B1(n1937), .A0N(top_core_KE_key_mem_5__10_), 
        .A1N(n1952), .Y(top_core_KE_n3493) );
  OAI2BB2X1 U25699 ( .B0(n1489), .B1(n1958), .A0N(top_core_KE_key_mem_6__10_), 
        .A1N(n1972), .Y(top_core_KE_n3622) );
  OAI2BB2X1 U25700 ( .B0(n1489), .B1(n1977), .A0N(top_core_KE_key_mem_7__10_), 
        .A1N(n1992), .Y(top_core_KE_n3751) );
  OAI2BB2X1 U25701 ( .B0(n1489), .B1(n2038), .A0N(top_core_KE_key_mem_10__10_), 
        .A1N(n2052), .Y(top_core_KE_n4138) );
  OAI2BB2X1 U25702 ( .B0(n1489), .B1(n2057), .A0N(top_core_KE_key_mem_11__10_), 
        .A1N(n2072), .Y(top_core_KE_n4267) );
  OAI2BB2X1 U25703 ( .B0(n1489), .B1(n2077), .A0N(top_core_KE_key_mem_12__10_), 
        .A1N(n2092), .Y(top_core_KE_n4396) );
  OAI2BB2X1 U25704 ( .B0(n1489), .B1(n2097), .A0N(top_core_KE_key_mem_13__10_), 
        .A1N(n2112), .Y(top_core_KE_n4525) );
  OAI2BB2X1 U25705 ( .B0(n1489), .B1(n2117), .A0N(top_core_KE_key_mem_14__10_), 
        .A1N(n2132), .Y(top_core_KE_n4654) );
  OAI2BB2X1 U25706 ( .B0(n1490), .B1(n1862), .A0N(top_core_KE_key_mem_1__9_), 
        .A1N(n1867), .Y(top_core_KE_n2978) );
  OAI2BB2X1 U25707 ( .B0(n1490), .B1(n1879), .A0N(top_core_KE_key_mem_2__9_), 
        .A1N(n1877), .Y(top_core_KE_n3107) );
  OAI2BB2X1 U25708 ( .B0(n1490), .B1(n1900), .A0N(top_core_KE_key_mem_3__9_), 
        .A1N(n1912), .Y(top_core_KE_n3236) );
  OAI2BB2X1 U25709 ( .B0(n1490), .B1(n1919), .A0N(top_core_KE_key_mem_4__9_), 
        .A1N(n1932), .Y(top_core_KE_n3365) );
  OAI2BB2X1 U25710 ( .B0(n1490), .B1(n1938), .A0N(top_core_KE_key_mem_5__9_), 
        .A1N(n1952), .Y(top_core_KE_n3494) );
  OAI2BB2X1 U25711 ( .B0(n1490), .B1(n1959), .A0N(top_core_KE_key_mem_6__9_), 
        .A1N(n1972), .Y(top_core_KE_n3623) );
  OAI2BB2X1 U25712 ( .B0(n1490), .B1(n1978), .A0N(top_core_KE_key_mem_7__9_), 
        .A1N(n1992), .Y(top_core_KE_n3752) );
  OAI2BB2X1 U25713 ( .B0(n1490), .B1(n2039), .A0N(top_core_KE_key_mem_10__9_), 
        .A1N(n2052), .Y(top_core_KE_n4139) );
  OAI2BB2X1 U25714 ( .B0(n1490), .B1(n2058), .A0N(top_core_KE_key_mem_11__9_), 
        .A1N(n2072), .Y(top_core_KE_n4268) );
  OAI2BB2X1 U25715 ( .B0(n1490), .B1(n2078), .A0N(top_core_KE_key_mem_12__9_), 
        .A1N(n2092), .Y(top_core_KE_n4397) );
  OAI2BB2X1 U25716 ( .B0(n1490), .B1(n2098), .A0N(top_core_KE_key_mem_13__9_), 
        .A1N(n2112), .Y(top_core_KE_n4526) );
  OAI2BB2X1 U25717 ( .B0(n1490), .B1(n2118), .A0N(top_core_KE_key_mem_14__9_), 
        .A1N(n2132), .Y(top_core_KE_n4655) );
  OAI2BB2X1 U25718 ( .B0(n1491), .B1(n1864), .A0N(top_core_KE_key_mem_1__8_), 
        .A1N(n1867), .Y(top_core_KE_n2979) );
  OAI2BB2X1 U25719 ( .B0(n1491), .B1(n1885), .A0N(top_core_KE_key_mem_2__8_), 
        .A1N(n1884), .Y(top_core_KE_n3108) );
  OAI2BB2X1 U25720 ( .B0(n1491), .B1(n1904), .A0N(top_core_KE_key_mem_3__8_), 
        .A1N(n1912), .Y(top_core_KE_n3237) );
  OAI2BB2X1 U25721 ( .B0(n1491), .B1(n1925), .A0N(top_core_KE_key_mem_4__8_), 
        .A1N(n1932), .Y(top_core_KE_n3366) );
  OAI2BB2X1 U25722 ( .B0(n1491), .B1(n1944), .A0N(top_core_KE_key_mem_5__8_), 
        .A1N(n1952), .Y(top_core_KE_n3495) );
  OAI2BB2X1 U25723 ( .B0(n1491), .B1(n1965), .A0N(top_core_KE_key_mem_6__8_), 
        .A1N(n1972), .Y(top_core_KE_n3624) );
  OAI2BB2X1 U25724 ( .B0(n1491), .B1(n1984), .A0N(top_core_KE_key_mem_7__8_), 
        .A1N(n1992), .Y(top_core_KE_n3753) );
  OAI2BB2X1 U25725 ( .B0(n1491), .B1(n2045), .A0N(top_core_KE_key_mem_10__8_), 
        .A1N(n2052), .Y(top_core_KE_n4140) );
  OAI2BB2X1 U25726 ( .B0(n1491), .B1(n2064), .A0N(top_core_KE_key_mem_11__8_), 
        .A1N(n2072), .Y(top_core_KE_n4269) );
  OAI2BB2X1 U25727 ( .B0(n1491), .B1(n2084), .A0N(top_core_KE_key_mem_12__8_), 
        .A1N(n2092), .Y(top_core_KE_n4398) );
  OAI2BB2X1 U25728 ( .B0(n1491), .B1(n2104), .A0N(top_core_KE_key_mem_13__8_), 
        .A1N(n2112), .Y(top_core_KE_n4527) );
  OAI2BB2X1 U25729 ( .B0(n1491), .B1(n2124), .A0N(top_core_KE_key_mem_14__8_), 
        .A1N(n2132), .Y(top_core_KE_n4656) );
  OAI2BB2X1 U25730 ( .B0(n1492), .B1(n1864), .A0N(top_core_KE_key_mem_1__7_), 
        .A1N(n1867), .Y(top_core_KE_n2980) );
  OAI2BB2X1 U25731 ( .B0(n1492), .B1(n1884), .A0N(top_core_KE_key_mem_2__7_), 
        .A1N(n1889), .Y(top_core_KE_n3109) );
  OAI2BB2X1 U25732 ( .B0(n1492), .B1(n1903), .A0N(top_core_KE_key_mem_3__7_), 
        .A1N(n1912), .Y(top_core_KE_n3238) );
  OAI2BB2X1 U25733 ( .B0(n1492), .B1(n1924), .A0N(top_core_KE_key_mem_4__7_), 
        .A1N(n1932), .Y(top_core_KE_n3367) );
  OAI2BB2X1 U25734 ( .B0(n1492), .B1(n1943), .A0N(top_core_KE_key_mem_5__7_), 
        .A1N(n1952), .Y(top_core_KE_n3496) );
  OAI2BB2X1 U25735 ( .B0(n1492), .B1(n1964), .A0N(top_core_KE_key_mem_6__7_), 
        .A1N(n1972), .Y(top_core_KE_n3625) );
  OAI2BB2X1 U25736 ( .B0(n1492), .B1(n1983), .A0N(top_core_KE_key_mem_7__7_), 
        .A1N(n1992), .Y(top_core_KE_n3754) );
  OAI2BB2X1 U25737 ( .B0(n1492), .B1(n2044), .A0N(top_core_KE_key_mem_10__7_), 
        .A1N(n2052), .Y(top_core_KE_n4141) );
  OAI2BB2X1 U25738 ( .B0(n1492), .B1(n2063), .A0N(top_core_KE_key_mem_11__7_), 
        .A1N(n2072), .Y(top_core_KE_n4270) );
  OAI2BB2X1 U25739 ( .B0(n1492), .B1(n2083), .A0N(top_core_KE_key_mem_12__7_), 
        .A1N(n2092), .Y(top_core_KE_n4399) );
  OAI2BB2X1 U25740 ( .B0(n1492), .B1(n2103), .A0N(top_core_KE_key_mem_13__7_), 
        .A1N(n2112), .Y(top_core_KE_n4528) );
  OAI2BB2X1 U25741 ( .B0(n1492), .B1(n2123), .A0N(top_core_KE_key_mem_14__7_), 
        .A1N(n2132), .Y(top_core_KE_n4657) );
  OAI2BB2X1 U25742 ( .B0(n1493), .B1(n1863), .A0N(top_core_KE_key_mem_1__6_), 
        .A1N(n1867), .Y(top_core_KE_n2981) );
  OAI2BB2X1 U25743 ( .B0(n1493), .B1(n1877), .A0N(top_core_KE_key_mem_2__6_), 
        .A1N(n1881), .Y(top_core_KE_n3110) );
  OAI2BB2X1 U25744 ( .B0(n1493), .B1(n1897), .A0N(top_core_KE_key_mem_3__6_), 
        .A1N(n1900), .Y(top_core_KE_n3239) );
  OAI2BB2X1 U25745 ( .B0(n1493), .B1(n1917), .A0N(top_core_KE_key_mem_4__6_), 
        .A1N(n1921), .Y(top_core_KE_n3368) );
  OAI2BB2X1 U25746 ( .B0(n1493), .B1(n1937), .A0N(top_core_KE_key_mem_5__6_), 
        .A1N(n1940), .Y(top_core_KE_n3497) );
  OAI2BB2X1 U25747 ( .B0(n1493), .B1(n1957), .A0N(top_core_KE_key_mem_6__6_), 
        .A1N(n1961), .Y(top_core_KE_n3626) );
  OAI2BB2X1 U25748 ( .B0(n1493), .B1(n1983), .A0N(top_core_KE_key_mem_7__6_), 
        .A1N(n1980), .Y(top_core_KE_n3755) );
  OAI2BB2X1 U25749 ( .B0(n1493), .B1(n2037), .A0N(top_core_KE_key_mem_10__6_), 
        .A1N(n2041), .Y(top_core_KE_n4142) );
  OAI2BB2X1 U25750 ( .B0(n1493), .B1(n2063), .A0N(top_core_KE_key_mem_11__6_), 
        .A1N(n2060), .Y(top_core_KE_n4271) );
  OAI2BB2X1 U25751 ( .B0(n1493), .B1(n2077), .A0N(top_core_KE_key_mem_12__6_), 
        .A1N(n2080), .Y(top_core_KE_n4400) );
  OAI2BB2X1 U25752 ( .B0(n1493), .B1(n2103), .A0N(top_core_KE_key_mem_13__6_), 
        .A1N(n2100), .Y(top_core_KE_n4529) );
  OAI2BB2X1 U25753 ( .B0(n1493), .B1(n2123), .A0N(top_core_KE_key_mem_14__6_), 
        .A1N(n2120), .Y(top_core_KE_n4658) );
  OAI2BB2X1 U25754 ( .B0(n1494), .B1(n1864), .A0N(top_core_KE_key_mem_1__5_), 
        .A1N(n1867), .Y(top_core_KE_n2982) );
  OAI2BB2X1 U25755 ( .B0(n1494), .B1(n1885), .A0N(top_core_KE_key_mem_2__5_), 
        .A1N(n1882), .Y(top_core_KE_n3111) );
  OAI2BB2X1 U25756 ( .B0(n1494), .B1(n1904), .A0N(top_core_KE_key_mem_3__5_), 
        .A1N(n1901), .Y(top_core_KE_n3240) );
  OAI2BB2X1 U25757 ( .B0(n1494), .B1(n1925), .A0N(top_core_KE_key_mem_4__5_), 
        .A1N(n1922), .Y(top_core_KE_n3369) );
  OAI2BB2X1 U25758 ( .B0(n1494), .B1(n1944), .A0N(top_core_KE_key_mem_5__5_), 
        .A1N(n1941), .Y(top_core_KE_n3498) );
  OAI2BB2X1 U25759 ( .B0(n1494), .B1(n1965), .A0N(top_core_KE_key_mem_6__5_), 
        .A1N(n1962), .Y(top_core_KE_n3627) );
  OAI2BB2X1 U25760 ( .B0(n1494), .B1(n1984), .A0N(top_core_KE_key_mem_7__5_), 
        .A1N(n1981), .Y(top_core_KE_n3756) );
  OAI2BB2X1 U25761 ( .B0(n1494), .B1(n2045), .A0N(top_core_KE_key_mem_10__5_), 
        .A1N(n2042), .Y(top_core_KE_n4143) );
  OAI2BB2X1 U25762 ( .B0(n1494), .B1(n2064), .A0N(top_core_KE_key_mem_11__5_), 
        .A1N(n2061), .Y(top_core_KE_n4272) );
  OAI2BB2X1 U25763 ( .B0(n1494), .B1(n2084), .A0N(top_core_KE_key_mem_12__5_), 
        .A1N(n2081), .Y(top_core_KE_n4401) );
  OAI2BB2X1 U25764 ( .B0(n1494), .B1(n2104), .A0N(top_core_KE_key_mem_13__5_), 
        .A1N(n2101), .Y(top_core_KE_n4530) );
  OAI2BB2X1 U25765 ( .B0(n1494), .B1(n2124), .A0N(top_core_KE_key_mem_14__5_), 
        .A1N(n2121), .Y(top_core_KE_n4659) );
  OAI2BB2X1 U25766 ( .B0(n1495), .B1(n1863), .A0N(top_core_KE_key_mem_1__4_), 
        .A1N(n1866), .Y(top_core_KE_n2983) );
  OAI2BB2X1 U25767 ( .B0(n1495), .B1(n1885), .A0N(top_core_KE_key_mem_2__4_), 
        .A1N(n1883), .Y(top_core_KE_n3112) );
  OAI2BB2X1 U25768 ( .B0(n1495), .B1(n1904), .A0N(top_core_KE_key_mem_3__4_), 
        .A1N(n1902), .Y(top_core_KE_n3241) );
  OAI2BB2X1 U25769 ( .B0(n1495), .B1(n1925), .A0N(top_core_KE_key_mem_4__4_), 
        .A1N(n1923), .Y(top_core_KE_n3370) );
  OAI2BB2X1 U25770 ( .B0(n1495), .B1(n1944), .A0N(top_core_KE_key_mem_5__4_), 
        .A1N(n1942), .Y(top_core_KE_n3499) );
  OAI2BB2X1 U25771 ( .B0(n1495), .B1(n1965), .A0N(top_core_KE_key_mem_6__4_), 
        .A1N(n1963), .Y(top_core_KE_n3628) );
  OAI2BB2X1 U25772 ( .B0(n1495), .B1(n1984), .A0N(top_core_KE_key_mem_7__4_), 
        .A1N(n1982), .Y(top_core_KE_n3757) );
  OAI2BB2X1 U25773 ( .B0(n1495), .B1(n2045), .A0N(top_core_KE_key_mem_10__4_), 
        .A1N(n2043), .Y(top_core_KE_n4144) );
  OAI2BB2X1 U25774 ( .B0(n1495), .B1(n2064), .A0N(top_core_KE_key_mem_11__4_), 
        .A1N(n2062), .Y(top_core_KE_n4273) );
  OAI2BB2X1 U25775 ( .B0(n1495), .B1(n2084), .A0N(top_core_KE_key_mem_12__4_), 
        .A1N(n2082), .Y(top_core_KE_n4402) );
  OAI2BB2X1 U25776 ( .B0(n1495), .B1(n2104), .A0N(top_core_KE_key_mem_13__4_), 
        .A1N(n2102), .Y(top_core_KE_n4531) );
  OAI2BB2X1 U25777 ( .B0(n1495), .B1(n2124), .A0N(top_core_KE_key_mem_14__4_), 
        .A1N(n2122), .Y(top_core_KE_n4660) );
  OAI2BB2X1 U25778 ( .B0(n1496), .B1(n1863), .A0N(top_core_KE_key_mem_1__3_), 
        .A1N(n1866), .Y(top_core_KE_n2984) );
  OAI2BB2X1 U25779 ( .B0(n1496), .B1(n1885), .A0N(top_core_KE_key_mem_2__3_), 
        .A1N(n1889), .Y(top_core_KE_n3113) );
  OAI2BB2X1 U25780 ( .B0(n1496), .B1(n1904), .A0N(top_core_KE_key_mem_3__3_), 
        .A1N(n1908), .Y(top_core_KE_n3242) );
  OAI2BB2X1 U25781 ( .B0(n1496), .B1(n1925), .A0N(top_core_KE_key_mem_4__3_), 
        .A1N(n1929), .Y(top_core_KE_n3371) );
  OAI2BB2X1 U25782 ( .B0(n1496), .B1(n1944), .A0N(top_core_KE_key_mem_5__3_), 
        .A1N(n1948), .Y(top_core_KE_n3500) );
  OAI2BB2X1 U25783 ( .B0(n1496), .B1(n1965), .A0N(top_core_KE_key_mem_6__3_), 
        .A1N(n1968), .Y(top_core_KE_n3629) );
  OAI2BB2X1 U25784 ( .B0(n1496), .B1(n1984), .A0N(top_core_KE_key_mem_7__3_), 
        .A1N(n1988), .Y(top_core_KE_n3758) );
  OAI2BB2X1 U25785 ( .B0(n1496), .B1(n2045), .A0N(top_core_KE_key_mem_10__3_), 
        .A1N(n2052), .Y(top_core_KE_n4145) );
  OAI2BB2X1 U25786 ( .B0(n1496), .B1(n2064), .A0N(top_core_KE_key_mem_11__3_), 
        .A1N(n2068), .Y(top_core_KE_n4274) );
  OAI2BB2X1 U25787 ( .B0(n1496), .B1(n2084), .A0N(top_core_KE_key_mem_12__3_), 
        .A1N(n2088), .Y(top_core_KE_n4403) );
  OAI2BB2X1 U25788 ( .B0(n1496), .B1(n2104), .A0N(top_core_KE_key_mem_13__3_), 
        .A1N(n2108), .Y(top_core_KE_n4532) );
  OAI2BB2X1 U25789 ( .B0(n1496), .B1(n2124), .A0N(top_core_KE_key_mem_14__3_), 
        .A1N(n2128), .Y(top_core_KE_n4661) );
  OAI2BB2X1 U25790 ( .B0(n1497), .B1(n1863), .A0N(top_core_KE_key_mem_1__2_), 
        .A1N(n1867), .Y(top_core_KE_n2985) );
  OAI2BB2X1 U25791 ( .B0(n1497), .B1(n1885), .A0N(top_core_KE_key_mem_2__2_), 
        .A1N(n1890), .Y(top_core_KE_n3114) );
  OAI2BB2X1 U25792 ( .B0(n1497), .B1(n1904), .A0N(top_core_KE_key_mem_3__2_), 
        .A1N(n1909), .Y(top_core_KE_n3243) );
  OAI2BB2X1 U25793 ( .B0(n1497), .B1(n1925), .A0N(top_core_KE_key_mem_4__2_), 
        .A1N(n1932), .Y(top_core_KE_n3372) );
  OAI2BB2X1 U25794 ( .B0(n1497), .B1(n1944), .A0N(top_core_KE_key_mem_5__2_), 
        .A1N(n1949), .Y(top_core_KE_n3501) );
  OAI2BB2X1 U25795 ( .B0(n1497), .B1(n1965), .A0N(top_core_KE_key_mem_6__2_), 
        .A1N(n1969), .Y(top_core_KE_n3630) );
  OAI2BB2X1 U25796 ( .B0(n1497), .B1(n1984), .A0N(top_core_KE_key_mem_7__2_), 
        .A1N(n1989), .Y(top_core_KE_n3759) );
  OAI2BB2X1 U25797 ( .B0(n1497), .B1(n2045), .A0N(top_core_KE_key_mem_10__2_), 
        .A1N(n2049), .Y(top_core_KE_n4146) );
  OAI2BB2X1 U25798 ( .B0(n1497), .B1(n2064), .A0N(top_core_KE_key_mem_11__2_), 
        .A1N(n2069), .Y(top_core_KE_n4275) );
  OAI2BB2X1 U25799 ( .B0(n1497), .B1(n2084), .A0N(top_core_KE_key_mem_12__2_), 
        .A1N(n2089), .Y(top_core_KE_n4404) );
  OAI2BB2X1 U25800 ( .B0(n1497), .B1(n2104), .A0N(top_core_KE_key_mem_13__2_), 
        .A1N(n2109), .Y(top_core_KE_n4533) );
  OAI2BB2X1 U25801 ( .B0(n1497), .B1(n2124), .A0N(top_core_KE_key_mem_14__2_), 
        .A1N(n2129), .Y(top_core_KE_n4662) );
  OAI2BB2X1 U25802 ( .B0(n1498), .B1(n1863), .A0N(top_core_KE_key_mem_1__1_), 
        .A1N(n1866), .Y(top_core_KE_n2986) );
  OAI2BB2X1 U25803 ( .B0(n1498), .B1(n1885), .A0N(top_core_KE_key_mem_2__1_), 
        .A1N(n1888), .Y(top_core_KE_n3115) );
  OAI2BB2X1 U25804 ( .B0(n1498), .B1(n1904), .A0N(top_core_KE_key_mem_3__1_), 
        .A1N(n1907), .Y(top_core_KE_n3244) );
  OAI2BB2X1 U25805 ( .B0(n1498), .B1(n1925), .A0N(top_core_KE_key_mem_4__1_), 
        .A1N(n1928), .Y(top_core_KE_n3373) );
  OAI2BB2X1 U25806 ( .B0(n1498), .B1(n1944), .A0N(top_core_KE_key_mem_5__1_), 
        .A1N(n1947), .Y(top_core_KE_n3502) );
  OAI2BB2X1 U25807 ( .B0(n1498), .B1(n1965), .A0N(top_core_KE_key_mem_6__1_), 
        .A1N(n1957), .Y(top_core_KE_n3631) );
  OAI2BB2X1 U25808 ( .B0(n1498), .B1(n1984), .A0N(top_core_KE_key_mem_7__1_), 
        .A1N(n1987), .Y(top_core_KE_n3760) );
  OAI2BB2X1 U25809 ( .B0(n1498), .B1(n2045), .A0N(top_core_KE_key_mem_10__1_), 
        .A1N(n2048), .Y(top_core_KE_n4147) );
  OAI2BB2X1 U25810 ( .B0(n1498), .B1(n2064), .A0N(top_core_KE_key_mem_11__1_), 
        .A1N(n2067), .Y(top_core_KE_n4276) );
  OAI2BB2X1 U25811 ( .B0(n1498), .B1(n2084), .A0N(top_core_KE_key_mem_12__1_), 
        .A1N(n2087), .Y(top_core_KE_n4405) );
  OAI2BB2X1 U25812 ( .B0(n1498), .B1(n2104), .A0N(top_core_KE_key_mem_13__1_), 
        .A1N(n2107), .Y(top_core_KE_n4534) );
  OAI2BB2X1 U25813 ( .B0(n1498), .B1(n2124), .A0N(top_core_KE_key_mem_14__1_), 
        .A1N(n2127), .Y(top_core_KE_n4663) );
  OAI2BB2X1 U25814 ( .B0(n1499), .B1(n1862), .A0N(top_core_KE_key_mem_1__0_), 
        .A1N(n1866), .Y(top_core_KE_n2987) );
  OAI2BB2X1 U25815 ( .B0(n1499), .B1(n1884), .A0N(top_core_KE_key_mem_2__0_), 
        .A1N(n1888), .Y(top_core_KE_n3116) );
  OAI2BB2X1 U25816 ( .B0(n1499), .B1(n1903), .A0N(top_core_KE_key_mem_3__0_), 
        .A1N(n1907), .Y(top_core_KE_n3245) );
  OAI2BB2X1 U25817 ( .B0(n1499), .B1(n1924), .A0N(top_core_KE_key_mem_4__0_), 
        .A1N(n1928), .Y(top_core_KE_n3374) );
  OAI2BB2X1 U25818 ( .B0(n1499), .B1(n1943), .A0N(top_core_KE_key_mem_5__0_), 
        .A1N(n1947), .Y(top_core_KE_n3503) );
  OAI2BB2X1 U25819 ( .B0(n1499), .B1(n1964), .A0N(top_core_KE_key_mem_6__0_), 
        .A1N(n1964), .Y(top_core_KE_n3632) );
  OAI2BB2X1 U25820 ( .B0(n1499), .B1(n1983), .A0N(top_core_KE_key_mem_7__0_), 
        .A1N(n1987), .Y(top_core_KE_n3761) );
  OAI2BB2X1 U25821 ( .B0(n1499), .B1(n2044), .A0N(top_core_KE_key_mem_10__0_), 
        .A1N(n2048), .Y(top_core_KE_n4148) );
  OAI2BB2X1 U25822 ( .B0(n1499), .B1(n2063), .A0N(top_core_KE_key_mem_11__0_), 
        .A1N(n2067), .Y(top_core_KE_n4277) );
  OAI2BB2X1 U25823 ( .B0(n1499), .B1(n2083), .A0N(top_core_KE_key_mem_12__0_), 
        .A1N(n2087), .Y(top_core_KE_n4406) );
  OAI2BB2X1 U25824 ( .B0(n1499), .B1(n2103), .A0N(top_core_KE_key_mem_13__0_), 
        .A1N(n2107), .Y(top_core_KE_n4535) );
  OAI2BB2X1 U25825 ( .B0(n1499), .B1(n2123), .A0N(top_core_KE_key_mem_14__0_), 
        .A1N(n2127), .Y(top_core_KE_n4664) );
  OAI2BB2X1 U25826 ( .B0(n1372), .B1(n2004), .A0N(top_core_KE_key_mem_8__127_), 
        .A1N(n2007), .Y(top_core_KE_n3763) );
  OAI2BB2X1 U25827 ( .B0(n1373), .B1(n1997), .A0N(top_core_KE_key_mem_8__126_), 
        .A1N(n2006), .Y(top_core_KE_n3764) );
  OAI2BB2X1 U25828 ( .B0(n1374), .B1(n2004), .A0N(top_core_KE_key_mem_8__125_), 
        .A1N(n2007), .Y(top_core_KE_n3765) );
  OAI2BB2X1 U25829 ( .B0(n1375), .B1(n2004), .A0N(top_core_KE_key_mem_8__124_), 
        .A1N(n2006), .Y(top_core_KE_n3766) );
  OAI2BB2X1 U25830 ( .B0(n1376), .B1(n1998), .A0N(top_core_KE_key_mem_8__123_), 
        .A1N(n2006), .Y(top_core_KE_n3767) );
  OAI2BB2X1 U25831 ( .B0(n1377), .B1(n2003), .A0N(top_core_KE_key_mem_8__122_), 
        .A1N(n2006), .Y(top_core_KE_n3768) );
  OAI2BB2X1 U25832 ( .B0(n1378), .B1(n2001), .A0N(top_core_KE_key_mem_8__121_), 
        .A1N(n2006), .Y(top_core_KE_n3769) );
  OAI2BB2X1 U25833 ( .B0(n1379), .B1(n2003), .A0N(top_core_KE_key_mem_8__120_), 
        .A1N(n2005), .Y(top_core_KE_n3770) );
  OAI2BB2X1 U25834 ( .B0(n1380), .B1(n2003), .A0N(top_core_KE_key_mem_8__119_), 
        .A1N(n2007), .Y(top_core_KE_n3771) );
  OAI2BB2X1 U25835 ( .B0(n1381), .B1(n2003), .A0N(top_core_KE_key_mem_8__118_), 
        .A1N(n2005), .Y(top_core_KE_n3772) );
  OAI2BB2X1 U25836 ( .B0(n1382), .B1(n2002), .A0N(top_core_KE_key_mem_8__117_), 
        .A1N(n2005), .Y(top_core_KE_n3773) );
  OAI2BB2X1 U25837 ( .B0(n1383), .B1(n2002), .A0N(top_core_KE_key_mem_8__116_), 
        .A1N(n2006), .Y(top_core_KE_n3774) );
  OAI2BB2X1 U25838 ( .B0(n1384), .B1(n2002), .A0N(top_core_KE_key_mem_8__115_), 
        .A1N(n2005), .Y(top_core_KE_n3775) );
  OAI2BB2X1 U25839 ( .B0(n1385), .B1(n2002), .A0N(top_core_KE_key_mem_8__114_), 
        .A1N(n2005), .Y(top_core_KE_n3776) );
  OAI2BB2X1 U25840 ( .B0(n1386), .B1(n2002), .A0N(top_core_KE_key_mem_8__113_), 
        .A1N(n2006), .Y(top_core_KE_n3777) );
  OAI2BB2X1 U25841 ( .B0(n1387), .B1(n2001), .A0N(top_core_KE_key_mem_8__112_), 
        .A1N(n2004), .Y(top_core_KE_n3778) );
  OAI2BB2X1 U25842 ( .B0(n1388), .B1(n2001), .A0N(top_core_KE_key_mem_8__111_), 
        .A1N(n2004), .Y(top_core_KE_n3779) );
  OAI2BB2X1 U25843 ( .B0(n1389), .B1(n2001), .A0N(top_core_KE_key_mem_8__110_), 
        .A1N(n2004), .Y(top_core_KE_n3780) );
  OAI2BB2X1 U25844 ( .B0(n1390), .B1(n2000), .A0N(top_core_KE_key_mem_8__109_), 
        .A1N(n2004), .Y(top_core_KE_n3781) );
  OAI2BB2X1 U25845 ( .B0(n1391), .B1(n2000), .A0N(top_core_KE_key_mem_8__108_), 
        .A1N(n2005), .Y(top_core_KE_n3782) );
  OAI2BB2X1 U25846 ( .B0(n1392), .B1(n2000), .A0N(top_core_KE_key_mem_8__107_), 
        .A1N(n2005), .Y(top_core_KE_n3783) );
  OAI2BB2X1 U25847 ( .B0(n1393), .B1(n2000), .A0N(top_core_KE_key_mem_8__106_), 
        .A1N(n2005), .Y(top_core_KE_n3784) );
  OAI2BB2X1 U25848 ( .B0(n1394), .B1(n1999), .A0N(top_core_KE_key_mem_8__105_), 
        .A1N(n2005), .Y(top_core_KE_n3785) );
  OAI2BB2X1 U25849 ( .B0(n1395), .B1(n1999), .A0N(top_core_KE_key_mem_8__104_), 
        .A1N(n2005), .Y(top_core_KE_n3786) );
  OAI2BB2X1 U25850 ( .B0(n1396), .B1(n1999), .A0N(top_core_KE_key_mem_8__103_), 
        .A1N(n2005), .Y(top_core_KE_n3787) );
  OAI2BB2X1 U25851 ( .B0(n1397), .B1(n1999), .A0N(top_core_KE_key_mem_8__102_), 
        .A1N(n2007), .Y(top_core_KE_n3788) );
  OAI2BB2X1 U25852 ( .B0(n1398), .B1(top_core_KE_n882), .A0N(
        top_core_KE_key_mem_8__101_), .A1N(n2005), .Y(top_core_KE_n3789) );
  OAI2BB2X1 U25853 ( .B0(n1399), .B1(top_core_KE_n882), .A0N(
        top_core_KE_key_mem_8__100_), .A1N(n2005), .Y(top_core_KE_n3790) );
  OAI2BB2X1 U25854 ( .B0(n1400), .B1(n1998), .A0N(top_core_KE_key_mem_8__99_), 
        .A1N(n2005), .Y(top_core_KE_n3791) );
  OAI2BB2X1 U25855 ( .B0(n1401), .B1(n2003), .A0N(top_core_KE_key_mem_8__98_), 
        .A1N(n2005), .Y(top_core_KE_n3792) );
  OAI2BB2X1 U25856 ( .B0(n1402), .B1(n1999), .A0N(top_core_KE_key_mem_8__97_), 
        .A1N(n2006), .Y(top_core_KE_n3793) );
  OAI2BB2X1 U25857 ( .B0(n1403), .B1(n1998), .A0N(top_core_KE_key_mem_8__96_), 
        .A1N(n2006), .Y(top_core_KE_n3794) );
  OAI2BB2X1 U25858 ( .B0(n1404), .B1(n2003), .A0N(top_core_KE_key_mem_8__95_), 
        .A1N(n2006), .Y(top_core_KE_n3795) );
  OAI2BB2X1 U25859 ( .B0(n1405), .B1(n2008), .A0N(top_core_KE_key_mem_8__94_), 
        .A1N(n2006), .Y(top_core_KE_n3796) );
  OAI2BB2X1 U25860 ( .B0(n1406), .B1(n1998), .A0N(top_core_KE_key_mem_8__93_), 
        .A1N(n2006), .Y(top_core_KE_n3797) );
  OAI2BB2X1 U25861 ( .B0(n1407), .B1(n1998), .A0N(top_core_KE_key_mem_8__92_), 
        .A1N(n2006), .Y(top_core_KE_n3798) );
  OAI2BB2X1 U25862 ( .B0(n1408), .B1(n1998), .A0N(top_core_KE_key_mem_8__91_), 
        .A1N(n2006), .Y(top_core_KE_n3799) );
  OAI2BB2X1 U25863 ( .B0(n1409), .B1(n1998), .A0N(top_core_KE_key_mem_8__90_), 
        .A1N(n2006), .Y(top_core_KE_n3800) );
  OAI2BB2X1 U25864 ( .B0(n1410), .B1(n1997), .A0N(top_core_KE_key_mem_8__89_), 
        .A1N(n2007), .Y(top_core_KE_n3801) );
  OAI2BB2X1 U25865 ( .B0(n1411), .B1(n1997), .A0N(top_core_KE_key_mem_8__88_), 
        .A1N(n2007), .Y(top_core_KE_n3802) );
  OAI2BB2X1 U25866 ( .B0(n1412), .B1(n1997), .A0N(top_core_KE_key_mem_8__87_), 
        .A1N(n2007), .Y(top_core_KE_n3803) );
  OAI2BB2X1 U25867 ( .B0(n1413), .B1(n1997), .A0N(top_core_KE_key_mem_8__86_), 
        .A1N(n2007), .Y(top_core_KE_n3804) );
  OAI2BB2X1 U25868 ( .B0(n1414), .B1(n2001), .A0N(top_core_KE_key_mem_8__85_), 
        .A1N(n2007), .Y(top_core_KE_n3805) );
  OAI2BB2X1 U25869 ( .B0(n1415), .B1(n1997), .A0N(top_core_KE_key_mem_8__84_), 
        .A1N(n2007), .Y(top_core_KE_n3806) );
  OAI2BB2X1 U25870 ( .B0(n1416), .B1(n1997), .A0N(top_core_KE_key_mem_8__83_), 
        .A1N(n2007), .Y(top_core_KE_n3807) );
  OAI2BB2X1 U25871 ( .B0(n1417), .B1(n1997), .A0N(top_core_KE_key_mem_8__82_), 
        .A1N(n2007), .Y(top_core_KE_n3808) );
  OAI2BB2X1 U25872 ( .B0(n1418), .B1(n1997), .A0N(top_core_KE_key_mem_8__81_), 
        .A1N(n2008), .Y(top_core_KE_n3809) );
  OAI2BB2X1 U25873 ( .B0(n1419), .B1(n1997), .A0N(top_core_KE_key_mem_8__80_), 
        .A1N(n2008), .Y(top_core_KE_n3810) );
  OAI2BB2X1 U25874 ( .B0(n1420), .B1(n1997), .A0N(top_core_KE_key_mem_8__79_), 
        .A1N(n2008), .Y(top_core_KE_n3811) );
  OAI2BB2X1 U25875 ( .B0(n1421), .B1(n1997), .A0N(top_core_KE_key_mem_8__78_), 
        .A1N(n2008), .Y(top_core_KE_n3812) );
  OAI2BB2X1 U25876 ( .B0(n1422), .B1(n1998), .A0N(top_core_KE_key_mem_8__77_), 
        .A1N(n2008), .Y(top_core_KE_n3813) );
  OAI2BB2X1 U25877 ( .B0(n1423), .B1(n1998), .A0N(top_core_KE_key_mem_8__76_), 
        .A1N(n2008), .Y(top_core_KE_n3814) );
  OAI2BB2X1 U25878 ( .B0(n1424), .B1(n1998), .A0N(top_core_KE_key_mem_8__75_), 
        .A1N(n2008), .Y(top_core_KE_n3815) );
  OAI2BB2X1 U25879 ( .B0(n1425), .B1(n1998), .A0N(top_core_KE_key_mem_8__74_), 
        .A1N(n2008), .Y(top_core_KE_n3816) );
  OAI2BB2X1 U25880 ( .B0(n1426), .B1(n1998), .A0N(top_core_KE_key_mem_8__73_), 
        .A1N(n2008), .Y(top_core_KE_n3817) );
  OAI2BB2X1 U25881 ( .B0(n1427), .B1(n1998), .A0N(top_core_KE_key_mem_8__72_), 
        .A1N(n2008), .Y(top_core_KE_n3818) );
  OAI2BB2X1 U25882 ( .B0(n1428), .B1(n1998), .A0N(top_core_KE_key_mem_8__71_), 
        .A1N(n2008), .Y(top_core_KE_n3819) );
  OAI2BB2X1 U25883 ( .B0(n1429), .B1(n1998), .A0N(top_core_KE_key_mem_8__70_), 
        .A1N(n2008), .Y(top_core_KE_n3820) );
  OAI2BB2X1 U25884 ( .B0(n1430), .B1(n2012), .A0N(top_core_KE_key_mem_8__69_), 
        .A1N(n2008), .Y(top_core_KE_n3821) );
  OAI2BB2X1 U25885 ( .B0(n1431), .B1(n2006), .A0N(top_core_KE_key_mem_8__68_), 
        .A1N(n2008), .Y(top_core_KE_n3822) );
  OAI2BB2X1 U25886 ( .B0(n1432), .B1(n2007), .A0N(top_core_KE_key_mem_8__67_), 
        .A1N(n2008), .Y(top_core_KE_n3823) );
  OAI2BB2X1 U25887 ( .B0(n1433), .B1(n2005), .A0N(top_core_KE_key_mem_8__66_), 
        .A1N(n2009), .Y(top_core_KE_n3824) );
  OAI2BB2X1 U25888 ( .B0(n1434), .B1(n2010), .A0N(top_core_KE_key_mem_8__65_), 
        .A1N(n2009), .Y(top_core_KE_n3825) );
  OAI2BB2X1 U25889 ( .B0(n1435), .B1(n2011), .A0N(top_core_KE_key_mem_8__64_), 
        .A1N(n2009), .Y(top_core_KE_n3826) );
  OAI2BB2X1 U25890 ( .B0(n1436), .B1(n2004), .A0N(top_core_KE_key_mem_8__63_), 
        .A1N(n2009), .Y(top_core_KE_n3827) );
  OAI2BB2X1 U25891 ( .B0(n1437), .B1(n2001), .A0N(top_core_KE_key_mem_8__62_), 
        .A1N(n2009), .Y(top_core_KE_n3828) );
  OAI2BB2X1 U25892 ( .B0(n1438), .B1(n2001), .A0N(top_core_KE_key_mem_8__61_), 
        .A1N(n2009), .Y(top_core_KE_n3829) );
  OAI2BB2X1 U25893 ( .B0(n1439), .B1(n2002), .A0N(top_core_KE_key_mem_8__60_), 
        .A1N(n2009), .Y(top_core_KE_n3830) );
  OAI2BB2X1 U25894 ( .B0(n1440), .B1(top_core_KE_n882), .A0N(
        top_core_KE_key_mem_8__59_), .A1N(n2009), .Y(top_core_KE_n3831) );
  OAI2BB2X1 U25895 ( .B0(n1441), .B1(n2000), .A0N(top_core_KE_key_mem_8__58_), 
        .A1N(n2009), .Y(top_core_KE_n3832) );
  OAI2BB2X1 U25896 ( .B0(n1442), .B1(n2002), .A0N(top_core_KE_key_mem_8__57_), 
        .A1N(n2009), .Y(top_core_KE_n3833) );
  OAI2BB2X1 U25897 ( .B0(n1443), .B1(n2004), .A0N(top_core_KE_key_mem_8__56_), 
        .A1N(n2009), .Y(top_core_KE_n3834) );
  OAI2BB2X1 U25898 ( .B0(n1444), .B1(n1997), .A0N(top_core_KE_key_mem_8__55_), 
        .A1N(n2009), .Y(top_core_KE_n3835) );
  OAI2BB2X1 U25899 ( .B0(n1445), .B1(n1999), .A0N(top_core_KE_key_mem_8__54_), 
        .A1N(n2009), .Y(top_core_KE_n3836) );
  OAI2BB2X1 U25900 ( .B0(n1446), .B1(n1999), .A0N(top_core_KE_key_mem_8__53_), 
        .A1N(n2009), .Y(top_core_KE_n3837) );
  OAI2BB2X1 U25901 ( .B0(n1447), .B1(n1999), .A0N(top_core_KE_key_mem_8__52_), 
        .A1N(n2009), .Y(top_core_KE_n3838) );
  OAI2BB2X1 U25902 ( .B0(n1448), .B1(n1999), .A0N(top_core_KE_key_mem_8__51_), 
        .A1N(n2010), .Y(top_core_KE_n3839) );
  OAI2BB2X1 U25903 ( .B0(n1449), .B1(n1999), .A0N(top_core_KE_key_mem_8__50_), 
        .A1N(n2010), .Y(top_core_KE_n3840) );
  OAI2BB2X1 U25904 ( .B0(n1450), .B1(n1999), .A0N(top_core_KE_key_mem_8__49_), 
        .A1N(n2010), .Y(top_core_KE_n3841) );
  OAI2BB2X1 U25905 ( .B0(n1451), .B1(n1999), .A0N(top_core_KE_key_mem_8__48_), 
        .A1N(n2010), .Y(top_core_KE_n3842) );
  OAI2BB2X1 U25906 ( .B0(n1452), .B1(n1999), .A0N(top_core_KE_key_mem_8__47_), 
        .A1N(n2010), .Y(top_core_KE_n3843) );
  OAI2BB2X1 U25907 ( .B0(n1453), .B1(n1999), .A0N(top_core_KE_key_mem_8__46_), 
        .A1N(n2010), .Y(top_core_KE_n3844) );
  OAI2BB2X1 U25908 ( .B0(n1454), .B1(n2000), .A0N(top_core_KE_key_mem_8__45_), 
        .A1N(n2010), .Y(top_core_KE_n3845) );
  OAI2BB2X1 U25909 ( .B0(n1455), .B1(n2000), .A0N(top_core_KE_key_mem_8__44_), 
        .A1N(n2010), .Y(top_core_KE_n3846) );
  OAI2BB2X1 U25910 ( .B0(n1456), .B1(n2000), .A0N(top_core_KE_key_mem_8__43_), 
        .A1N(n2010), .Y(top_core_KE_n3847) );
  OAI2BB2X1 U25911 ( .B0(n1457), .B1(n2000), .A0N(top_core_KE_key_mem_8__42_), 
        .A1N(n2010), .Y(top_core_KE_n3848) );
  OAI2BB2X1 U25912 ( .B0(n1458), .B1(n2000), .A0N(top_core_KE_key_mem_8__41_), 
        .A1N(n2010), .Y(top_core_KE_n3849) );
  OAI2BB2X1 U25913 ( .B0(n1459), .B1(n2000), .A0N(top_core_KE_key_mem_8__40_), 
        .A1N(n2010), .Y(top_core_KE_n3850) );
  OAI2BB2X1 U25914 ( .B0(n1460), .B1(n2000), .A0N(top_core_KE_key_mem_8__39_), 
        .A1N(n2010), .Y(top_core_KE_n3851) );
  OAI2BB2X1 U25915 ( .B0(n1461), .B1(n2000), .A0N(top_core_KE_key_mem_8__38_), 
        .A1N(n2010), .Y(top_core_KE_n3852) );
  OAI2BB2X1 U25916 ( .B0(n1462), .B1(n2001), .A0N(top_core_KE_key_mem_8__37_), 
        .A1N(n2010), .Y(top_core_KE_n3853) );
  OAI2BB2X1 U25917 ( .B0(n1463), .B1(n2001), .A0N(top_core_KE_key_mem_8__36_), 
        .A1N(n2011), .Y(top_core_KE_n3854) );
  OAI2BB2X1 U25918 ( .B0(n1464), .B1(n2001), .A0N(top_core_KE_key_mem_8__35_), 
        .A1N(n2011), .Y(top_core_KE_n3855) );
  OAI2BB2X1 U25919 ( .B0(n1465), .B1(n2001), .A0N(top_core_KE_key_mem_8__34_), 
        .A1N(n2011), .Y(top_core_KE_n3856) );
  OAI2BB2X1 U25920 ( .B0(n1466), .B1(n2001), .A0N(top_core_KE_key_mem_8__33_), 
        .A1N(n2011), .Y(top_core_KE_n3857) );
  OAI2BB2X1 U25921 ( .B0(n1467), .B1(n2001), .A0N(top_core_KE_key_mem_8__32_), 
        .A1N(n2011), .Y(top_core_KE_n3858) );
  OAI2BB2X1 U25922 ( .B0(n1468), .B1(n2001), .A0N(top_core_KE_key_mem_8__31_), 
        .A1N(n2011), .Y(top_core_KE_n3859) );
  OAI2BB2X1 U25923 ( .B0(n1469), .B1(n2001), .A0N(top_core_KE_key_mem_8__30_), 
        .A1N(n2011), .Y(top_core_KE_n3860) );
  OAI2BB2X1 U25924 ( .B0(n1470), .B1(n2002), .A0N(top_core_KE_key_mem_8__29_), 
        .A1N(n2011), .Y(top_core_KE_n3861) );
  OAI2BB2X1 U25925 ( .B0(n1471), .B1(n2002), .A0N(top_core_KE_key_mem_8__28_), 
        .A1N(n2011), .Y(top_core_KE_n3862) );
  OAI2BB2X1 U25926 ( .B0(n1472), .B1(n2002), .A0N(top_core_KE_key_mem_8__27_), 
        .A1N(n2011), .Y(top_core_KE_n3863) );
  OAI2BB2X1 U25927 ( .B0(n1473), .B1(n2002), .A0N(top_core_KE_key_mem_8__26_), 
        .A1N(n2011), .Y(top_core_KE_n3864) );
  OAI2BB2X1 U25928 ( .B0(n1474), .B1(n2002), .A0N(top_core_KE_key_mem_8__25_), 
        .A1N(n2011), .Y(top_core_KE_n3865) );
  OAI2BB2X1 U25929 ( .B0(n1475), .B1(n2002), .A0N(top_core_KE_key_mem_8__24_), 
        .A1N(n2011), .Y(top_core_KE_n3866) );
  OAI2BB2X1 U25930 ( .B0(n1476), .B1(n2003), .A0N(top_core_KE_key_mem_8__23_), 
        .A1N(n2011), .Y(top_core_KE_n3867) );
  OAI2BB2X1 U25931 ( .B0(n1477), .B1(n2003), .A0N(top_core_KE_key_mem_8__22_), 
        .A1N(n2011), .Y(top_core_KE_n3868) );
  OAI2BB2X1 U25932 ( .B0(n1478), .B1(n2002), .A0N(top_core_KE_key_mem_8__21_), 
        .A1N(n2012), .Y(top_core_KE_n3869) );
  OAI2BB2X1 U25933 ( .B0(n1479), .B1(n2003), .A0N(top_core_KE_key_mem_8__20_), 
        .A1N(n2012), .Y(top_core_KE_n3870) );
  OAI2BB2X1 U25934 ( .B0(n1480), .B1(n2003), .A0N(top_core_KE_key_mem_8__19_), 
        .A1N(n2012), .Y(top_core_KE_n3871) );
  OAI2BB2X1 U25935 ( .B0(n1481), .B1(n2003), .A0N(top_core_KE_key_mem_8__18_), 
        .A1N(n2012), .Y(top_core_KE_n3872) );
  OAI2BB2X1 U25936 ( .B0(n1482), .B1(n2003), .A0N(top_core_KE_key_mem_8__17_), 
        .A1N(n2012), .Y(top_core_KE_n3873) );
  OAI2BB2X1 U25937 ( .B0(n1483), .B1(n2002), .A0N(top_core_KE_key_mem_8__16_), 
        .A1N(n2012), .Y(top_core_KE_n3874) );
  OAI2BB2X1 U25938 ( .B0(n1484), .B1(n2003), .A0N(top_core_KE_key_mem_8__15_), 
        .A1N(n2012), .Y(top_core_KE_n3875) );
  OAI2BB2X1 U25939 ( .B0(n1485), .B1(n2000), .A0N(top_core_KE_key_mem_8__14_), 
        .A1N(n2012), .Y(top_core_KE_n3876) );
  OAI2BB2X1 U25940 ( .B0(n1486), .B1(n2004), .A0N(top_core_KE_key_mem_8__13_), 
        .A1N(n2012), .Y(top_core_KE_n3877) );
  OAI2BB2X1 U25941 ( .B0(n1487), .B1(n2003), .A0N(top_core_KE_key_mem_8__12_), 
        .A1N(n2012), .Y(top_core_KE_n3878) );
  OAI2BB2X1 U25942 ( .B0(n1488), .B1(n1999), .A0N(top_core_KE_key_mem_8__11_), 
        .A1N(n2012), .Y(top_core_KE_n3879) );
  OAI2BB2X1 U25943 ( .B0(n1489), .B1(n1997), .A0N(top_core_KE_key_mem_8__10_), 
        .A1N(n2012), .Y(top_core_KE_n3880) );
  OAI2BB2X1 U25944 ( .B0(n1490), .B1(n2000), .A0N(top_core_KE_key_mem_8__9_), 
        .A1N(n2012), .Y(top_core_KE_n3881) );
  OAI2BB2X1 U25945 ( .B0(n1491), .B1(n2004), .A0N(top_core_KE_key_mem_8__8_), 
        .A1N(n2012), .Y(top_core_KE_n3882) );
  OAI2BB2X1 U25946 ( .B0(n1492), .B1(n2003), .A0N(top_core_KE_key_mem_8__7_), 
        .A1N(n2012), .Y(top_core_KE_n3883) );
  OAI2BB2X1 U25947 ( .B0(n1493), .B1(n1998), .A0N(top_core_KE_key_mem_8__6_), 
        .A1N(n2000), .Y(top_core_KE_n3884) );
  OAI2BB2X1 U25948 ( .B0(n1494), .B1(n2004), .A0N(top_core_KE_key_mem_8__5_), 
        .A1N(n2001), .Y(top_core_KE_n3885) );
  OAI2BB2X1 U25949 ( .B0(n1495), .B1(n2004), .A0N(top_core_KE_key_mem_8__4_), 
        .A1N(n2002), .Y(top_core_KE_n3886) );
  OAI2BB2X1 U25950 ( .B0(n1496), .B1(n2004), .A0N(top_core_KE_key_mem_8__3_), 
        .A1N(n2008), .Y(top_core_KE_n3887) );
  OAI2BB2X1 U25951 ( .B0(n1497), .B1(n2004), .A0N(top_core_KE_key_mem_8__2_), 
        .A1N(n2009), .Y(top_core_KE_n3888) );
  OAI2BB2X1 U25952 ( .B0(n1498), .B1(n2004), .A0N(top_core_KE_key_mem_8__1_), 
        .A1N(n2007), .Y(top_core_KE_n3889) );
  OAI2BB2X1 U25953 ( .B0(n1499), .B1(n2003), .A0N(top_core_KE_key_mem_8__0_), 
        .A1N(n2007), .Y(top_core_KE_n3890) );
  OAI2BB2X1 U25954 ( .B0(n1372), .B1(n2024), .A0N(top_core_KE_key_mem_9__127_), 
        .A1N(n2027), .Y(top_core_KE_n3892) );
  OAI2BB2X1 U25955 ( .B0(n1373), .B1(n2018), .A0N(top_core_KE_key_mem_9__126_), 
        .A1N(n2026), .Y(top_core_KE_n3893) );
  OAI2BB2X1 U25956 ( .B0(n1374), .B1(n2024), .A0N(top_core_KE_key_mem_9__125_), 
        .A1N(n2027), .Y(top_core_KE_n3894) );
  OAI2BB2X1 U25957 ( .B0(n1375), .B1(n2024), .A0N(top_core_KE_key_mem_9__124_), 
        .A1N(n2026), .Y(top_core_KE_n3895) );
  OAI2BB2X1 U25958 ( .B0(n1376), .B1(n2017), .A0N(top_core_KE_key_mem_9__123_), 
        .A1N(n2026), .Y(top_core_KE_n3896) );
  OAI2BB2X1 U25959 ( .B0(n1377), .B1(n2023), .A0N(top_core_KE_key_mem_9__122_), 
        .A1N(n2026), .Y(top_core_KE_n3897) );
  OAI2BB2X1 U25960 ( .B0(n1378), .B1(n2021), .A0N(top_core_KE_key_mem_9__121_), 
        .A1N(n2026), .Y(top_core_KE_n3898) );
  OAI2BB2X1 U25961 ( .B0(n1379), .B1(n2023), .A0N(top_core_KE_key_mem_9__120_), 
        .A1N(n2025), .Y(top_core_KE_n3899) );
  OAI2BB2X1 U25962 ( .B0(n1380), .B1(n2023), .A0N(top_core_KE_key_mem_9__119_), 
        .A1N(n2027), .Y(top_core_KE_n3900) );
  OAI2BB2X1 U25963 ( .B0(n1381), .B1(n2023), .A0N(top_core_KE_key_mem_9__118_), 
        .A1N(n2025), .Y(top_core_KE_n3901) );
  OAI2BB2X1 U25964 ( .B0(n1382), .B1(n2022), .A0N(top_core_KE_key_mem_9__117_), 
        .A1N(n2025), .Y(top_core_KE_n3902) );
  OAI2BB2X1 U25965 ( .B0(n1383), .B1(n2022), .A0N(top_core_KE_key_mem_9__116_), 
        .A1N(n2026), .Y(top_core_KE_n3903) );
  OAI2BB2X1 U25966 ( .B0(n1384), .B1(n2022), .A0N(top_core_KE_key_mem_9__115_), 
        .A1N(n2025), .Y(top_core_KE_n3904) );
  OAI2BB2X1 U25967 ( .B0(n1385), .B1(n2022), .A0N(top_core_KE_key_mem_9__114_), 
        .A1N(n2025), .Y(top_core_KE_n3905) );
  OAI2BB2X1 U25968 ( .B0(n1386), .B1(n2022), .A0N(top_core_KE_key_mem_9__113_), 
        .A1N(n2026), .Y(top_core_KE_n3906) );
  OAI2BB2X1 U25969 ( .B0(n1387), .B1(n2021), .A0N(top_core_KE_key_mem_9__112_), 
        .A1N(n2024), .Y(top_core_KE_n3907) );
  OAI2BB2X1 U25970 ( .B0(n1388), .B1(n2021), .A0N(top_core_KE_key_mem_9__111_), 
        .A1N(n2024), .Y(top_core_KE_n3908) );
  OAI2BB2X1 U25971 ( .B0(n1389), .B1(n2021), .A0N(top_core_KE_key_mem_9__110_), 
        .A1N(n2024), .Y(top_core_KE_n3909) );
  OAI2BB2X1 U25972 ( .B0(n1390), .B1(n2020), .A0N(top_core_KE_key_mem_9__109_), 
        .A1N(n2024), .Y(top_core_KE_n3910) );
  OAI2BB2X1 U25973 ( .B0(n1391), .B1(n2020), .A0N(top_core_KE_key_mem_9__108_), 
        .A1N(n2025), .Y(top_core_KE_n3911) );
  OAI2BB2X1 U25974 ( .B0(n1392), .B1(n2020), .A0N(top_core_KE_key_mem_9__107_), 
        .A1N(n2025), .Y(top_core_KE_n3912) );
  OAI2BB2X1 U25975 ( .B0(n1393), .B1(n2020), .A0N(top_core_KE_key_mem_9__106_), 
        .A1N(n2025), .Y(top_core_KE_n3913) );
  OAI2BB2X1 U25976 ( .B0(n1394), .B1(n2019), .A0N(top_core_KE_key_mem_9__105_), 
        .A1N(n2025), .Y(top_core_KE_n3914) );
  OAI2BB2X1 U25977 ( .B0(n1395), .B1(n2019), .A0N(top_core_KE_key_mem_9__104_), 
        .A1N(n2025), .Y(top_core_KE_n3915) );
  OAI2BB2X1 U25978 ( .B0(n1396), .B1(n2019), .A0N(top_core_KE_key_mem_9__103_), 
        .A1N(n2025), .Y(top_core_KE_n3916) );
  OAI2BB2X1 U25979 ( .B0(n1397), .B1(n2019), .A0N(top_core_KE_key_mem_9__102_), 
        .A1N(n2027), .Y(top_core_KE_n3917) );
  OAI2BB2X1 U25980 ( .B0(n1398), .B1(top_core_KE_n885), .A0N(
        top_core_KE_key_mem_9__101_), .A1N(n2025), .Y(top_core_KE_n3918) );
  OAI2BB2X1 U25981 ( .B0(n1399), .B1(top_core_KE_n885), .A0N(
        top_core_KE_key_mem_9__100_), .A1N(n2025), .Y(top_core_KE_n3919) );
  OAI2BB2X1 U25982 ( .B0(n1400), .B1(n2017), .A0N(top_core_KE_key_mem_9__99_), 
        .A1N(n2025), .Y(top_core_KE_n3920) );
  OAI2BB2X1 U25983 ( .B0(n1401), .B1(n2023), .A0N(top_core_KE_key_mem_9__98_), 
        .A1N(n2025), .Y(top_core_KE_n3921) );
  OAI2BB2X1 U25984 ( .B0(n1402), .B1(n2018), .A0N(top_core_KE_key_mem_9__97_), 
        .A1N(n2026), .Y(top_core_KE_n3922) );
  OAI2BB2X1 U25985 ( .B0(n1403), .B1(n2018), .A0N(top_core_KE_key_mem_9__96_), 
        .A1N(n2026), .Y(top_core_KE_n3923) );
  OAI2BB2X1 U25986 ( .B0(n1404), .B1(n2018), .A0N(top_core_KE_key_mem_9__95_), 
        .A1N(n2026), .Y(top_core_KE_n3924) );
  OAI2BB2X1 U25987 ( .B0(n1405), .B1(n2018), .A0N(top_core_KE_key_mem_9__94_), 
        .A1N(n2026), .Y(top_core_KE_n3925) );
  OAI2BB2X1 U25988 ( .B0(n1406), .B1(n2017), .A0N(top_core_KE_key_mem_9__93_), 
        .A1N(n2026), .Y(top_core_KE_n3926) );
  OAI2BB2X1 U25989 ( .B0(n1407), .B1(n2017), .A0N(top_core_KE_key_mem_9__92_), 
        .A1N(n2026), .Y(top_core_KE_n3927) );
  OAI2BB2X1 U25990 ( .B0(n1408), .B1(n2017), .A0N(top_core_KE_key_mem_9__91_), 
        .A1N(n2026), .Y(top_core_KE_n3928) );
  OAI2BB2X1 U25991 ( .B0(n1409), .B1(n2017), .A0N(top_core_KE_key_mem_9__90_), 
        .A1N(n2026), .Y(top_core_KE_n3929) );
  OAI2BB2X1 U25992 ( .B0(n1410), .B1(n2020), .A0N(top_core_KE_key_mem_9__89_), 
        .A1N(n2027), .Y(top_core_KE_n3930) );
  OAI2BB2X1 U25993 ( .B0(n1411), .B1(n2019), .A0N(top_core_KE_key_mem_9__88_), 
        .A1N(n2027), .Y(top_core_KE_n3931) );
  OAI2BB2X1 U25994 ( .B0(n1412), .B1(n2018), .A0N(top_core_KE_key_mem_9__87_), 
        .A1N(n2027), .Y(top_core_KE_n3932) );
  OAI2BB2X1 U25995 ( .B0(n1413), .B1(n2017), .A0N(top_core_KE_key_mem_9__86_), 
        .A1N(n2027), .Y(top_core_KE_n3933) );
  OAI2BB2X1 U25996 ( .B0(n1414), .B1(n2021), .A0N(top_core_KE_key_mem_9__85_), 
        .A1N(n2027), .Y(top_core_KE_n3934) );
  OAI2BB2X1 U25997 ( .B0(n1415), .B1(n2028), .A0N(top_core_KE_key_mem_9__84_), 
        .A1N(n2027), .Y(top_core_KE_n3935) );
  OAI2BB2X1 U25998 ( .B0(n1416), .B1(n2029), .A0N(top_core_KE_key_mem_9__83_), 
        .A1N(n2027), .Y(top_core_KE_n3936) );
  OAI2BB2X1 U25999 ( .B0(n1417), .B1(n2032), .A0N(top_core_KE_key_mem_9__82_), 
        .A1N(n2027), .Y(top_core_KE_n3937) );
  OAI2BB2X1 U26000 ( .B0(n1418), .B1(n2032), .A0N(top_core_KE_key_mem_9__81_), 
        .A1N(n2028), .Y(top_core_KE_n3938) );
  OAI2BB2X1 U26001 ( .B0(n1419), .B1(n2026), .A0N(top_core_KE_key_mem_9__80_), 
        .A1N(n2028), .Y(top_core_KE_n3939) );
  OAI2BB2X1 U26002 ( .B0(n1420), .B1(n2027), .A0N(top_core_KE_key_mem_9__79_), 
        .A1N(n2028), .Y(top_core_KE_n3940) );
  OAI2BB2X1 U26003 ( .B0(n1421), .B1(n2030), .A0N(top_core_KE_key_mem_9__78_), 
        .A1N(n2028), .Y(top_core_KE_n3941) );
  OAI2BB2X1 U26004 ( .B0(n1422), .B1(n2017), .A0N(top_core_KE_key_mem_9__77_), 
        .A1N(n2028), .Y(top_core_KE_n3942) );
  OAI2BB2X1 U26005 ( .B0(n1423), .B1(n2017), .A0N(top_core_KE_key_mem_9__76_), 
        .A1N(n2028), .Y(top_core_KE_n3943) );
  OAI2BB2X1 U26006 ( .B0(n1424), .B1(n2017), .A0N(top_core_KE_key_mem_9__75_), 
        .A1N(n2028), .Y(top_core_KE_n3944) );
  OAI2BB2X1 U26007 ( .B0(n1425), .B1(n2017), .A0N(top_core_KE_key_mem_9__74_), 
        .A1N(n2028), .Y(top_core_KE_n3945) );
  OAI2BB2X1 U26008 ( .B0(n1426), .B1(n2017), .A0N(top_core_KE_key_mem_9__73_), 
        .A1N(n2028), .Y(top_core_KE_n3946) );
  OAI2BB2X1 U26009 ( .B0(n1427), .B1(n2017), .A0N(top_core_KE_key_mem_9__72_), 
        .A1N(n2028), .Y(top_core_KE_n3947) );
  OAI2BB2X1 U26010 ( .B0(n1428), .B1(n2017), .A0N(top_core_KE_key_mem_9__71_), 
        .A1N(n2028), .Y(top_core_KE_n3948) );
  OAI2BB2X1 U26011 ( .B0(n1429), .B1(n2017), .A0N(top_core_KE_key_mem_9__70_), 
        .A1N(n2028), .Y(top_core_KE_n3949) );
  OAI2BB2X1 U26012 ( .B0(n1430), .B1(n2018), .A0N(top_core_KE_key_mem_9__69_), 
        .A1N(n2028), .Y(top_core_KE_n3950) );
  OAI2BB2X1 U26013 ( .B0(n1431), .B1(n2018), .A0N(top_core_KE_key_mem_9__68_), 
        .A1N(n2028), .Y(top_core_KE_n3951) );
  OAI2BB2X1 U26014 ( .B0(n1432), .B1(n2018), .A0N(top_core_KE_key_mem_9__67_), 
        .A1N(n2028), .Y(top_core_KE_n3952) );
  OAI2BB2X1 U26015 ( .B0(n1433), .B1(n2018), .A0N(top_core_KE_key_mem_9__66_), 
        .A1N(n2029), .Y(top_core_KE_n3953) );
  OAI2BB2X1 U26016 ( .B0(n1434), .B1(n2018), .A0N(top_core_KE_key_mem_9__65_), 
        .A1N(n2029), .Y(top_core_KE_n3954) );
  OAI2BB2X1 U26017 ( .B0(n1435), .B1(n2018), .A0N(top_core_KE_key_mem_9__64_), 
        .A1N(n2029), .Y(top_core_KE_n3955) );
  OAI2BB2X1 U26018 ( .B0(n1436), .B1(n2018), .A0N(top_core_KE_key_mem_9__63_), 
        .A1N(n2029), .Y(top_core_KE_n3956) );
  OAI2BB2X1 U26019 ( .B0(n1437), .B1(n2018), .A0N(top_core_KE_key_mem_9__62_), 
        .A1N(n2029), .Y(top_core_KE_n3957) );
  OAI2BB2X1 U26020 ( .B0(n1438), .B1(n2021), .A0N(top_core_KE_key_mem_9__61_), 
        .A1N(n2029), .Y(top_core_KE_n3958) );
  OAI2BB2X1 U26021 ( .B0(n1439), .B1(n2022), .A0N(top_core_KE_key_mem_9__60_), 
        .A1N(n2029), .Y(top_core_KE_n3959) );
  OAI2BB2X1 U26022 ( .B0(n1440), .B1(top_core_KE_n885), .A0N(
        top_core_KE_key_mem_9__59_), .A1N(n2029), .Y(top_core_KE_n3960) );
  OAI2BB2X1 U26023 ( .B0(n1441), .B1(n2020), .A0N(top_core_KE_key_mem_9__58_), 
        .A1N(n2029), .Y(top_core_KE_n3961) );
  OAI2BB2X1 U26024 ( .B0(n1442), .B1(n2018), .A0N(top_core_KE_key_mem_9__57_), 
        .A1N(n2029), .Y(top_core_KE_n3962) );
  OAI2BB2X1 U26025 ( .B0(n1443), .B1(n2024), .A0N(top_core_KE_key_mem_9__56_), 
        .A1N(n2029), .Y(top_core_KE_n3963) );
  OAI2BB2X1 U26026 ( .B0(n1444), .B1(n2031), .A0N(top_core_KE_key_mem_9__55_), 
        .A1N(n2029), .Y(top_core_KE_n3964) );
  OAI2BB2X1 U26027 ( .B0(n1445), .B1(n2019), .A0N(top_core_KE_key_mem_9__54_), 
        .A1N(n2029), .Y(top_core_KE_n3965) );
  OAI2BB2X1 U26028 ( .B0(n1446), .B1(n2019), .A0N(top_core_KE_key_mem_9__53_), 
        .A1N(n2029), .Y(top_core_KE_n3966) );
  OAI2BB2X1 U26029 ( .B0(n1447), .B1(n2019), .A0N(top_core_KE_key_mem_9__52_), 
        .A1N(n2029), .Y(top_core_KE_n3967) );
  OAI2BB2X1 U26030 ( .B0(n1448), .B1(n2019), .A0N(top_core_KE_key_mem_9__51_), 
        .A1N(n2030), .Y(top_core_KE_n3968) );
  OAI2BB2X1 U26031 ( .B0(n1449), .B1(n2019), .A0N(top_core_KE_key_mem_9__50_), 
        .A1N(n2030), .Y(top_core_KE_n3969) );
  OAI2BB2X1 U26032 ( .B0(n1450), .B1(n2019), .A0N(top_core_KE_key_mem_9__49_), 
        .A1N(n2030), .Y(top_core_KE_n3970) );
  OAI2BB2X1 U26033 ( .B0(n1451), .B1(n2019), .A0N(top_core_KE_key_mem_9__48_), 
        .A1N(n2030), .Y(top_core_KE_n3971) );
  OAI2BB2X1 U26034 ( .B0(n1452), .B1(n2019), .A0N(top_core_KE_key_mem_9__47_), 
        .A1N(n2030), .Y(top_core_KE_n3972) );
  OAI2BB2X1 U26035 ( .B0(n1453), .B1(n2019), .A0N(top_core_KE_key_mem_9__46_), 
        .A1N(n2030), .Y(top_core_KE_n3973) );
  OAI2BB2X1 U26036 ( .B0(n1454), .B1(n2020), .A0N(top_core_KE_key_mem_9__45_), 
        .A1N(n2030), .Y(top_core_KE_n3974) );
  OAI2BB2X1 U26037 ( .B0(n1455), .B1(n2020), .A0N(top_core_KE_key_mem_9__44_), 
        .A1N(n2030), .Y(top_core_KE_n3975) );
  OAI2BB2X1 U26038 ( .B0(n1456), .B1(n2020), .A0N(top_core_KE_key_mem_9__43_), 
        .A1N(n2030), .Y(top_core_KE_n3976) );
  OAI2BB2X1 U26039 ( .B0(n1457), .B1(n2020), .A0N(top_core_KE_key_mem_9__42_), 
        .A1N(n2030), .Y(top_core_KE_n3977) );
  OAI2BB2X1 U26040 ( .B0(n1458), .B1(n2020), .A0N(top_core_KE_key_mem_9__41_), 
        .A1N(n2030), .Y(top_core_KE_n3978) );
  OAI2BB2X1 U26041 ( .B0(n1459), .B1(n2020), .A0N(top_core_KE_key_mem_9__40_), 
        .A1N(n2030), .Y(top_core_KE_n3979) );
  OAI2BB2X1 U26042 ( .B0(n1460), .B1(n2020), .A0N(top_core_KE_key_mem_9__39_), 
        .A1N(n2030), .Y(top_core_KE_n3980) );
  OAI2BB2X1 U26043 ( .B0(n1461), .B1(n2020), .A0N(top_core_KE_key_mem_9__38_), 
        .A1N(n2030), .Y(top_core_KE_n3981) );
  OAI2BB2X1 U26044 ( .B0(n1462), .B1(n2021), .A0N(top_core_KE_key_mem_9__37_), 
        .A1N(n2030), .Y(top_core_KE_n3982) );
  OAI2BB2X1 U26045 ( .B0(n1463), .B1(n2021), .A0N(top_core_KE_key_mem_9__36_), 
        .A1N(n2031), .Y(top_core_KE_n3983) );
  OAI2BB2X1 U26046 ( .B0(n1464), .B1(n2021), .A0N(top_core_KE_key_mem_9__35_), 
        .A1N(n2031), .Y(top_core_KE_n3984) );
  OAI2BB2X1 U26047 ( .B0(n1465), .B1(n2021), .A0N(top_core_KE_key_mem_9__34_), 
        .A1N(n2031), .Y(top_core_KE_n3985) );
  OAI2BB2X1 U26048 ( .B0(n1466), .B1(n2021), .A0N(top_core_KE_key_mem_9__33_), 
        .A1N(n2031), .Y(top_core_KE_n3986) );
  OAI2BB2X1 U26049 ( .B0(n1467), .B1(n2021), .A0N(top_core_KE_key_mem_9__32_), 
        .A1N(n2031), .Y(top_core_KE_n3987) );
  OAI2BB2X1 U26050 ( .B0(n1468), .B1(n2021), .A0N(top_core_KE_key_mem_9__31_), 
        .A1N(n2031), .Y(top_core_KE_n3988) );
  OAI2BB2X1 U26051 ( .B0(n1469), .B1(n2021), .A0N(top_core_KE_key_mem_9__30_), 
        .A1N(n2031), .Y(top_core_KE_n3989) );
  OAI2BB2X1 U26052 ( .B0(n1470), .B1(n2022), .A0N(top_core_KE_key_mem_9__29_), 
        .A1N(n2031), .Y(top_core_KE_n3990) );
  OAI2BB2X1 U26053 ( .B0(n1471), .B1(n2022), .A0N(top_core_KE_key_mem_9__28_), 
        .A1N(n2031), .Y(top_core_KE_n3991) );
  OAI2BB2X1 U26054 ( .B0(n1472), .B1(n2022), .A0N(top_core_KE_key_mem_9__27_), 
        .A1N(n2031), .Y(top_core_KE_n3992) );
  OAI2BB2X1 U26055 ( .B0(n1473), .B1(n2022), .A0N(top_core_KE_key_mem_9__26_), 
        .A1N(n2031), .Y(top_core_KE_n3993) );
  OAI2BB2X1 U26056 ( .B0(n1474), .B1(n2022), .A0N(top_core_KE_key_mem_9__25_), 
        .A1N(n2031), .Y(top_core_KE_n3994) );
  OAI2BB2X1 U26057 ( .B0(n1475), .B1(n2022), .A0N(top_core_KE_key_mem_9__24_), 
        .A1N(n2031), .Y(top_core_KE_n3995) );
  OAI2BB2X1 U26058 ( .B0(n1476), .B1(n2023), .A0N(top_core_KE_key_mem_9__23_), 
        .A1N(n2031), .Y(top_core_KE_n3996) );
  OAI2BB2X1 U26059 ( .B0(n1477), .B1(n2023), .A0N(top_core_KE_key_mem_9__22_), 
        .A1N(n2031), .Y(top_core_KE_n3997) );
  OAI2BB2X1 U26060 ( .B0(n1478), .B1(n2022), .A0N(top_core_KE_key_mem_9__21_), 
        .A1N(n2032), .Y(top_core_KE_n3998) );
  OAI2BB2X1 U26061 ( .B0(n1479), .B1(n2023), .A0N(top_core_KE_key_mem_9__20_), 
        .A1N(n2032), .Y(top_core_KE_n3999) );
  OAI2BB2X1 U26062 ( .B0(n1480), .B1(n2023), .A0N(top_core_KE_key_mem_9__19_), 
        .A1N(n2032), .Y(top_core_KE_n4000) );
  OAI2BB2X1 U26063 ( .B0(n1481), .B1(n2023), .A0N(top_core_KE_key_mem_9__18_), 
        .A1N(n2032), .Y(top_core_KE_n4001) );
  OAI2BB2X1 U26064 ( .B0(n1482), .B1(n2023), .A0N(top_core_KE_key_mem_9__17_), 
        .A1N(n2032), .Y(top_core_KE_n4002) );
  OAI2BB2X1 U26065 ( .B0(n1483), .B1(n2022), .A0N(top_core_KE_key_mem_9__16_), 
        .A1N(n2032), .Y(top_core_KE_n4003) );
  OAI2BB2X1 U26066 ( .B0(n1484), .B1(n2023), .A0N(top_core_KE_key_mem_9__15_), 
        .A1N(n2032), .Y(top_core_KE_n4004) );
  OAI2BB2X1 U26067 ( .B0(n1485), .B1(n2020), .A0N(top_core_KE_key_mem_9__14_), 
        .A1N(n2032), .Y(top_core_KE_n4005) );
  OAI2BB2X1 U26068 ( .B0(n1486), .B1(n2024), .A0N(top_core_KE_key_mem_9__13_), 
        .A1N(n2032), .Y(top_core_KE_n4006) );
  OAI2BB2X1 U26069 ( .B0(n1487), .B1(n2023), .A0N(top_core_KE_key_mem_9__12_), 
        .A1N(n2032), .Y(top_core_KE_n4007) );
  OAI2BB2X1 U26070 ( .B0(n1488), .B1(n2019), .A0N(top_core_KE_key_mem_9__11_), 
        .A1N(n2032), .Y(top_core_KE_n4008) );
  OAI2BB2X1 U26071 ( .B0(n1489), .B1(n2024), .A0N(top_core_KE_key_mem_9__10_), 
        .A1N(n2032), .Y(top_core_KE_n4009) );
  OAI2BB2X1 U26072 ( .B0(n1490), .B1(n2018), .A0N(top_core_KE_key_mem_9__9_), 
        .A1N(n2032), .Y(top_core_KE_n4010) );
  OAI2BB2X1 U26073 ( .B0(n1491), .B1(n2024), .A0N(top_core_KE_key_mem_9__8_), 
        .A1N(n2032), .Y(top_core_KE_n4011) );
  OAI2BB2X1 U26074 ( .B0(n1492), .B1(n2023), .A0N(top_core_KE_key_mem_9__7_), 
        .A1N(n2032), .Y(top_core_KE_n4012) );
  OAI2BB2X1 U26075 ( .B0(n1493), .B1(n2017), .A0N(top_core_KE_key_mem_9__6_), 
        .A1N(n2020), .Y(top_core_KE_n4013) );
  OAI2BB2X1 U26076 ( .B0(n1494), .B1(n2024), .A0N(top_core_KE_key_mem_9__5_), 
        .A1N(n2021), .Y(top_core_KE_n4014) );
  OAI2BB2X1 U26077 ( .B0(n1495), .B1(n2024), .A0N(top_core_KE_key_mem_9__4_), 
        .A1N(n2022), .Y(top_core_KE_n4015) );
  OAI2BB2X1 U26078 ( .B0(n1496), .B1(n2024), .A0N(top_core_KE_key_mem_9__3_), 
        .A1N(n2028), .Y(top_core_KE_n4016) );
  OAI2BB2X1 U26079 ( .B0(n1497), .B1(n2024), .A0N(top_core_KE_key_mem_9__2_), 
        .A1N(n2029), .Y(top_core_KE_n4017) );
  OAI2BB2X1 U26080 ( .B0(n1498), .B1(n2024), .A0N(top_core_KE_key_mem_9__1_), 
        .A1N(n2027), .Y(top_core_KE_n4018) );
  OAI2BB2X1 U26081 ( .B0(n1499), .B1(n2023), .A0N(top_core_KE_key_mem_9__0_), 
        .A1N(n2027), .Y(top_core_KE_n4019) );
  OAI2BB2X1 U26082 ( .B0(n1371), .B1(n1877), .A0N(top_core_KE_key_mem_2__128_), 
        .A1N(n1888), .Y(top_core_KE_n2988) );
  OAI2BB2X1 U26083 ( .B0(n1371), .B1(n1897), .A0N(top_core_KE_key_mem_3__128_), 
        .A1N(n1907), .Y(top_core_KE_n3117) );
  OAI2BB2X1 U26084 ( .B0(n1371), .B1(n1917), .A0N(top_core_KE_key_mem_4__128_), 
        .A1N(n1928), .Y(top_core_KE_n3246) );
  OAI2BB2X1 U26085 ( .B0(n1371), .B1(n1937), .A0N(top_core_KE_key_mem_5__128_), 
        .A1N(n1947), .Y(top_core_KE_n3375) );
  OAI2BB2X1 U26086 ( .B0(n1371), .B1(n1957), .A0N(top_core_KE_key_mem_6__128_), 
        .A1N(n1968), .Y(top_core_KE_n3504) );
  OAI2BB2X1 U26087 ( .B0(n1371), .B1(n1978), .A0N(top_core_KE_key_mem_7__128_), 
        .A1N(n1987), .Y(top_core_KE_n3633) );
  OAI2BB2X1 U26088 ( .B0(n1371), .B1(n2037), .A0N(top_core_KE_key_mem_10__128_), .A1N(n2048), .Y(top_core_KE_n4020) );
  OAI2BB2X1 U26089 ( .B0(n1371), .B1(n2058), .A0N(top_core_KE_key_mem_11__128_), .A1N(n2067), .Y(top_core_KE_n4149) );
  OAI2BB2X1 U26090 ( .B0(n1371), .B1(n2077), .A0N(top_core_KE_key_mem_12__128_), .A1N(n2087), .Y(top_core_KE_n4278) );
  OAI2BB2X1 U26091 ( .B0(n1371), .B1(n2098), .A0N(top_core_KE_key_mem_13__128_), .A1N(n2107), .Y(top_core_KE_n4407) );
  OAI2BB2X1 U26092 ( .B0(n1371), .B1(n2118), .A0N(top_core_KE_key_mem_14__128_), .A1N(n2127), .Y(top_core_KE_n4536) );
  OAI2BB2X1 U26093 ( .B0(n1371), .B1(n1861), .A0N(top_core_KE_key_mem_1__128_), 
        .A1N(n1866), .Y(top_core_KE_n2859) );
  OAI2BB2X1 U26094 ( .B0(n1371), .B1(n1997), .A0N(top_core_KE_key_mem_8__128_), 
        .A1N(n2007), .Y(top_core_KE_n3762) );
  OAI2BB2X1 U26095 ( .B0(n1371), .B1(n2026), .A0N(top_core_KE_key_mem_9__128_), 
        .A1N(n2027), .Y(top_core_KE_n3891) );
  AND2X2 U26096 ( .A(n3570), .B(top_core_Core_Full), .Y(top_core_EC_n1009) );
  INVX1 U26097 ( .A(top_core_KE_rcon_reg_3_), .Y(n7002) );
  INVX1 U26098 ( .A(top_core_KE_rcon_reg_2_), .Y(n7003) );
  INVX1 U26099 ( .A(top_core_KE_rcon_reg_0_), .Y(n7005) );
  INVX1 U26100 ( .A(top_core_KE_prev_key0_reg_62_), .Y(n6405) );
  INVX1 U26101 ( .A(top_core_KE_prev_key0_reg_61_), .Y(n6513) );
  INVX1 U26102 ( .A(top_core_KE_prev_key0_reg_60_), .Y(n6583) );
  INVX1 U26103 ( .A(top_core_KE_prev_key0_reg_59_), .Y(n6647) );
  INVX1 U26104 ( .A(top_core_KE_prev_key0_reg_58_), .Y(n6671) );
  INVX1 U26105 ( .A(top_core_KE_prev_key0_reg_57_), .Y(n6310) );
  INVX1 U26106 ( .A(top_core_KE_prev_key0_reg_56_), .Y(n6692) );
  INVX1 U26107 ( .A(top_core_KE_prev_key0_reg_55_), .Y(n6332) );
  INVX1 U26108 ( .A(top_core_KE_prev_key0_reg_54_), .Y(n6396) );
  INVX1 U26109 ( .A(top_core_KE_prev_key0_reg_53_), .Y(n6444) );
  INVX1 U26110 ( .A(top_core_KE_prev_key0_reg_52_), .Y(n6535) );
  INVX1 U26111 ( .A(top_core_KE_prev_key0_reg_51_), .Y(n6630) );
  INVX1 U26112 ( .A(top_core_KE_prev_key0_reg_50_), .Y(n6663) );
  INVX1 U26113 ( .A(top_core_KE_prev_key0_reg_49_), .Y(n6678) );
  INVX1 U26114 ( .A(top_core_KE_prev_key0_reg_48_), .Y(n6685) );
  INVX1 U26115 ( .A(top_core_KE_prev_key0_reg_47_), .Y(n6323) );
  INVX1 U26116 ( .A(top_core_KE_prev_key0_reg_46_), .Y(n6388) );
  INVX1 U26117 ( .A(top_core_KE_prev_key0_reg_45_), .Y(n6810) );
  INVX1 U26118 ( .A(top_core_KE_prev_key0_reg_44_), .Y(n6877) );
  INVX1 U26119 ( .A(top_core_KE_prev_key0_reg_43_), .Y(n6938) );
  INVX1 U26120 ( .A(top_core_KE_prev_key0_reg_42_), .Y(n6959) );
  INVX1 U26121 ( .A(top_core_KE_prev_key0_reg_34_), .Y(n6953) );
  INVX1 U26122 ( .A(top_core_KE_prev_key0_reg_33_), .Y(n6965) );
  INVX1 U26123 ( .A(top_core_KE_prev_key0_reg_32_), .Y(n6975) );
  XNOR2X1 U26124 ( .A(top_core_KE_n2515), .B(top_core_KE_n2350), .Y(
        top_core_KE_n1369) );
  XNOR2X1 U26125 ( .A(top_core_KE_prev_key1_reg_62_), .B(n6484), .Y(
        top_core_KE_n2515) );
  XNOR2X1 U26126 ( .A(top_core_KE_n2518), .B(top_core_KE_n2356), .Y(
        top_core_KE_n1377) );
  XNOR2X1 U26127 ( .A(top_core_KE_prev_key1_reg_61_), .B(n6485), .Y(
        top_core_KE_n2518) );
  XNOR2X1 U26128 ( .A(top_core_KE_n2521), .B(top_core_KE_n2362), .Y(
        top_core_KE_n1385) );
  XNOR2X1 U26129 ( .A(top_core_KE_prev_key1_reg_60_), .B(n6486), .Y(
        top_core_KE_n2521) );
  XNOR2X1 U26130 ( .A(top_core_KE_n2524), .B(top_core_KE_n2368), .Y(
        top_core_KE_n1393) );
  XNOR2X1 U26131 ( .A(top_core_KE_prev_key1_reg_59_), .B(n6489), .Y(
        top_core_KE_n2524) );
  XNOR2X1 U26132 ( .A(top_core_KE_n2527), .B(top_core_KE_n2374), .Y(
        top_core_KE_n1401) );
  XNOR2X1 U26133 ( .A(top_core_KE_prev_key1_reg_58_), .B(n6492), .Y(
        top_core_KE_n2527) );
  XNOR2X1 U26134 ( .A(top_core_KE_n2530), .B(top_core_KE_n2380), .Y(
        top_core_KE_n1409) );
  XNOR2X1 U26135 ( .A(top_core_KE_prev_key1_reg_57_), .B(n6496), .Y(
        top_core_KE_n2530) );
  XNOR2X1 U26136 ( .A(top_core_KE_n2533), .B(top_core_KE_n2386), .Y(
        top_core_KE_n1417) );
  XNOR2X1 U26137 ( .A(top_core_KE_prev_key1_reg_56_), .B(n6499), .Y(
        top_core_KE_n2533) );
  XNOR2X1 U26138 ( .A(top_core_KE_n2560), .B(top_core_KE_n2561), .Y(
        top_core_KE_n1617) );
  XNOR2X1 U26139 ( .A(n1370), .B(top_core_KE_prev_key1_reg_63_), .Y(
        top_core_KE_n2560) );
  XNOR2X1 U26140 ( .A(top_core_KE_n2183), .B(top_core_KE_n2344), .Y(
        top_core_KE_n2561) );
  XNOR2X1 U26141 ( .A(top_core_KE_n2565), .B(top_core_KE_n2566), .Y(
        top_core_KE_n1625) );
  XNOR2X1 U26142 ( .A(n1368), .B(top_core_KE_prev_key1_reg_62_), .Y(
        top_core_KE_n2565) );
  XNOR2X1 U26143 ( .A(top_core_KE_n2514), .B(top_core_KE_n2350), .Y(
        top_core_KE_n2566) );
  XNOR2X1 U26144 ( .A(top_core_KE_n2570), .B(top_core_KE_n2571), .Y(
        top_core_KE_n1633) );
  XNOR2X1 U26145 ( .A(n1754), .B(top_core_KE_prev_key1_reg_61_), .Y(
        top_core_KE_n2570) );
  XNOR2X1 U26146 ( .A(top_core_KE_n2517), .B(top_core_KE_n2356), .Y(
        top_core_KE_n2571) );
  XNOR2X1 U26147 ( .A(top_core_KE_n2575), .B(top_core_KE_n2576), .Y(
        top_core_KE_n1641) );
  XNOR2X1 U26148 ( .A(n1364), .B(top_core_KE_prev_key1_reg_60_), .Y(
        top_core_KE_n2575) );
  XNOR2X1 U26149 ( .A(top_core_KE_n2520), .B(top_core_KE_n2362), .Y(
        top_core_KE_n2576) );
  XNOR2X1 U26150 ( .A(top_core_KE_n2580), .B(top_core_KE_n2581), .Y(
        top_core_KE_n1649) );
  XNOR2X1 U26151 ( .A(n1360), .B(top_core_KE_prev_key1_reg_59_), .Y(
        top_core_KE_n2580) );
  XNOR2X1 U26152 ( .A(top_core_KE_n2523), .B(top_core_KE_n2368), .Y(
        top_core_KE_n2581) );
  XNOR2X1 U26153 ( .A(top_core_KE_n2585), .B(top_core_KE_n2586), .Y(
        top_core_KE_n1657) );
  XNOR2X1 U26154 ( .A(n1358), .B(top_core_KE_prev_key1_reg_58_), .Y(
        top_core_KE_n2585) );
  XNOR2X1 U26155 ( .A(top_core_KE_n2526), .B(top_core_KE_n2374), .Y(
        top_core_KE_n2586) );
  XNOR2X1 U26156 ( .A(top_core_KE_n2590), .B(top_core_KE_n2591), .Y(
        top_core_KE_n1665) );
  XNOR2X1 U26157 ( .A(n1760), .B(top_core_KE_prev_key1_reg_57_), .Y(
        top_core_KE_n2590) );
  XNOR2X1 U26158 ( .A(top_core_KE_n2529), .B(top_core_KE_n2380), .Y(
        top_core_KE_n2591) );
  XNOR2X1 U26159 ( .A(top_core_KE_n2595), .B(top_core_KE_n2596), .Y(
        top_core_KE_n1673) );
  XNOR2X1 U26160 ( .A(n1767), .B(top_core_KE_prev_key1_reg_56_), .Y(
        top_core_KE_n2595) );
  XNOR2X1 U26161 ( .A(top_core_KE_n2532), .B(top_core_KE_n2386), .Y(
        top_core_KE_n2596) );
  OAI2BB2XL U26163 ( .B0(n4196), .B1(n2), .A0N(n2), .A1N(top_core_EC_rounds_2_), .Y(top_core_EC_n1297) );
  OAI2BB2XL U26164 ( .B0(n4197), .B1(n2), .A0N(n2), .A1N(top_core_EC_rounds_3_), .Y(top_core_EC_n1298) );
  INVX1 U26165 ( .A(top_core_KE_prev_key0_reg_41_), .Y(n6970) );
  INVX1 U26166 ( .A(top_core_KE_prev_key0_reg_40_), .Y(n6980) );
  INVX1 U26167 ( .A(top_core_KE_prev_key0_reg_39_), .Y(n6319) );
  INVX1 U26168 ( .A(top_core_KE_prev_key0_reg_38_), .Y(n6380) );
  INVX1 U26169 ( .A(top_core_KE_prev_key0_reg_37_), .Y(n6747) );
  INVX1 U26170 ( .A(top_core_KE_prev_key0_reg_36_), .Y(n6831) );
  INVX1 U26171 ( .A(top_core_KE_prev_key0_reg_35_), .Y(n6923) );
  BUFX3 U26172 ( .A(top_core_KE_prev_key1_reg_75_), .Y(n1347) );
  BUFX3 U26173 ( .A(top_core_KE_prev_key1_reg_67_), .Y(n1349) );
  BUFX3 U26174 ( .A(top_core_KE_prev_key1_reg_83_), .Y(n1363) );
  AOI2BB2X1 U26175 ( .B0(top_core_KE_CipherKey0_63_), .B1(n2217), .A0N(n2190), 
        .A1N(top_core_KE_n1358), .Y(top_core_KE_n1357) );
  INVX1 U26176 ( .A(top_core_EC_round_result_r_1_), .Y(n6303) );
  INVX1 U26177 ( .A(top_core_EC_round_result_r_18_), .Y(n6286) );
  INVX1 U26178 ( .A(top_core_EC_round_result_r_2_), .Y(n6302) );
  INVX1 U26179 ( .A(top_core_EC_round_result_r_34_), .Y(n6270) );
  INVX1 U26180 ( .A(top_core_EC_round_result_r_50_), .Y(n6254) );
  INVX1 U26181 ( .A(top_core_EC_round_result_r_16_), .Y(n6288) );
  INVX1 U26182 ( .A(top_core_EC_round_result_r_0_), .Y(n6304) );
  INVX1 U26183 ( .A(top_core_EC_round_result_r_19_), .Y(n6285) );
  INVX1 U26184 ( .A(top_core_EC_round_result_r_3_), .Y(n6301) );
  INVX1 U26185 ( .A(top_core_EC_round_result_r_7_), .Y(n6297) );
  INVX1 U26186 ( .A(top_core_EC_round_result_r_32_), .Y(n6272) );
  INVX1 U26187 ( .A(top_core_EC_round_result_r_48_), .Y(n6256) );
  INVX1 U26188 ( .A(top_core_EC_round_result_r_51_), .Y(n6253) );
  INVX1 U26189 ( .A(top_core_EC_round_result_r_35_), .Y(n6269) );
  INVX1 U26190 ( .A(top_core_EC_round_result_r_17_), .Y(n6287) );
  INVX1 U26191 ( .A(top_core_EC_round_result_r_10_), .Y(n6294) );
  INVX1 U26192 ( .A(top_core_EC_round_result_r_11_), .Y(n6293) );
  INVX1 U26193 ( .A(top_core_EC_round_result_r_20_), .Y(n6284) );
  INVX1 U26194 ( .A(top_core_EC_round_result_r_4_), .Y(n6300) );
  INVX1 U26195 ( .A(top_core_EC_round_result_r_21_), .Y(n6283) );
  INVX1 U26196 ( .A(top_core_EC_round_result_r_5_), .Y(n6299) );
  INVX1 U26197 ( .A(top_core_EC_round_result_r_22_), .Y(n6282) );
  INVX1 U26198 ( .A(top_core_EC_round_result_r_6_), .Y(n6298) );
  INVX1 U26199 ( .A(top_core_EC_round_result_r_23_), .Y(n6281) );
  INVX1 U26200 ( .A(top_core_EC_round_result_r_49_), .Y(n6255) );
  INVX1 U26201 ( .A(top_core_EC_round_result_r_33_), .Y(n6271) );
  INVX1 U26202 ( .A(top_core_EC_round_result_r_52_), .Y(n6252) );
  INVX1 U26203 ( .A(top_core_EC_round_result_r_53_), .Y(n6251) );
  INVX1 U26204 ( .A(top_core_EC_round_result_r_36_), .Y(n6268) );
  INVX1 U26205 ( .A(top_core_EC_round_result_r_54_), .Y(n6250) );
  INVX1 U26206 ( .A(top_core_EC_round_result_r_37_), .Y(n6267) );
  INVX1 U26207 ( .A(top_core_EC_round_result_r_55_), .Y(n6249) );
  INVX1 U26208 ( .A(top_core_EC_round_result_r_39_), .Y(n6265) );
  INVX1 U26209 ( .A(top_core_EC_round_result_r_38_), .Y(n6266) );
  INVX1 U26210 ( .A(top_core_EC_round_result_r_8_), .Y(n6296) );
  INVX1 U26211 ( .A(top_core_EC_round_result_r_13_), .Y(n6291) );
  INVX1 U26212 ( .A(top_core_EC_round_result_r_14_), .Y(n6290) );
  INVX1 U26213 ( .A(top_core_EC_round_result_r_29_), .Y(n6275) );
  INVX1 U26214 ( .A(top_core_EC_round_result_r_30_), .Y(n6274) );
  INVX1 U26215 ( .A(top_core_EC_round_result_r_40_), .Y(n6264) );
  INVX1 U26216 ( .A(top_core_EC_round_result_r_42_), .Y(n6262) );
  INVX1 U26217 ( .A(top_core_EC_round_result_r_43_), .Y(n6261) );
  INVX1 U26218 ( .A(top_core_EC_round_result_r_45_), .Y(n6259) );
  INVX1 U26219 ( .A(top_core_EC_round_result_r_46_), .Y(n6258) );
  INVX1 U26220 ( .A(top_core_EC_round_result_r_47_), .Y(n6257) );
  INVX1 U26221 ( .A(top_core_EC_round_result_r_15_), .Y(n6289) );
  INVX1 U26222 ( .A(top_core_EC_round_result_r_31_), .Y(n6273) );
  INVX1 U26223 ( .A(top_core_EC_round_result_r_24_), .Y(n6280) );
  INVX1 U26224 ( .A(top_core_EC_round_result_r_26_), .Y(n6278) );
  INVX1 U26225 ( .A(top_core_EC_round_result_r_27_), .Y(n6277) );
  INVX1 U26226 ( .A(top_core_EC_round_result_r_9_), .Y(n6295) );
  INVX1 U26227 ( .A(top_core_EC_round_result_r_12_), .Y(n6292) );
  INVX1 U26228 ( .A(top_core_EC_round_result_r_25_), .Y(n6279) );
  INVX1 U26229 ( .A(top_core_EC_round_result_r_28_), .Y(n6276) );
  INVX1 U26230 ( .A(top_core_EC_round_result_r_56_), .Y(n6248) );
  INVX1 U26231 ( .A(top_core_EC_round_result_r_41_), .Y(n6263) );
  INVX1 U26232 ( .A(top_core_EC_round_result_r_44_), .Y(n6260) );
  INVX1 U26233 ( .A(top_core_EC_round_result_r_57_), .Y(n6247) );
  BUFX3 U26234 ( .A(top_core_KE_prev_key1_reg_31_), .Y(n1370) );
  BUFX3 U26235 ( .A(top_core_KE_prev_key1_reg_91_), .Y(n1361) );
  INVX1 U26236 ( .A(top_core_EC_round_result_r_81_), .Y(n6223) );
  INVX1 U26237 ( .A(top_core_EC_round_result_r_113_), .Y(n6191) );
  INVX1 U26238 ( .A(top_core_EC_round_result_r_80_), .Y(n6224) );
  INVX1 U26239 ( .A(top_core_EC_round_result_r_74_), .Y(n6230) );
  INVX1 U26240 ( .A(top_core_EC_round_result_r_112_), .Y(n6192) );
  INVX1 U26241 ( .A(top_core_EC_round_result_r_122_), .Y(n6182) );
  INVX1 U26242 ( .A(top_core_EC_round_result_r_82_), .Y(n6222) );
  INVX1 U26243 ( .A(top_core_EC_round_result_r_114_), .Y(n6190) );
  INVX1 U26244 ( .A(top_core_EC_round_result_r_89_), .Y(n6215) );
  INVX1 U26245 ( .A(top_core_EC_round_result_r_66_), .Y(n6238) );
  INVX1 U26246 ( .A(top_core_EC_round_result_r_65_), .Y(n6239) );
  INVX1 U26247 ( .A(top_core_EC_round_result_r_121_), .Y(n6183) );
  INVX1 U26248 ( .A(top_core_EC_round_result_r_98_), .Y(n6206) );
  INVX1 U26249 ( .A(top_core_EC_round_result_r_97_), .Y(n6207) );
  INVX1 U26250 ( .A(top_core_EC_round_result_r_90_), .Y(n6214) );
  INVX1 U26251 ( .A(top_core_EC_round_result_r_104_), .Y(n6200) );
  INVX1 U26252 ( .A(top_core_EC_round_result_r_105_), .Y(n6199) );
  INVX1 U26253 ( .A(top_core_EC_round_result_r_85_), .Y(n6219) );
  INVX1 U26254 ( .A(top_core_EC_round_result_r_84_), .Y(n6220) );
  INVX1 U26255 ( .A(top_core_EC_round_result_r_120_), .Y(n6184) );
  INVX1 U26256 ( .A(top_core_EC_round_result_r_72_), .Y(n6232) );
  INVX1 U26257 ( .A(top_core_EC_round_result_r_73_), .Y(n6231) );
  INVX1 U26258 ( .A(top_core_EC_round_result_r_117_), .Y(n6187) );
  INVX1 U26259 ( .A(top_core_EC_round_result_r_116_), .Y(n6188) );
  INVX1 U26260 ( .A(top_core_EC_round_result_r_64_), .Y(n6240) );
  INVX1 U26261 ( .A(top_core_EC_round_result_r_96_), .Y(n6208) );
  INVX1 U26262 ( .A(top_core_EC_round_result_r_88_), .Y(n6216) );
  INVX1 U26263 ( .A(top_core_EC_round_result_r_106_), .Y(n6198) );
  INVX1 U26264 ( .A(top_core_EC_round_result_r_58_), .Y(n6246) );
  INVX1 U26265 ( .A(top_core_EC_round_result_r_124_), .Y(n6180) );
  INVX1 U26266 ( .A(top_core_EC_round_result_r_77_), .Y(n6227) );
  INVX1 U26267 ( .A(top_core_EC_round_result_r_76_), .Y(n6228) );
  INVX1 U26268 ( .A(top_core_EC_round_result_r_125_), .Y(n6179) );
  INVX1 U26269 ( .A(top_core_EC_round_result_r_109_), .Y(n6195) );
  INVX1 U26270 ( .A(top_core_EC_round_result_r_108_), .Y(n6196) );
  INVX1 U26271 ( .A(top_core_EC_round_result_r_86_), .Y(n6218) );
  INVX1 U26272 ( .A(top_core_EC_round_result_r_61_), .Y(n6243) );
  INVX1 U26273 ( .A(top_core_EC_round_result_r_118_), .Y(n6186) );
  INVX1 U26274 ( .A(top_core_EC_round_result_r_68_), .Y(n6236) );
  INVX1 U26275 ( .A(top_core_EC_round_result_r_69_), .Y(n6235) );
  INVX1 U26276 ( .A(top_core_EC_round_result_r_100_), .Y(n6204) );
  INVX1 U26277 ( .A(top_core_EC_round_result_r_101_), .Y(n6203) );
  INVX1 U26278 ( .A(top_core_EC_round_result_r_92_), .Y(n6212) );
  INVX1 U26279 ( .A(top_core_EC_round_result_r_60_), .Y(n6244) );
  INVX1 U26280 ( .A(top_core_EC_round_result_r_93_), .Y(n6211) );
  INVX1 U26281 ( .A(top_core_EC_round_result_r_78_), .Y(n6226) );
  INVX1 U26282 ( .A(top_core_EC_round_result_r_110_), .Y(n6194) );
  INVX1 U26283 ( .A(top_core_EC_round_result_r_83_), .Y(n6221) );
  INVX1 U26284 ( .A(top_core_EC_round_result_r_62_), .Y(n6242) );
  INVX1 U26285 ( .A(top_core_EC_round_result_r_126_), .Y(n6178) );
  INVX1 U26286 ( .A(top_core_EC_round_result_r_115_), .Y(n6189) );
  INVX1 U26287 ( .A(top_core_EC_round_result_r_70_), .Y(n6234) );
  INVX1 U26288 ( .A(top_core_EC_round_result_r_102_), .Y(n6202) );
  INVX1 U26289 ( .A(top_core_EC_round_result_r_94_), .Y(n6210) );
  INVX1 U26290 ( .A(top_core_EC_round_result_r_75_), .Y(n6229) );
  INVX1 U26291 ( .A(top_core_EC_round_result_r_123_), .Y(n6181) );
  INVX1 U26292 ( .A(top_core_EC_round_result_r_67_), .Y(n6237) );
  INVX1 U26293 ( .A(top_core_EC_round_result_r_107_), .Y(n6197) );
  INVX1 U26294 ( .A(top_core_EC_round_result_r_59_), .Y(n6245) );
  INVX1 U26295 ( .A(top_core_EC_round_result_r_99_), .Y(n6205) );
  INVX1 U26296 ( .A(top_core_EC_round_result_r_91_), .Y(n6213) );
  INVX1 U26297 ( .A(top_core_EC_round_result_r_87_), .Y(n6217) );
  INVX1 U26298 ( .A(top_core_EC_round_result_r_119_), .Y(n6185) );
  INVX1 U26299 ( .A(top_core_EC_round_result_r_71_), .Y(n6233) );
  INVX1 U26300 ( .A(top_core_EC_round_result_r_111_), .Y(n6193) );
  INVX1 U26301 ( .A(top_core_EC_round_result_r_63_), .Y(n6241) );
  INVX1 U26302 ( .A(top_core_EC_round_result_r_127_), .Y(n6177) );
  INVX1 U26303 ( .A(top_core_EC_round_result_r_103_), .Y(n6201) );
  INVX1 U26304 ( .A(top_core_EC_round_result_r_79_), .Y(n6225) );
  INVX1 U26305 ( .A(top_core_EC_round_result_r_95_), .Y(n6209) );
  BUFX3 U26306 ( .A(top_core_KE_round_ctr_reg_3_), .Y(n1334) );
  BUFX3 U26307 ( .A(top_core_KE_prev_key1_reg_15_), .Y(n1338) );
  BUFX3 U26308 ( .A(top_core_KE_prev_key1_reg_7_), .Y(n1335) );
  BUFX3 U26309 ( .A(top_core_KE_prev_key1_reg_23_), .Y(n1339) );
  INVX1 U26310 ( .A(top_core_KE_prev_key0_reg_9_), .Y(n6974) );
  INVX1 U26311 ( .A(top_core_KE_prev_key0_reg_8_), .Y(n6984) );
  INVX1 U26312 ( .A(top_core_KE_prev_key0_reg_7_), .Y(n6996) );
  INVX1 U26313 ( .A(top_core_KE_prev_key0_reg_6_), .Y(n6387) );
  INVX1 U26314 ( .A(top_core_KE_prev_key0_reg_5_), .Y(n6784) );
  INVX1 U26315 ( .A(top_core_KE_prev_key0_reg_4_), .Y(n6856) );
  INVX1 U26316 ( .A(top_core_KE_prev_key0_reg_3_), .Y(n6932) );
  INVX1 U26317 ( .A(top_core_KE_prev_key0_reg_31_), .Y(n6345) );
  INVX1 U26318 ( .A(top_core_KE_prev_key0_reg_30_), .Y(n6438) );
  INVX1 U26319 ( .A(top_core_KE_prev_key0_reg_29_), .Y(n6526) );
  INVX1 U26320 ( .A(top_core_KE_prev_key0_reg_28_), .Y(n6609) );
  INVX1 U26321 ( .A(top_core_KE_prev_key0_reg_27_), .Y(n6657) );
  INVX1 U26322 ( .A(top_core_KE_prev_key0_reg_26_), .Y(n6676) );
  INVX1 U26323 ( .A(top_core_KE_prev_key0_reg_25_), .Y(n6318) );
  INVX1 U26324 ( .A(top_core_KE_prev_key0_reg_24_), .Y(n6697) );
  INVX1 U26325 ( .A(top_core_KE_prev_key0_reg_23_), .Y(n6991) );
  INVX1 U26326 ( .A(top_core_KE_prev_key0_reg_22_), .Y(n6404) );
  INVX1 U26327 ( .A(top_core_KE_prev_key0_reg_21_), .Y(n6482) );
  INVX1 U26328 ( .A(top_core_KE_prev_key0_reg_20_), .Y(n6562) );
  INVX1 U26329 ( .A(top_core_KE_prev_key0_reg_19_), .Y(n6641) );
  INVX1 U26330 ( .A(top_core_KE_prev_key0_reg_18_), .Y(n6669) );
  INVX1 U26331 ( .A(top_core_KE_prev_key0_reg_17_), .Y(n6684) );
  INVX1 U26332 ( .A(top_core_KE_prev_key0_reg_16_), .Y(n6691) );
  INVX1 U26333 ( .A(top_core_KE_prev_key0_reg_15_), .Y(n6331) );
  INVX1 U26334 ( .A(top_core_KE_prev_key0_reg_14_), .Y(n6720) );
  INVX1 U26335 ( .A(top_core_KE_prev_key0_reg_13_), .Y(n6822) );
  INVX1 U26336 ( .A(top_core_KE_prev_key0_reg_12_), .Y(n6902) );
  INVX1 U26337 ( .A(top_core_KE_prev_key0_reg_11_), .Y(n6947) );
  INVX1 U26338 ( .A(top_core_KE_prev_key0_reg_10_), .Y(n6963) );
  INVX1 U26339 ( .A(top_core_KE_prev_key0_reg_2_), .Y(n6957) );
  INVX1 U26340 ( .A(top_core_KE_prev_key0_reg_1_), .Y(n6969) );
  INVX1 U26341 ( .A(top_core_KE_prev_key0_reg_0_), .Y(n6979) );
  NAND3X1 U26342 ( .A(top_core_KE_n2375), .B(top_core_KE_n2376), .C(
        top_core_KE_n2377), .Y(top_core_KE_n4830) );
  AOI222X1 U26343 ( .A0(n1652), .A1(n2299), .B0(n2309), .B1(
        top_core_KE_CipherKey0_25_), .C0(n2355), .C1(n6312), .Y(
        top_core_KE_n2377) );
  AOI22X1 U26344 ( .A0(top_core_KE_n2181), .A1(top_core_KE_n1177), .B0(n2338), 
        .B1(top_core_KE_n1179), .Y(top_core_KE_n2375) );
  AOI22X1 U26345 ( .A0(n2314), .A1(top_core_KE_n2378), .B0(n2319), .B1(
        top_core_KE_CipherKey0_89_), .Y(top_core_KE_n2376) );
  NAND3X1 U26346 ( .A(top_core_KE_n2467), .B(top_core_KE_n2468), .C(
        top_core_KE_n2469), .Y(top_core_KE_n4848) );
  AOI222X1 U26347 ( .A0(n1336), .A1(n2303), .B0(n2307), .B1(
        top_core_KE_CipherKey0_7_), .C0(n2351), .C1(top_core_KE_n1301), .Y(
        top_core_KE_n2469) );
  AOI22X1 U26348 ( .A0(n2329), .A1(top_core_KE_n1303), .B0(n2339), .B1(
        top_core_KE_n1305), .Y(top_core_KE_n2467) );
  AOI22X1 U26349 ( .A0(n2312), .A1(top_core_KE_n2470), .B0(n2320), .B1(
        top_core_KE_CipherKey0_71_), .Y(top_core_KE_n2468) );
  NAND3X1 U26350 ( .A(top_core_KE_n2427), .B(top_core_KE_n2428), .C(
        top_core_KE_n2429), .Y(top_core_KE_n4840) );
  AOI222X1 U26351 ( .A0(n1337), .A1(n2303), .B0(n2308), .B1(
        top_core_KE_CipherKey0_15_), .C0(n2354), .C1(top_core_KE_n1245), .Y(
        top_core_KE_n2429) );
  AOI22X1 U26352 ( .A0(n2329), .A1(top_core_KE_n1247), .B0(n2339), .B1(
        top_core_KE_n1249), .Y(top_core_KE_n2427) );
  AOI22X1 U26353 ( .A0(n2313), .A1(top_core_KE_n2430), .B0(n2320), .B1(
        top_core_KE_CipherKey0_79_), .Y(top_core_KE_n2428) );
  NAND3X1 U26354 ( .A(top_core_KE_n2387), .B(top_core_KE_n2388), .C(
        top_core_KE_n2389), .Y(top_core_KE_n4832) );
  AOI222X1 U26355 ( .A0(n1340), .A1(n2300), .B0(n2308), .B1(
        top_core_KE_CipherKey0_23_), .C0(n2362), .C1(top_core_KE_n1189), .Y(
        top_core_KE_n2389) );
  AOI22X1 U26356 ( .A0(top_core_KE_n2181), .A1(top_core_KE_n1191), .B0(n2337), 
        .B1(top_core_KE_n1193), .Y(top_core_KE_n2387) );
  AOI22X1 U26357 ( .A0(n2313), .A1(top_core_KE_n2390), .B0(n2319), .B1(
        top_core_KE_CipherKey0_87_), .Y(top_core_KE_n2388) );
  NAND3X1 U26358 ( .A(top_core_KE_n2339), .B(top_core_KE_n2340), .C(
        top_core_KE_n2341), .Y(top_core_KE_n4824) );
  AOI222X1 U26359 ( .A0(n1341), .A1(n2297), .B0(n2309), .B1(
        top_core_KE_CipherKey0_31_), .C0(n2357), .C1(n6339), .Y(
        top_core_KE_n2341) );
  AOI22X1 U26360 ( .A0(n2328), .A1(top_core_KE_n1135), .B0(n2338), .B1(
        top_core_KE_n1137), .Y(top_core_KE_n2339) );
  AOI22X1 U26361 ( .A0(n2314), .A1(top_core_KE_n2342), .B0(n2318), .B1(
        top_core_KE_CipherKey0_95_), .Y(top_core_KE_n2340) );
  NAND3X1 U26362 ( .A(top_core_KE_n2472), .B(top_core_KE_n2473), .C(
        top_core_KE_n2474), .Y(top_core_KE_n4849) );
  AOI222X1 U26363 ( .A0(n1342), .A1(n2292), .B0(n2307), .B1(
        top_core_KE_CipherKey0_6_), .C0(n2351), .C1(top_core_KE_n1308), .Y(
        top_core_KE_n2474) );
  AOI22X1 U26364 ( .A0(n2329), .A1(top_core_KE_n1310), .B0(n2339), .B1(
        top_core_KE_n1312), .Y(top_core_KE_n2472) );
  AOI22X1 U26365 ( .A0(n2312), .A1(top_core_KE_n2475), .B0(n2320), .B1(
        top_core_KE_CipherKey0_70_), .Y(top_core_KE_n2473) );
  NAND3X1 U26366 ( .A(top_core_KE_n2294), .B(top_core_KE_n2295), .C(
        top_core_KE_n2296), .Y(top_core_KE_n4815) );
  AOI222X1 U26367 ( .A0(top_core_KE_prev_key1_reg_104_), .A1(n2301), .B0(
        top_core_KE_n2176), .B1(top_core_KE_CipherKey0_40_), .C0(n767), .C1(
        n6741), .Y(top_core_KE_n2296) );
  AOI22X1 U26368 ( .A0(n2312), .A1(top_core_KE_n2297), .B0(top_core_KE_n2179), 
        .B1(top_core_KE_CipherKey0_104_), .Y(top_core_KE_n2295) );
  AOI22X1 U26369 ( .A0(n2327), .A1(top_core_KE_n1072), .B0(n2337), .B1(
        top_core_KE_n1074), .Y(top_core_KE_n2294) );
  NAND3X1 U26370 ( .A(top_core_KE_n2462), .B(top_core_KE_n2463), .C(
        top_core_KE_n2464), .Y(top_core_KE_n4847) );
  AOI222X1 U26371 ( .A0(n1717), .A1(n2302), .B0(n2307), .B1(
        top_core_KE_CipherKey0_8_), .C0(n2351), .C1(top_core_KE_n1294), .Y(
        top_core_KE_n2464) );
  AOI22X1 U26372 ( .A0(n2329), .A1(top_core_KE_n1296), .B0(n2339), .B1(
        top_core_KE_n1298), .Y(top_core_KE_n2462) );
  AOI22X1 U26373 ( .A0(n2312), .A1(top_core_KE_n2465), .B0(n2320), .B1(
        top_core_KE_CipherKey0_72_), .Y(top_core_KE_n2463) );
  NAND3X1 U26374 ( .A(top_core_KE_n2334), .B(top_core_KE_n2335), .C(
        top_core_KE_n2336), .Y(top_core_KE_n4823) );
  AOI222X1 U26375 ( .A0(top_core_KE_prev_key1_reg_96_), .A1(n2299), .B0(n2309), 
        .B1(top_core_KE_CipherKey0_32_), .C0(n2357), .C1(n6798), .Y(
        top_core_KE_n2336) );
  AOI22X1 U26376 ( .A0(n2314), .A1(top_core_KE_n2337), .B0(n2318), .B1(
        top_core_KE_CipherKey0_96_), .Y(top_core_KE_n2335) );
  AOI22X1 U26377 ( .A0(n2328), .A1(top_core_KE_n1128), .B0(n2338), .B1(
        top_core_KE_n1130), .Y(top_core_KE_n2334) );
  NAND3X1 U26378 ( .A(top_core_KE_n2502), .B(top_core_KE_n2503), .C(
        top_core_KE_n2504), .Y(top_core_KE_n4855) );
  AOI222X1 U26379 ( .A0(n1746), .A1(n2284), .B0(n2307), .B1(
        top_core_KE_CipherKey0_0_), .C0(n2360), .C1(top_core_KE_n1350), .Y(
        top_core_KE_n2504) );
  AOI22X1 U26380 ( .A0(n2330), .A1(top_core_KE_n1352), .B0(n2340), .B1(
        top_core_KE_n1354), .Y(top_core_KE_n2502) );
  AOI22X1 U26381 ( .A0(n2312), .A1(top_core_KE_n2507), .B0(n2321), .B1(
        top_core_KE_CipherKey0_64_), .Y(top_core_KE_n2503) );
  NAND3X1 U26382 ( .A(top_core_KE_n2289), .B(top_core_KE_n2290), .C(
        top_core_KE_n2291), .Y(top_core_KE_n4814) );
  AOI222X1 U26383 ( .A0(top_core_KE_prev_key1_reg_105_), .A1(n2299), .B0(
        top_core_KE_n2176), .B1(top_core_KE_CipherKey0_41_), .C0(n767), .C1(
        n6738), .Y(top_core_KE_n2291) );
  AOI22X1 U26384 ( .A0(n2313), .A1(top_core_KE_n2292), .B0(top_core_KE_n2179), 
        .B1(top_core_KE_CipherKey0_105_), .Y(top_core_KE_n2290) );
  AOI22X1 U26385 ( .A0(n2327), .A1(top_core_KE_n1065), .B0(n2337), .B1(
        top_core_KE_n1067), .Y(top_core_KE_n2289) );
  NAND3X1 U26386 ( .A(top_core_KE_n2457), .B(top_core_KE_n2458), .C(
        top_core_KE_n2459), .Y(top_core_KE_n4846) );
  AOI222X1 U26387 ( .A0(n1710), .A1(n2293), .B0(n2307), .B1(
        top_core_KE_CipherKey0_9_), .C0(n2352), .C1(top_core_KE_n1287), .Y(
        top_core_KE_n2459) );
  AOI22X1 U26388 ( .A0(n2329), .A1(top_core_KE_n1289), .B0(n2339), .B1(
        top_core_KE_n1291), .Y(top_core_KE_n2457) );
  AOI22X1 U26389 ( .A0(n2312), .A1(top_core_KE_n2460), .B0(n2320), .B1(
        top_core_KE_CipherKey0_73_), .Y(top_core_KE_n2458) );
  NAND3X1 U26390 ( .A(top_core_KE_n2329), .B(top_core_KE_n2330), .C(
        top_core_KE_n2331), .Y(top_core_KE_n4822) );
  AOI222X1 U26391 ( .A0(top_core_KE_prev_key1_reg_97_), .A1(n2297), .B0(n2309), 
        .B1(top_core_KE_CipherKey0_33_), .C0(n2358), .C1(n6796), .Y(
        top_core_KE_n2331) );
  AOI22X1 U26392 ( .A0(n2314), .A1(top_core_KE_n2332), .B0(n2318), .B1(
        top_core_KE_CipherKey0_97_), .Y(top_core_KE_n2330) );
  AOI22X1 U26393 ( .A0(n2328), .A1(top_core_KE_n1121), .B0(n2338), .B1(
        top_core_KE_n1123), .Y(top_core_KE_n2329) );
  NAND3X1 U26394 ( .A(top_core_KE_n2497), .B(top_core_KE_n2498), .C(
        top_core_KE_n2499), .Y(top_core_KE_n4854) );
  AOI222X1 U26395 ( .A0(n1739), .A1(n2304), .B0(n2307), .B1(
        top_core_KE_CipherKey0_1_), .C0(n2355), .C1(top_core_KE_n1343), .Y(
        top_core_KE_n2499) );
  AOI22X1 U26396 ( .A0(n2330), .A1(top_core_KE_n1345), .B0(n2340), .B1(
        top_core_KE_n1347), .Y(top_core_KE_n2497) );
  AOI22X1 U26397 ( .A0(n2312), .A1(top_core_KE_n2500), .B0(n2321), .B1(
        top_core_KE_CipherKey0_65_), .Y(top_core_KE_n2498) );
  NAND3X1 U26398 ( .A(top_core_KE_n2284), .B(top_core_KE_n2285), .C(
        top_core_KE_n2286), .Y(top_core_KE_n4813) );
  AOI222X1 U26399 ( .A0(top_core_KE_prev_key1_reg_106_), .A1(n2294), .B0(
        top_core_KE_n2176), .B1(top_core_KE_CipherKey0_42_), .C0(n2359), .C1(
        n6730), .Y(top_core_KE_n2286) );
  AOI22X1 U26400 ( .A0(n2314), .A1(top_core_KE_n2287), .B0(n2317), .B1(
        top_core_KE_CipherKey0_106_), .Y(top_core_KE_n2285) );
  AOI22X1 U26401 ( .A0(n2327), .A1(top_core_KE_n1058), .B0(n2337), .B1(
        top_core_KE_n1060), .Y(top_core_KE_n2284) );
  NAND3X1 U26402 ( .A(top_core_KE_n2452), .B(top_core_KE_n2453), .C(
        top_core_KE_n2454), .Y(top_core_KE_n4845) );
  AOI222X1 U26403 ( .A0(n1703), .A1(top_core_KE_n2175), .B0(n2307), .B1(
        top_core_KE_CipherKey0_10_), .C0(n2352), .C1(top_core_KE_n1280), .Y(
        top_core_KE_n2454) );
  AOI22X1 U26404 ( .A0(n2329), .A1(top_core_KE_n1282), .B0(n2339), .B1(
        top_core_KE_n1284), .Y(top_core_KE_n2452) );
  AOI22X1 U26405 ( .A0(n2312), .A1(top_core_KE_n2455), .B0(n2320), .B1(
        top_core_KE_CipherKey0_74_), .Y(top_core_KE_n2453) );
  NAND3X1 U26406 ( .A(top_core_KE_n2324), .B(top_core_KE_n2325), .C(
        top_core_KE_n2326), .Y(top_core_KE_n4821) );
  AOI222X1 U26407 ( .A0(top_core_KE_prev_key1_reg_98_), .A1(n2297), .B0(n2309), 
        .B1(top_core_KE_CipherKey0_34_), .C0(n2358), .C1(n6793), .Y(
        top_core_KE_n2326) );
  AOI22X1 U26408 ( .A0(n2314), .A1(top_core_KE_n2327), .B0(n2318), .B1(
        top_core_KE_CipherKey0_98_), .Y(top_core_KE_n2325) );
  AOI22X1 U26409 ( .A0(n2328), .A1(top_core_KE_n1114), .B0(n2338), .B1(
        top_core_KE_n1116), .Y(top_core_KE_n2324) );
  NAND3X1 U26410 ( .A(top_core_KE_n2492), .B(top_core_KE_n2493), .C(
        top_core_KE_n2494), .Y(top_core_KE_n4853) );
  AOI222X1 U26411 ( .A0(n1732), .A1(n2304), .B0(n2307), .B1(
        top_core_KE_CipherKey0_2_), .C0(n2356), .C1(top_core_KE_n1336), .Y(
        top_core_KE_n2494) );
  AOI22X1 U26412 ( .A0(n2330), .A1(top_core_KE_n1338), .B0(n2340), .B1(
        top_core_KE_n1340), .Y(top_core_KE_n2492) );
  AOI22X1 U26413 ( .A0(n2312), .A1(top_core_KE_n2495), .B0(n2321), .B1(
        top_core_KE_CipherKey0_66_), .Y(top_core_KE_n2493) );
  NAND3X1 U26414 ( .A(top_core_KE_n2279), .B(top_core_KE_n2280), .C(
        top_core_KE_n2281), .Y(top_core_KE_n4812) );
  AOI222X1 U26415 ( .A0(top_core_KE_prev_key1_reg_107_), .A1(n2295), .B0(
        top_core_KE_n2176), .B1(top_core_KE_CipherKey0_43_), .C0(n2359), .C1(
        n6734), .Y(top_core_KE_n2281) );
  AOI22X1 U26416 ( .A0(n2315), .A1(top_core_KE_n2282), .B0(n2318), .B1(
        top_core_KE_CipherKey0_107_), .Y(top_core_KE_n2280) );
  AOI22X1 U26417 ( .A0(n2327), .A1(top_core_KE_n1051), .B0(n2337), .B1(
        top_core_KE_n1053), .Y(top_core_KE_n2279) );
  NAND3X1 U26418 ( .A(top_core_KE_n2447), .B(top_core_KE_n2448), .C(
        top_core_KE_n2449), .Y(top_core_KE_n4844) );
  AOI222X1 U26419 ( .A0(n1347), .A1(n2291), .B0(n2307), .B1(
        top_core_KE_CipherKey0_11_), .C0(n2352), .C1(top_core_KE_n1273), .Y(
        top_core_KE_n2449) );
  AOI22X1 U26420 ( .A0(n2329), .A1(top_core_KE_n1275), .B0(n2339), .B1(
        top_core_KE_n1277), .Y(top_core_KE_n2447) );
  AOI22X1 U26421 ( .A0(n2312), .A1(top_core_KE_n2450), .B0(n2320), .B1(
        top_core_KE_CipherKey0_75_), .Y(top_core_KE_n2448) );
  NAND3X1 U26422 ( .A(top_core_KE_n2319), .B(top_core_KE_n2320), .C(
        top_core_KE_n2321), .Y(top_core_KE_n4820) );
  AOI222X1 U26423 ( .A0(top_core_KE_prev_key1_reg_99_), .A1(n2297), .B0(n2309), 
        .B1(top_core_KE_CipherKey0_35_), .C0(n2358), .C1(n6791), .Y(
        top_core_KE_n2321) );
  AOI22X1 U26424 ( .A0(n2314), .A1(top_core_KE_n2322), .B0(n2318), .B1(
        top_core_KE_CipherKey0_99_), .Y(top_core_KE_n2320) );
  AOI22X1 U26425 ( .A0(n2328), .A1(top_core_KE_n1107), .B0(n2338), .B1(
        top_core_KE_n1109), .Y(top_core_KE_n2319) );
  NAND3X1 U26426 ( .A(top_core_KE_n2487), .B(top_core_KE_n2488), .C(
        top_core_KE_n2489), .Y(top_core_KE_n4852) );
  AOI222X1 U26427 ( .A0(n1349), .A1(n2304), .B0(n2307), .B1(
        top_core_KE_CipherKey0_3_), .C0(n2352), .C1(top_core_KE_n1329), .Y(
        top_core_KE_n2489) );
  AOI22X1 U26428 ( .A0(n2330), .A1(top_core_KE_n1331), .B0(n2340), .B1(
        top_core_KE_n1333), .Y(top_core_KE_n2487) );
  AOI22X1 U26429 ( .A0(n2312), .A1(top_core_KE_n2490), .B0(n2321), .B1(
        top_core_KE_CipherKey0_67_), .Y(top_core_KE_n2488) );
  NAND3X1 U26430 ( .A(top_core_KE_n2274), .B(top_core_KE_n2275), .C(
        top_core_KE_n2276), .Y(top_core_KE_n4811) );
  AOI222X1 U26431 ( .A0(top_core_KE_prev_key1_reg_108_), .A1(n2294), .B0(
        top_core_KE_n2176), .B1(top_core_KE_CipherKey0_44_), .C0(n2359), .C1(
        n6727), .Y(top_core_KE_n2276) );
  AOI22X1 U26432 ( .A0(n2312), .A1(top_core_KE_n2277), .B0(n2320), .B1(
        top_core_KE_CipherKey0_108_), .Y(top_core_KE_n2275) );
  AOI22X1 U26433 ( .A0(n2327), .A1(top_core_KE_n1044), .B0(n2337), .B1(
        top_core_KE_n1046), .Y(top_core_KE_n2274) );
  NAND3X1 U26434 ( .A(top_core_KE_n2442), .B(top_core_KE_n2443), .C(
        top_core_KE_n2444), .Y(top_core_KE_n4843) );
  AOI222X1 U26435 ( .A0(n1351), .A1(n2304), .B0(n2308), .B1(
        top_core_KE_CipherKey0_12_), .C0(n2353), .C1(top_core_KE_n1266), .Y(
        top_core_KE_n2444) );
  AOI22X1 U26436 ( .A0(n2329), .A1(top_core_KE_n1268), .B0(n2339), .B1(
        top_core_KE_n1270), .Y(top_core_KE_n2442) );
  AOI22X1 U26437 ( .A0(n2313), .A1(top_core_KE_n2445), .B0(n2320), .B1(
        top_core_KE_CipherKey0_76_), .Y(top_core_KE_n2443) );
  NAND3X1 U26438 ( .A(top_core_KE_n2314), .B(top_core_KE_n2315), .C(
        top_core_KE_n2316), .Y(top_core_KE_n4819) );
  AOI222X1 U26439 ( .A0(top_core_KE_prev_key1_reg_100_), .A1(n2296), .B0(n2310), .B1(top_core_KE_CipherKey0_36_), .C0(n767), .C1(n6789), .Y(top_core_KE_n2316) );
  AOI22X1 U26440 ( .A0(n2313), .A1(top_core_KE_n2317), .B0(n2318), .B1(
        top_core_KE_CipherKey0_100_), .Y(top_core_KE_n2315) );
  AOI22X1 U26441 ( .A0(n2328), .A1(top_core_KE_n1100), .B0(n2338), .B1(
        top_core_KE_n1102), .Y(top_core_KE_n2314) );
  NAND3X1 U26442 ( .A(top_core_KE_n2482), .B(top_core_KE_n2483), .C(
        top_core_KE_n2484), .Y(top_core_KE_n4851) );
  AOI222X1 U26443 ( .A0(n1353), .A1(n2304), .B0(n2307), .B1(
        top_core_KE_CipherKey0_4_), .C0(n767), .C1(top_core_KE_n1322), .Y(
        top_core_KE_n2484) );
  AOI22X1 U26444 ( .A0(n2329), .A1(top_core_KE_n1324), .B0(n2339), .B1(
        top_core_KE_n1326), .Y(top_core_KE_n2482) );
  AOI22X1 U26445 ( .A0(n2312), .A1(top_core_KE_n2485), .B0(n2320), .B1(
        top_core_KE_CipherKey0_68_), .Y(top_core_KE_n2483) );
  NAND3X1 U26446 ( .A(top_core_KE_n2269), .B(top_core_KE_n2270), .C(
        top_core_KE_n2271), .Y(top_core_KE_n4810) );
  AOI222X1 U26447 ( .A0(top_core_KE_prev_key1_reg_109_), .A1(n2296), .B0(n2307), .B1(top_core_KE_CipherKey0_45_), .C0(n2360), .C1(n6724), .Y(
        top_core_KE_n2271) );
  AOI22X1 U26448 ( .A0(n2314), .A1(top_core_KE_n2272), .B0(n2319), .B1(
        top_core_KE_CipherKey0_109_), .Y(top_core_KE_n2270) );
  AOI22X1 U26449 ( .A0(n2327), .A1(top_core_KE_n1037), .B0(n2337), .B1(
        top_core_KE_n1039), .Y(top_core_KE_n2269) );
  NAND3X1 U26450 ( .A(top_core_KE_n2437), .B(top_core_KE_n2438), .C(
        top_core_KE_n2439), .Y(top_core_KE_n4842) );
  AOI222X1 U26451 ( .A0(n1696), .A1(n2303), .B0(n2308), .B1(
        top_core_KE_CipherKey0_13_), .C0(n2353), .C1(top_core_KE_n1259), .Y(
        top_core_KE_n2439) );
  AOI22X1 U26452 ( .A0(n2329), .A1(top_core_KE_n1261), .B0(n2339), .B1(
        top_core_KE_n1263), .Y(top_core_KE_n2437) );
  AOI22X1 U26453 ( .A0(n2313), .A1(top_core_KE_n2440), .B0(n2320), .B1(
        top_core_KE_CipherKey0_77_), .Y(top_core_KE_n2438) );
  NAND3X1 U26454 ( .A(top_core_KE_n2309), .B(top_core_KE_n2310), .C(
        top_core_KE_n2311), .Y(top_core_KE_n4818) );
  AOI222X1 U26455 ( .A0(top_core_KE_prev_key1_reg_101_), .A1(n2296), .B0(n2308), .B1(top_core_KE_CipherKey0_37_), .C0(n2356), .C1(n6782), .Y(
        top_core_KE_n2311) );
  AOI22X1 U26456 ( .A0(n2315), .A1(top_core_KE_n2312), .B0(n2318), .B1(
        top_core_KE_CipherKey0_101_), .Y(top_core_KE_n2310) );
  AOI22X1 U26457 ( .A0(n2328), .A1(top_core_KE_n1093), .B0(n2338), .B1(
        top_core_KE_n1095), .Y(top_core_KE_n2309) );
  NAND3X1 U26458 ( .A(top_core_KE_n2477), .B(top_core_KE_n2478), .C(
        top_core_KE_n2479), .Y(top_core_KE_n4850) );
  AOI222X1 U26459 ( .A0(n1725), .A1(n2303), .B0(n2307), .B1(
        top_core_KE_CipherKey0_5_), .C0(n767), .C1(top_core_KE_n1315), .Y(
        top_core_KE_n2479) );
  AOI22X1 U26460 ( .A0(n2329), .A1(top_core_KE_n1317), .B0(n2339), .B1(
        top_core_KE_n1319), .Y(top_core_KE_n2477) );
  AOI22X1 U26461 ( .A0(n2312), .A1(top_core_KE_n2480), .B0(n2320), .B1(
        top_core_KE_CipherKey0_69_), .Y(top_core_KE_n2478) );
  NAND3X1 U26462 ( .A(top_core_KE_n2264), .B(top_core_KE_n2265), .C(
        top_core_KE_n2266), .Y(top_core_KE_n4809) );
  AOI222X1 U26463 ( .A0(top_core_KE_prev_key1_reg_110_), .A1(n2295), .B0(n2309), .B1(top_core_KE_CipherKey0_46_), .C0(n2360), .C1(n6718), .Y(
        top_core_KE_n2266) );
  AOI22X1 U26464 ( .A0(n2312), .A1(top_core_KE_n2267), .B0(n2317), .B1(
        top_core_KE_CipherKey0_110_), .Y(top_core_KE_n2265) );
  AOI22X1 U26465 ( .A0(n2327), .A1(top_core_KE_n1030), .B0(n2337), .B1(
        top_core_KE_n1032), .Y(top_core_KE_n2264) );
  NAND3X1 U26466 ( .A(top_core_KE_n2432), .B(top_core_KE_n2433), .C(
        top_core_KE_n2434), .Y(top_core_KE_n4841) );
  AOI222X1 U26467 ( .A0(n1355), .A1(n2303), .B0(n2308), .B1(
        top_core_KE_CipherKey0_14_), .C0(n2353), .C1(top_core_KE_n1252), .Y(
        top_core_KE_n2434) );
  AOI22X1 U26468 ( .A0(n2329), .A1(top_core_KE_n1254), .B0(n2339), .B1(
        top_core_KE_n1256), .Y(top_core_KE_n2432) );
  AOI22X1 U26469 ( .A0(n2313), .A1(top_core_KE_n2435), .B0(n2320), .B1(
        top_core_KE_CipherKey0_78_), .Y(top_core_KE_n2433) );
  NAND3X1 U26470 ( .A(top_core_KE_n2392), .B(top_core_KE_n2393), .C(
        top_core_KE_n2394), .Y(top_core_KE_n4833) );
  AOI222X1 U26471 ( .A0(n1356), .A1(n2300), .B0(n2308), .B1(
        top_core_KE_CipherKey0_22_), .C0(n2358), .C1(top_core_KE_n1196), .Y(
        top_core_KE_n2394) );
  AOI22X1 U26472 ( .A0(top_core_KE_n2181), .A1(top_core_KE_n1198), .B0(n2339), 
        .B1(top_core_KE_n1200), .Y(top_core_KE_n2392) );
  AOI22X1 U26473 ( .A0(n2313), .A1(top_core_KE_n2395), .B0(n2319), .B1(
        top_core_KE_CipherKey0_86_), .Y(top_core_KE_n2393) );
  NAND3X1 U26474 ( .A(top_core_KE_n2214), .B(top_core_KE_n2215), .C(
        top_core_KE_n2216), .Y(top_core_KE_n4799) );
  AOI222X1 U26475 ( .A0(top_core_KE_prev_key1_reg_120_), .A1(n2291), .B0(n2310), .B1(top_core_KE_CipherKey0_56_), .C0(n2362), .C1(n6357), .Y(
        top_core_KE_n2216) );
  AOI22X1 U26476 ( .A0(n2328), .A1(top_core_KE_n960), .B0(top_core_KE_n2182), 
        .B1(top_core_KE_n962), .Y(top_core_KE_n2214) );
  AOI22X1 U26477 ( .A0(n2315), .A1(top_core_KE_n2217), .B0(n2317), .B1(
        top_core_KE_CipherKey0_120_), .Y(top_core_KE_n2215) );
  NAND3X1 U26478 ( .A(top_core_KE_n2381), .B(top_core_KE_n2382), .C(
        top_core_KE_n2383), .Y(top_core_KE_n4831) );
  AOI222X1 U26479 ( .A0(n1659), .A1(n2300), .B0(n2309), .B1(
        top_core_KE_CipherKey0_24_), .C0(n2355), .C1(n6356), .Y(
        top_core_KE_n2383) );
  AOI22X1 U26480 ( .A0(top_core_KE_n2181), .A1(top_core_KE_n1184), .B0(n2338), 
        .B1(top_core_KE_n1186), .Y(top_core_KE_n2381) );
  AOI22X1 U26481 ( .A0(n2314), .A1(top_core_KE_n2384), .B0(n2319), .B1(
        top_core_KE_CipherKey0_88_), .Y(top_core_KE_n2382) );
  NAND3X1 U26482 ( .A(top_core_KE_n2254), .B(top_core_KE_n2255), .C(
        top_core_KE_n2256), .Y(top_core_KE_n4807) );
  AOI222X1 U26483 ( .A0(top_core_KE_prev_key1_reg_112_), .A1(n2295), .B0(n2310), .B1(top_core_KE_CipherKey0_48_), .C0(n767), .C1(top_core_KE_n1014), .Y(
        top_core_KE_n2256) );
  AOI22X1 U26484 ( .A0(n2315), .A1(top_core_KE_n2257), .B0(n2318), .B1(
        top_core_KE_CipherKey0_112_), .Y(top_core_KE_n2255) );
  AOI22X1 U26485 ( .A0(n2327), .A1(top_core_KE_n1016), .B0(n2337), .B1(
        top_core_KE_n1018), .Y(top_core_KE_n2254) );
  NAND3X1 U26486 ( .A(top_core_KE_n2422), .B(top_core_KE_n2423), .C(
        top_core_KE_n2424), .Y(top_core_KE_n4839) );
  AOI222X1 U26487 ( .A0(n1688), .A1(n2302), .B0(n2308), .B1(
        top_core_KE_CipherKey0_16_), .C0(n2354), .C1(top_core_KE_n1238), .Y(
        top_core_KE_n2424) );
  AOI22X1 U26488 ( .A0(top_core_KE_n2181), .A1(top_core_KE_n1240), .B0(n2337), 
        .B1(top_core_KE_n1242), .Y(top_core_KE_n2422) );
  AOI22X1 U26489 ( .A0(n2313), .A1(top_core_KE_n2425), .B0(n2319), .B1(
        top_core_KE_CipherKey0_80_), .Y(top_core_KE_n2423) );
  NAND3X1 U26490 ( .A(top_core_KE_n2249), .B(top_core_KE_n2250), .C(
        top_core_KE_n2251), .Y(top_core_KE_n4806) );
  AOI222X1 U26491 ( .A0(top_core_KE_prev_key1_reg_113_), .A1(n2295), .B0(n2310), .B1(top_core_KE_CipherKey0_49_), .C0(n2359), .C1(top_core_KE_n1007), .Y(
        top_core_KE_n2251) );
  AOI22X1 U26492 ( .A0(n2315), .A1(top_core_KE_n2252), .B0(n2320), .B1(
        top_core_KE_CipherKey0_113_), .Y(top_core_KE_n2250) );
  AOI22X1 U26493 ( .A0(n2327), .A1(top_core_KE_n1009), .B0(n2337), .B1(
        top_core_KE_n1011), .Y(top_core_KE_n2249) );
  NAND3X1 U26494 ( .A(top_core_KE_n2417), .B(top_core_KE_n2418), .C(
        top_core_KE_n2419), .Y(top_core_KE_n4838) );
  AOI222X1 U26495 ( .A0(n1681), .A1(n2302), .B0(n2308), .B1(
        top_core_KE_CipherKey0_17_), .C0(n2354), .C1(top_core_KE_n1231), .Y(
        top_core_KE_n2419) );
  AOI22X1 U26496 ( .A0(top_core_KE_n2181), .A1(top_core_KE_n1233), .B0(n2339), 
        .B1(top_core_KE_n1235), .Y(top_core_KE_n2417) );
  AOI22X1 U26497 ( .A0(n2313), .A1(top_core_KE_n2420), .B0(n2319), .B1(
        top_core_KE_CipherKey0_81_), .Y(top_core_KE_n2418) );
  NAND3X1 U26498 ( .A(top_core_KE_n2204), .B(top_core_KE_n2205), .C(
        top_core_KE_n2206), .Y(top_core_KE_n4797) );
  AOI222X1 U26499 ( .A0(top_core_KE_prev_key1_reg_122_), .A1(n2293), .B0(n2310), .B1(top_core_KE_CipherKey0_58_), .C0(n2361), .C1(n6371), .Y(
        top_core_KE_n2206) );
  AOI22X1 U26500 ( .A0(n2327), .A1(top_core_KE_n946), .B0(top_core_KE_n2182), 
        .B1(top_core_KE_n948), .Y(top_core_KE_n2204) );
  AOI22X1 U26501 ( .A0(n2315), .A1(top_core_KE_n2207), .B0(n2317), .B1(
        top_core_KE_CipherKey0_122_), .Y(top_core_KE_n2205) );
  NAND3X1 U26502 ( .A(top_core_KE_n2369), .B(top_core_KE_n2370), .C(
        top_core_KE_n2371), .Y(top_core_KE_n4829) );
  AOI222X1 U26503 ( .A0(n1649), .A1(n2299), .B0(n2309), .B1(
        top_core_KE_CipherKey0_26_), .C0(n2355), .C1(n6370), .Y(
        top_core_KE_n2371) );
  AOI22X1 U26504 ( .A0(top_core_KE_n2181), .A1(top_core_KE_n1170), .B0(n2338), 
        .B1(top_core_KE_n1172), .Y(top_core_KE_n2369) );
  AOI22X1 U26505 ( .A0(n2314), .A1(top_core_KE_n2372), .B0(n2319), .B1(
        top_core_KE_CipherKey0_90_), .Y(top_core_KE_n2370) );
  NAND3X1 U26506 ( .A(top_core_KE_n2244), .B(top_core_KE_n2245), .C(
        top_core_KE_n2246), .Y(top_core_KE_n4805) );
  AOI222X1 U26507 ( .A0(top_core_KE_prev_key1_reg_114_), .A1(n2295), .B0(n2310), .B1(top_core_KE_CipherKey0_50_), .C0(n2357), .C1(top_core_KE_n1000), .Y(
        top_core_KE_n2246) );
  AOI22X1 U26508 ( .A0(n2315), .A1(top_core_KE_n2247), .B0(n2319), .B1(
        top_core_KE_CipherKey0_114_), .Y(top_core_KE_n2245) );
  AOI22X1 U26509 ( .A0(n2327), .A1(top_core_KE_n1002), .B0(n2337), .B1(
        top_core_KE_n1004), .Y(top_core_KE_n2244) );
  NAND3X1 U26510 ( .A(top_core_KE_n2412), .B(top_core_KE_n2413), .C(
        top_core_KE_n2414), .Y(top_core_KE_n4837) );
  AOI222X1 U26511 ( .A0(n1674), .A1(n2302), .B0(n2308), .B1(
        top_core_KE_CipherKey0_18_), .C0(n2361), .C1(top_core_KE_n1224), .Y(
        top_core_KE_n2414) );
  AOI22X1 U26512 ( .A0(top_core_KE_n2181), .A1(top_core_KE_n1226), .B0(n2337), 
        .B1(top_core_KE_n1228), .Y(top_core_KE_n2412) );
  AOI22X1 U26513 ( .A0(n2313), .A1(top_core_KE_n2415), .B0(n2319), .B1(
        top_core_KE_CipherKey0_82_), .Y(top_core_KE_n2413) );
  NAND3X1 U26514 ( .A(top_core_KE_n2199), .B(top_core_KE_n2200), .C(
        top_core_KE_n2201), .Y(top_core_KE_n4796) );
  AOI222X1 U26515 ( .A0(top_core_KE_prev_key1_reg_123_), .A1(n2293), .B0(n2310), .B1(top_core_KE_CipherKey0_59_), .C0(n2361), .C1(n6367), .Y(
        top_core_KE_n2201) );
  AOI22X1 U26516 ( .A0(n2329), .A1(top_core_KE_n939), .B0(top_core_KE_n2182), 
        .B1(top_core_KE_n941), .Y(top_core_KE_n2199) );
  AOI22X1 U26517 ( .A0(n2315), .A1(top_core_KE_n2202), .B0(n2317), .B1(
        top_core_KE_CipherKey0_123_), .Y(top_core_KE_n2200) );
  NAND3X1 U26518 ( .A(top_core_KE_n2363), .B(top_core_KE_n2364), .C(
        top_core_KE_n2365), .Y(top_core_KE_n4828) );
  AOI222X1 U26519 ( .A0(n1361), .A1(n2299), .B0(n2309), .B1(
        top_core_KE_CipherKey0_27_), .C0(n2356), .C1(n6366), .Y(
        top_core_KE_n2365) );
  AOI22X1 U26520 ( .A0(top_core_KE_n2181), .A1(top_core_KE_n1163), .B0(n2339), 
        .B1(top_core_KE_n1165), .Y(top_core_KE_n2363) );
  AOI22X1 U26521 ( .A0(n2314), .A1(top_core_KE_n2366), .B0(n2319), .B1(
        top_core_KE_CipherKey0_91_), .Y(top_core_KE_n2364) );
  NAND3X1 U26522 ( .A(top_core_KE_n2239), .B(top_core_KE_n2240), .C(
        top_core_KE_n2241), .Y(top_core_KE_n4804) );
  AOI222X1 U26523 ( .A0(top_core_KE_prev_key1_reg_115_), .A1(n2294), .B0(n2310), .B1(top_core_KE_CipherKey0_51_), .C0(n2353), .C1(top_core_KE_n993), .Y(
        top_core_KE_n2241) );
  AOI22X1 U26524 ( .A0(n2315), .A1(top_core_KE_n2242), .B0(n2317), .B1(
        top_core_KE_CipherKey0_115_), .Y(top_core_KE_n2240) );
  AOI22X1 U26525 ( .A0(n2327), .A1(top_core_KE_n995), .B0(n2337), .B1(
        top_core_KE_n997), .Y(top_core_KE_n2239) );
  NAND3X1 U26526 ( .A(top_core_KE_n2407), .B(top_core_KE_n2408), .C(
        top_core_KE_n2409), .Y(top_core_KE_n4836) );
  AOI222X1 U26527 ( .A0(n1363), .A1(n2301), .B0(n2308), .B1(
        top_core_KE_CipherKey0_19_), .C0(n2351), .C1(top_core_KE_n1217), .Y(
        top_core_KE_n2409) );
  AOI22X1 U26528 ( .A0(n2328), .A1(top_core_KE_n1219), .B0(n2340), .B1(
        top_core_KE_n1221), .Y(top_core_KE_n2407) );
  AOI22X1 U26529 ( .A0(n2313), .A1(top_core_KE_n2410), .B0(n2319), .B1(
        top_core_KE_CipherKey0_83_), .Y(top_core_KE_n2408) );
  NAND3X1 U26530 ( .A(top_core_KE_n2194), .B(top_core_KE_n2195), .C(
        top_core_KE_n2196), .Y(top_core_KE_n4795) );
  AOI222X1 U26531 ( .A0(top_core_KE_prev_key1_reg_124_), .A1(n2284), .B0(
        top_core_KE_n2176), .B1(top_core_KE_CipherKey0_60_), .C0(n2362), .C1(
        n6353), .Y(top_core_KE_n2196) );
  AOI22X1 U26532 ( .A0(n2328), .A1(top_core_KE_n932), .B0(top_core_KE_n2182), 
        .B1(top_core_KE_n934), .Y(top_core_KE_n2194) );
  AOI22X1 U26533 ( .A0(n2312), .A1(top_core_KE_n2197), .B0(n2317), .B1(
        top_core_KE_CipherKey0_124_), .Y(top_core_KE_n2195) );
  NAND3X1 U26534 ( .A(top_core_KE_n2357), .B(top_core_KE_n2358), .C(
        top_core_KE_n2359), .Y(top_core_KE_n4827) );
  AOI222X1 U26535 ( .A0(n1365), .A1(n2298), .B0(n2309), .B1(
        top_core_KE_CipherKey0_28_), .C0(n2356), .C1(n6352), .Y(
        top_core_KE_n2359) );
  AOI22X1 U26536 ( .A0(n2328), .A1(top_core_KE_n1156), .B0(n2338), .B1(
        top_core_KE_n1158), .Y(top_core_KE_n2357) );
  AOI22X1 U26537 ( .A0(n2314), .A1(top_core_KE_n2360), .B0(n2318), .B1(
        top_core_KE_CipherKey0_92_), .Y(top_core_KE_n2358) );
  NAND3X1 U26538 ( .A(top_core_KE_n2234), .B(top_core_KE_n2235), .C(
        top_core_KE_n2236), .Y(top_core_KE_n4803) );
  AOI222X1 U26539 ( .A0(top_core_KE_prev_key1_reg_116_), .A1(n2294), .B0(n2310), .B1(top_core_KE_CipherKey0_52_), .C0(n2354), .C1(top_core_KE_n986), .Y(
        top_core_KE_n2236) );
  AOI22X1 U26540 ( .A0(n2315), .A1(top_core_KE_n2237), .B0(n2317), .B1(
        top_core_KE_CipherKey0_116_), .Y(top_core_KE_n2235) );
  AOI22X1 U26541 ( .A0(n2327), .A1(top_core_KE_n988), .B0(top_core_KE_n2182), 
        .B1(top_core_KE_n990), .Y(top_core_KE_n2234) );
  NAND3X1 U26542 ( .A(top_core_KE_n2402), .B(top_core_KE_n2403), .C(
        top_core_KE_n2404), .Y(top_core_KE_n4835) );
  AOI222X1 U26543 ( .A0(n1367), .A1(n2301), .B0(n2308), .B1(
        top_core_KE_CipherKey0_20_), .C0(n2358), .C1(top_core_KE_n1210), .Y(
        top_core_KE_n2404) );
  AOI22X1 U26544 ( .A0(n2327), .A1(top_core_KE_n1212), .B0(n2338), .B1(
        top_core_KE_n1214), .Y(top_core_KE_n2402) );
  AOI22X1 U26545 ( .A0(n2313), .A1(top_core_KE_n2405), .B0(n2319), .B1(
        top_core_KE_CipherKey0_84_), .Y(top_core_KE_n2403) );
  NAND3X1 U26546 ( .A(top_core_KE_n2189), .B(top_core_KE_n2190), .C(
        top_core_KE_n2191), .Y(top_core_KE_n4794) );
  AOI222X1 U26547 ( .A0(top_core_KE_prev_key1_reg_125_), .A1(n2291), .B0(
        top_core_KE_n2176), .B1(top_core_KE_CipherKey0_61_), .C0(n2362), .C1(
        n6363), .Y(top_core_KE_n2191) );
  AOI22X1 U26548 ( .A0(n2329), .A1(top_core_KE_n925), .B0(top_core_KE_n2182), 
        .B1(top_core_KE_n927), .Y(top_core_KE_n2189) );
  AOI22X1 U26549 ( .A0(n2313), .A1(top_core_KE_n2192), .B0(n2317), .B1(
        top_core_KE_CipherKey0_125_), .Y(top_core_KE_n2190) );
  NAND3X1 U26550 ( .A(top_core_KE_n2351), .B(top_core_KE_n2352), .C(
        top_core_KE_n2353), .Y(top_core_KE_n4826) );
  AOI222X1 U26551 ( .A0(n1640), .A1(n2298), .B0(n2309), .B1(
        top_core_KE_CipherKey0_29_), .C0(n2356), .C1(n6362), .Y(
        top_core_KE_n2353) );
  AOI22X1 U26552 ( .A0(n2328), .A1(top_core_KE_n1149), .B0(n2338), .B1(
        top_core_KE_n1151), .Y(top_core_KE_n2351) );
  AOI22X1 U26553 ( .A0(n2314), .A1(top_core_KE_n2354), .B0(n2318), .B1(
        top_core_KE_CipherKey0_93_), .Y(top_core_KE_n2352) );
  NAND3X1 U26554 ( .A(top_core_KE_n2229), .B(top_core_KE_n2230), .C(
        top_core_KE_n2231), .Y(top_core_KE_n4802) );
  AOI222X1 U26555 ( .A0(top_core_KE_prev_key1_reg_117_), .A1(n2294), .B0(n2310), .B1(top_core_KE_CipherKey0_53_), .C0(n2361), .C1(top_core_KE_n979), .Y(
        top_core_KE_n2231) );
  AOI22X1 U26556 ( .A0(n2315), .A1(top_core_KE_n2232), .B0(n2317), .B1(
        top_core_KE_CipherKey0_117_), .Y(top_core_KE_n2230) );
  AOI22X1 U26557 ( .A0(n2328), .A1(top_core_KE_n981), .B0(top_core_KE_n2182), 
        .B1(top_core_KE_n983), .Y(top_core_KE_n2229) );
  NAND3X1 U26558 ( .A(top_core_KE_n2397), .B(top_core_KE_n2398), .C(
        top_core_KE_n2399), .Y(top_core_KE_n4834) );
  AOI222X1 U26559 ( .A0(n1667), .A1(n2301), .B0(n2308), .B1(
        top_core_KE_CipherKey0_21_), .C0(n2360), .C1(top_core_KE_n1203), .Y(
        top_core_KE_n2399) );
  AOI22X1 U26560 ( .A0(n2329), .A1(top_core_KE_n1205), .B0(n2337), .B1(
        top_core_KE_n1207), .Y(top_core_KE_n2397) );
  AOI22X1 U26561 ( .A0(n2313), .A1(top_core_KE_n2400), .B0(n2319), .B1(
        top_core_KE_CipherKey0_85_), .Y(top_core_KE_n2398) );
  NAND3X1 U26562 ( .A(top_core_KE_n2184), .B(top_core_KE_n2185), .C(
        top_core_KE_n2186), .Y(top_core_KE_n4793) );
  AOI222X1 U26563 ( .A0(top_core_KE_prev_key1_reg_126_), .A1(n2293), .B0(
        top_core_KE_n2176), .B1(top_core_KE_CipherKey0_62_), .C0(n2362), .C1(
        n6349), .Y(top_core_KE_n2186) );
  AOI22X1 U26564 ( .A0(n2327), .A1(top_core_KE_n917), .B0(top_core_KE_n2182), 
        .B1(top_core_KE_n920), .Y(top_core_KE_n2184) );
  AOI22X1 U26565 ( .A0(n2314), .A1(top_core_KE_n2187), .B0(n2317), .B1(
        top_core_KE_CipherKey0_126_), .Y(top_core_KE_n2185) );
  NAND3X1 U26566 ( .A(top_core_KE_n2345), .B(top_core_KE_n2346), .C(
        top_core_KE_n2347), .Y(top_core_KE_n4825) );
  AOI222X1 U26567 ( .A0(n1369), .A1(n2298), .B0(n2309), .B1(
        top_core_KE_CipherKey0_30_), .C0(n2357), .C1(n6348), .Y(
        top_core_KE_n2347) );
  AOI22X1 U26568 ( .A0(n2328), .A1(top_core_KE_n1142), .B0(n2338), .B1(
        top_core_KE_n1144), .Y(top_core_KE_n2345) );
  AOI22X1 U26569 ( .A0(n2314), .A1(top_core_KE_n2348), .B0(n2318), .B1(
        top_core_KE_CipherKey0_94_), .Y(top_core_KE_n2346) );
  NAND3X1 U26570 ( .A(top_core_KE_n2224), .B(top_core_KE_n2225), .C(
        top_core_KE_n2226), .Y(top_core_KE_n4801) );
  AOI222X1 U26571 ( .A0(top_core_KE_prev_key1_reg_118_), .A1(n2292), .B0(n2310), .B1(top_core_KE_CipherKey0_54_), .C0(n2351), .C1(top_core_KE_n972), .Y(
        top_core_KE_n2226) );
  AOI22X1 U26572 ( .A0(n2315), .A1(top_core_KE_n2227), .B0(n2317), .B1(
        top_core_KE_CipherKey0_118_), .Y(top_core_KE_n2225) );
  AOI22X1 U26573 ( .A0(n2329), .A1(top_core_KE_n974), .B0(top_core_KE_n2182), 
        .B1(top_core_KE_n976), .Y(top_core_KE_n2224) );
  NAND3X1 U26574 ( .A(top_core_KE_n2219), .B(top_core_KE_n2220), .C(
        top_core_KE_n2221), .Y(top_core_KE_n4800) );
  AOI222X1 U26575 ( .A0(top_core_KE_prev_key1_reg_119_), .A1(top_core_KE_n2175), .B0(n2310), .B1(top_core_KE_CipherKey0_55_), .C0(n2352), .C1(
        top_core_KE_n965), .Y(top_core_KE_n2221) );
  AOI22X1 U26576 ( .A0(n2315), .A1(top_core_KE_n2222), .B0(n2317), .B1(
        top_core_KE_CipherKey0_119_), .Y(top_core_KE_n2220) );
  AOI22X1 U26577 ( .A0(n2330), .A1(top_core_KE_n967), .B0(n2338), .B1(
        top_core_KE_n969), .Y(top_core_KE_n2219) );
  NAND3X1 U26578 ( .A(top_core_KE_n2304), .B(top_core_KE_n2305), .C(
        top_core_KE_n2306), .Y(top_core_KE_n4817) );
  AOI222X1 U26579 ( .A0(top_core_KE_prev_key1_reg_102_), .A1(n2296), .B0(n2310), .B1(top_core_KE_CipherKey0_38_), .C0(n2357), .C1(n6385), .Y(
        top_core_KE_n2306) );
  AOI22X1 U26580 ( .A0(n2313), .A1(top_core_KE_n2307), .B0(n2318), .B1(
        top_core_KE_CipherKey0_102_), .Y(top_core_KE_n2305) );
  AOI22X1 U26581 ( .A0(n2328), .A1(top_core_KE_n1086), .B0(n2338), .B1(
        top_core_KE_n1088), .Y(top_core_KE_n2304) );
  NAND3X1 U26582 ( .A(top_core_KE_n2299), .B(top_core_KE_n2300), .C(
        top_core_KE_n2301), .Y(top_core_KE_n4816) );
  AOI222X1 U26583 ( .A0(top_core_KE_prev_key1_reg_103_), .A1(n2298), .B0(n2307), .B1(top_core_KE_CipherKey0_39_), .C0(n2359), .C1(n6378), .Y(
        top_core_KE_n2301) );
  AOI22X1 U26584 ( .A0(n2314), .A1(top_core_KE_n2302), .B0(n2318), .B1(
        top_core_KE_CipherKey0_103_), .Y(top_core_KE_n2300) );
  AOI22X1 U26585 ( .A0(n2328), .A1(top_core_KE_n1079), .B0(n2338), .B1(
        top_core_KE_n1081), .Y(top_core_KE_n2299) );
  NAND3X1 U26586 ( .A(top_core_KE_n2172), .B(top_core_KE_n2173), .C(
        top_core_KE_n2174), .Y(top_core_KE_n4792) );
  AOI222X1 U26587 ( .A0(top_core_KE_prev_key1_reg_127_), .A1(n2298), .B0(
        top_core_KE_n2176), .B1(top_core_KE_CipherKey0_63_), .C0(n767), .C1(
        top_core_KE_n902), .Y(top_core_KE_n2174) );
  AOI22X1 U26588 ( .A0(n2328), .A1(top_core_KE_n903), .B0(n2337), .B1(
        top_core_KE_n909), .Y(top_core_KE_n2172) );
  AOI22X1 U26589 ( .A0(n2315), .A1(top_core_KE_n2178), .B0(n2317), .B1(
        top_core_KE_CipherKey0_127_), .Y(top_core_KE_n2173) );
  NAND3X1 U26590 ( .A(top_core_KE_n2259), .B(top_core_KE_n2260), .C(
        top_core_KE_n2261), .Y(top_core_KE_n4808) );
  AOI222X1 U26591 ( .A0(top_core_KE_prev_key1_reg_111_), .A1(n2300), .B0(n2308), .B1(top_core_KE_CipherKey0_47_), .C0(n2360), .C1(n6329), .Y(
        top_core_KE_n2261) );
  AOI22X1 U26592 ( .A0(n2315), .A1(top_core_KE_n2262), .B0(n2318), .B1(
        top_core_KE_CipherKey0_111_), .Y(top_core_KE_n2260) );
  AOI22X1 U26593 ( .A0(n2327), .A1(top_core_KE_n1023), .B0(n2337), .B1(
        top_core_KE_n1025), .Y(top_core_KE_n2259) );
  NAND3X1 U26594 ( .A(top_core_KE_n2209), .B(top_core_KE_n2210), .C(
        top_core_KE_n2211), .Y(top_core_KE_n4798) );
  AOI222X1 U26595 ( .A0(top_core_KE_prev_key1_reg_121_), .A1(n2293), .B0(n2310), .B1(top_core_KE_CipherKey0_57_), .C0(n2361), .C1(n6315), .Y(
        top_core_KE_n2211) );
  AOI22X1 U26596 ( .A0(n2327), .A1(top_core_KE_n953), .B0(n2339), .B1(
        top_core_KE_n955), .Y(top_core_KE_n2209) );
  AOI22X1 U26597 ( .A0(n2315), .A1(top_core_KE_n2212), .B0(n2317), .B1(
        top_core_KE_CipherKey0_121_), .Y(top_core_KE_n2210) );
  BUFX3 U26598 ( .A(top_core_KE_prev_key1_reg_27_), .Y(n1360) );
  BUFX3 U26599 ( .A(top_core_KE_round_ctr_reg_2_), .Y(n1333) );
  INVX1 U26600 ( .A(top_core_KE_prev_key1_reg_63_), .Y(n6338) );
  BUFX3 U26601 ( .A(top_core_KE_prev_key1_reg_11_), .Y(n1346) );
  BUFX3 U26602 ( .A(top_core_KE_prev_key1_reg_3_), .Y(n1348) );
  BUFX3 U26603 ( .A(top_core_KE_prev_key1_reg_19_), .Y(n1362) );
  XNOR2X1 U26604 ( .A(n7246), .B(n3989), .Y(top_core_EC_n1034) );
  INVX1 U26605 ( .A(top_core_op), .Y(n4256) );
  BUFX3 U26606 ( .A(top_core_KE_round_ctr_reg_1_), .Y(n1332) );
  INVX1 U26607 ( .A(top_core_Nr[1]), .Y(n4195) );
  INVX1 U26608 ( .A(top_core_Nr[2]), .Y(n4196) );
  INVX1 U26609 ( .A(top_core_Nr[3]), .Y(n4197) );
  AOI221X1 U26610 ( .A0(top_core_KE_n965), .A1(n2196), .B0(n2213), .B1(
        top_core_KE_CipherKey0_119_), .C0(top_core_KE_n966), .Y(
        top_core_KE_n964) );
  OAI2BB2X1 U26611 ( .B0(n6394), .B1(n2228), .A0N(n1633), .A1N(
        top_core_KE_n967), .Y(top_core_KE_n966) );
  AOI221X1 U26612 ( .A0(top_core_KE_n972), .A1(n2196), .B0(n2215), .B1(
        top_core_KE_CipherKey0_118_), .C0(top_core_KE_n973), .Y(
        top_core_KE_n971) );
  OAI2BB2X1 U26613 ( .B0(n6402), .B1(n2228), .A0N(n1633), .A1N(
        top_core_KE_n974), .Y(top_core_KE_n973) );
  AOI221X1 U26614 ( .A0(top_core_KE_n979), .A1(n2197), .B0(n2212), .B1(
        top_core_KE_CipherKey0_117_), .C0(top_core_KE_n980), .Y(
        top_core_KE_n978) );
  OAI2BB2X1 U26615 ( .B0(n6480), .B1(n2229), .A0N(n1633), .A1N(
        top_core_KE_n981), .Y(top_core_KE_n980) );
  AOI221X1 U26616 ( .A0(top_core_KE_n986), .A1(n2197), .B0(n2212), .B1(
        top_core_KE_CipherKey0_116_), .C0(top_core_KE_n987), .Y(
        top_core_KE_n985) );
  OAI2BB2X1 U26617 ( .B0(n6560), .B1(n2229), .A0N(n1633), .A1N(
        top_core_KE_n988), .Y(top_core_KE_n987) );
  AOI221X1 U26618 ( .A0(top_core_KE_n993), .A1(n2197), .B0(n2212), .B1(
        top_core_KE_CipherKey0_115_), .C0(top_core_KE_n994), .Y(
        top_core_KE_n992) );
  OAI2BB2X1 U26619 ( .B0(n6639), .B1(n2235), .A0N(n1633), .A1N(
        top_core_KE_n995), .Y(top_core_KE_n994) );
  AOI221X1 U26620 ( .A0(top_core_KE_n1000), .A1(n2198), .B0(n2213), .B1(
        top_core_KE_CipherKey0_114_), .C0(top_core_KE_n1001), .Y(
        top_core_KE_n999) );
  OAI2BB2X1 U26621 ( .B0(n6667), .B1(n2228), .A0N(n1633), .A1N(
        top_core_KE_n1002), .Y(top_core_KE_n1001) );
  AOI221X1 U26622 ( .A0(top_core_KE_n1007), .A1(n2198), .B0(n2213), .B1(
        top_core_KE_CipherKey0_113_), .C0(top_core_KE_n1008), .Y(
        top_core_KE_n1006) );
  OAI2BB2X1 U26623 ( .B0(n6682), .B1(n2230), .A0N(n1633), .A1N(
        top_core_KE_n1009), .Y(top_core_KE_n1008) );
  AOI221X1 U26624 ( .A0(top_core_KE_n1014), .A1(n2198), .B0(n2213), .B1(
        top_core_KE_CipherKey0_112_), .C0(top_core_KE_n1015), .Y(
        top_core_KE_n1013) );
  OAI2BB2X1 U26625 ( .B0(n6689), .B1(n2230), .A0N(n1633), .A1N(
        top_core_KE_n1016), .Y(top_core_KE_n1015) );
  AOI221X1 U26626 ( .A0(top_core_KE_n1189), .A1(n2199), .B0(n2214), .B1(
        top_core_KE_CipherKey0_87_), .C0(top_core_KE_n1190), .Y(
        top_core_KE_n1188) );
  OAI2BB2X1 U26627 ( .B0(top_core_KE_n635), .B1(n2235), .A0N(n1632), .A1N(
        top_core_KE_n1191), .Y(top_core_KE_n1190) );
  AOI221X1 U26628 ( .A0(top_core_KE_n1196), .A1(n2199), .B0(n2215), .B1(
        top_core_KE_CipherKey0_86_), .C0(top_core_KE_n1197), .Y(
        top_core_KE_n1195) );
  OAI2BB2X1 U26629 ( .B0(top_core_KE_n636), .B1(n2228), .A0N(n1633), .A1N(
        top_core_KE_n1198), .Y(top_core_KE_n1197) );
  AOI221X1 U26630 ( .A0(top_core_KE_n1203), .A1(n2199), .B0(n2214), .B1(
        top_core_KE_CipherKey0_85_), .C0(top_core_KE_n1204), .Y(
        top_core_KE_n1202) );
  OAI2BB2X1 U26631 ( .B0(top_core_KE_n637), .B1(n2233), .A0N(n1632), .A1N(
        top_core_KE_n1205), .Y(top_core_KE_n1204) );
  AOI221X1 U26632 ( .A0(top_core_KE_n1210), .A1(n2199), .B0(n2214), .B1(
        top_core_KE_CipherKey0_84_), .C0(top_core_KE_n1211), .Y(
        top_core_KE_n1209) );
  OAI2BB2X1 U26633 ( .B0(top_core_KE_n638), .B1(n2234), .A0N(n1633), .A1N(
        top_core_KE_n1212), .Y(top_core_KE_n1211) );
  AOI221X1 U26634 ( .A0(top_core_KE_n1217), .A1(n2200), .B0(n2216), .B1(
        top_core_KE_CipherKey0_83_), .C0(top_core_KE_n1218), .Y(
        top_core_KE_n1216) );
  OAI2BB2X1 U26635 ( .B0(top_core_KE_n639), .B1(n2229), .A0N(n1632), .A1N(
        top_core_KE_n1219), .Y(top_core_KE_n1218) );
  AOI221X1 U26636 ( .A0(top_core_KE_n1224), .A1(n2200), .B0(n2211), .B1(
        top_core_KE_CipherKey0_82_), .C0(top_core_KE_n1225), .Y(
        top_core_KE_n1223) );
  OAI2BB2X1 U26637 ( .B0(top_core_KE_n640), .B1(n2231), .A0N(n1632), .A1N(
        top_core_KE_n1226), .Y(top_core_KE_n1225) );
  AOI221X1 U26638 ( .A0(top_core_KE_n1231), .A1(n2200), .B0(n2214), .B1(
        top_core_KE_CipherKey0_81_), .C0(top_core_KE_n1232), .Y(
        top_core_KE_n1230) );
  OAI2BB2X1 U26639 ( .B0(top_core_KE_n641), .B1(n2230), .A0N(n1633), .A1N(
        top_core_KE_n1233), .Y(top_core_KE_n1232) );
  AOI221X1 U26640 ( .A0(top_core_KE_n1238), .A1(n2197), .B0(n2215), .B1(
        top_core_KE_CipherKey0_80_), .C0(top_core_KE_n1239), .Y(
        top_core_KE_n1237) );
  OAI2BB2X1 U26641 ( .B0(top_core_KE_n642), .B1(n2232), .A0N(n1632), .A1N(
        top_core_KE_n1240), .Y(top_core_KE_n1239) );
  AOI221X1 U26642 ( .A0(top_core_KE_n1245), .A1(n2203), .B0(n2215), .B1(
        top_core_KE_CipherKey0_79_), .C0(top_core_KE_n1246), .Y(
        top_core_KE_n1244) );
  OAI2BB2X1 U26643 ( .B0(top_core_KE_n643), .B1(n2221), .A0N(n1632), .A1N(
        top_core_KE_n1247), .Y(top_core_KE_n1246) );
  AOI221X1 U26644 ( .A0(top_core_KE_n1252), .A1(n2201), .B0(n2216), .B1(
        top_core_KE_CipherKey0_78_), .C0(top_core_KE_n1253), .Y(
        top_core_KE_n1251) );
  OAI2BB2X1 U26645 ( .B0(top_core_KE_n644), .B1(n2232), .A0N(n1633), .A1N(
        top_core_KE_n1254), .Y(top_core_KE_n1253) );
  AOI221X1 U26646 ( .A0(top_core_KE_n1259), .A1(n2201), .B0(n2216), .B1(
        top_core_KE_CipherKey0_77_), .C0(top_core_KE_n1260), .Y(
        top_core_KE_n1258) );
  OAI2BB2X1 U26647 ( .B0(top_core_KE_n645), .B1(n2233), .A0N(n1632), .A1N(
        top_core_KE_n1261), .Y(top_core_KE_n1260) );
  AOI221X1 U26648 ( .A0(top_core_KE_n1266), .A1(n2201), .B0(n2216), .B1(
        top_core_KE_CipherKey0_76_), .C0(top_core_KE_n1267), .Y(
        top_core_KE_n1265) );
  OAI2BB2X1 U26649 ( .B0(top_core_KE_n646), .B1(n2234), .A0N(n1632), .A1N(
        top_core_KE_n1268), .Y(top_core_KE_n1267) );
  AOI221X1 U26650 ( .A0(top_core_KE_n1273), .A1(n2202), .B0(n2217), .B1(
        top_core_KE_CipherKey0_75_), .C0(top_core_KE_n1274), .Y(
        top_core_KE_n1272) );
  OAI2BB2X1 U26651 ( .B0(top_core_KE_n647), .B1(n2231), .A0N(n1632), .A1N(
        top_core_KE_n1275), .Y(top_core_KE_n1274) );
  AOI221X1 U26652 ( .A0(top_core_KE_n1280), .A1(n2202), .B0(n2217), .B1(
        top_core_KE_CipherKey0_74_), .C0(top_core_KE_n1281), .Y(
        top_core_KE_n1279) );
  OAI2BB2X1 U26653 ( .B0(top_core_KE_n648), .B1(n2231), .A0N(n1632), .A1N(
        top_core_KE_n1282), .Y(top_core_KE_n1281) );
  AOI221X1 U26654 ( .A0(top_core_KE_n1287), .A1(n2202), .B0(n2217), .B1(
        top_core_KE_CipherKey0_73_), .C0(top_core_KE_n1288), .Y(
        top_core_KE_n1286) );
  OAI2BB2X1 U26655 ( .B0(top_core_KE_n649), .B1(n2229), .A0N(n1632), .A1N(
        top_core_KE_n1289), .Y(top_core_KE_n1288) );
  AOI221X1 U26656 ( .A0(top_core_KE_n1294), .A1(n2198), .B0(n2218), .B1(
        top_core_KE_CipherKey0_72_), .C0(top_core_KE_n1295), .Y(
        top_core_KE_n1293) );
  OAI2BB2X1 U26657 ( .B0(top_core_KE_n650), .B1(n2231), .A0N(n1633), .A1N(
        top_core_KE_n1296), .Y(top_core_KE_n1295) );
  AOI221X1 U26658 ( .A0(top_core_KE_n1301), .A1(n2201), .B0(n2218), .B1(
        top_core_KE_CipherKey0_71_), .C0(top_core_KE_n1302), .Y(
        top_core_KE_n1300) );
  OAI2BB2X1 U26659 ( .B0(top_core_KE_n651), .B1(n2235), .A0N(n1632), .A1N(
        top_core_KE_n1303), .Y(top_core_KE_n1302) );
  AOI221X1 U26660 ( .A0(top_core_KE_n1308), .A1(n2201), .B0(n2218), .B1(
        top_core_KE_CipherKey0_70_), .C0(top_core_KE_n1309), .Y(
        top_core_KE_n1307) );
  OAI2BB2X1 U26661 ( .B0(top_core_KE_n652), .B1(n2221), .A0N(n1632), .A1N(
        top_core_KE_n1310), .Y(top_core_KE_n1309) );
  AOI221X1 U26662 ( .A0(top_core_KE_n1315), .A1(n2203), .B0(n2218), .B1(
        top_core_KE_CipherKey0_69_), .C0(top_core_KE_n1316), .Y(
        top_core_KE_n1314) );
  OAI2BB2X1 U26663 ( .B0(top_core_KE_n653), .B1(n2221), .A0N(n1629), .A1N(
        top_core_KE_n1317), .Y(top_core_KE_n1316) );
  AOI221X1 U26664 ( .A0(top_core_KE_n1322), .A1(n2203), .B0(n2214), .B1(
        top_core_KE_CipherKey0_68_), .C0(top_core_KE_n1323), .Y(
        top_core_KE_n1321) );
  OAI2BB2X1 U26665 ( .B0(top_core_KE_n654), .B1(n2232), .A0N(n1632), .A1N(
        top_core_KE_n1324), .Y(top_core_KE_n1323) );
  AOI221X1 U26666 ( .A0(top_core_KE_n1329), .A1(n2203), .B0(n2212), .B1(
        top_core_KE_CipherKey0_67_), .C0(top_core_KE_n1330), .Y(
        top_core_KE_n1328) );
  OAI2BB2X1 U26667 ( .B0(top_core_KE_n655), .B1(n2232), .A0N(n1630), .A1N(
        top_core_KE_n1331), .Y(top_core_KE_n1330) );
  AOI221X1 U26668 ( .A0(top_core_KE_n1336), .A1(n2200), .B0(n2219), .B1(
        top_core_KE_CipherKey0_66_), .C0(top_core_KE_n1337), .Y(
        top_core_KE_n1335) );
  OAI2BB2X1 U26669 ( .B0(top_core_KE_n656), .B1(n2232), .A0N(n1633), .A1N(
        top_core_KE_n1338), .Y(top_core_KE_n1337) );
  AOI221X1 U26670 ( .A0(top_core_KE_n1343), .A1(n2196), .B0(n2219), .B1(
        top_core_KE_CipherKey0_65_), .C0(top_core_KE_n1344), .Y(
        top_core_KE_n1342) );
  OAI2BB2X1 U26671 ( .B0(top_core_KE_n657), .B1(n2229), .A0N(n1628), .A1N(
        top_core_KE_n1345), .Y(top_core_KE_n1344) );
  AOI221X1 U26672 ( .A0(top_core_KE_n1350), .A1(n2196), .B0(n2217), .B1(
        top_core_KE_CipherKey0_64_), .C0(top_core_KE_n1351), .Y(
        top_core_KE_n1349) );
  OAI2BB2X1 U26673 ( .B0(top_core_KE_n658), .B1(n2231), .A0N(n1632), .A1N(
        top_core_KE_n1352), .Y(top_core_KE_n1351) );
  XNOR2X1 U26674 ( .A(top_core_Key[113]), .B(top_core_EC_round_result_9_), .Y(
        n768) );
  XNOR2X1 U26675 ( .A(top_core_Key[120]), .B(top_core_EC_round_result_0_), .Y(
        n769) );
  XNOR2X1 U26676 ( .A(top_core_Key[82]), .B(top_core_EC_round_result_42_), .Y(
        n770) );
  XNOR2X1 U26677 ( .A(top_core_Key[121]), .B(top_core_EC_round_result_1_), .Y(
        n771) );
  XNOR2X1 U26678 ( .A(top_core_Key[41]), .B(top_core_EC_round_result_81_), .Y(
        n772) );
  XNOR2X1 U26679 ( .A(top_core_Key[9]), .B(top_core_EC_round_result_113_), .Y(
        n773) );
  XNOR2X1 U26680 ( .A(top_core_Key[89]), .B(top_core_EC_round_result_33_), .Y(
        n774) );
  XNOR2X1 U26681 ( .A(top_core_Key[40]), .B(top_core_EC_round_result_80_), .Y(
        n775) );
  XNOR2X1 U26682 ( .A(top_core_Key[50]), .B(top_core_EC_round_result_74_), .Y(
        n776) );
  XNOR2X1 U26683 ( .A(top_core_Key[8]), .B(top_core_EC_round_result_112_), .Y(
        n777) );
  XNOR2X1 U26684 ( .A(top_core_Key[88]), .B(top_core_EC_round_result_32_), .Y(
        n778) );
  XNOR2X1 U26685 ( .A(top_core_Key[2]), .B(top_core_EC_round_result_122_), .Y(
        n779) );
  XNOR2X1 U26686 ( .A(top_core_Key[122]), .B(top_core_EC_round_result_2_), .Y(
        n780) );
  XNOR2X1 U26687 ( .A(top_core_Key[65]), .B(top_core_EC_round_result_57_), .Y(
        n781) );
  XNOR2X1 U26688 ( .A(top_core_Key[42]), .B(top_core_EC_round_result_82_), .Y(
        n782) );
  XNOR2X1 U26689 ( .A(top_core_Key[10]), .B(top_core_EC_round_result_114_), 
        .Y(n783) );
  XNOR2X1 U26690 ( .A(top_core_Key[90]), .B(top_core_EC_round_result_34_), .Y(
        n784) );
  XNOR2X1 U26691 ( .A(top_core_Key[98]), .B(top_core_EC_round_result_26_), .Y(
        n785) );
  XNOR2X1 U26692 ( .A(top_core_Key[33]), .B(top_core_EC_round_result_89_), .Y(
        n786) );
  XNOR2X1 U26693 ( .A(top_core_Key[58]), .B(top_core_EC_round_result_66_), .Y(
        n787) );
  XNOR2X1 U26694 ( .A(top_core_Key[57]), .B(top_core_EC_round_result_65_), .Y(
        n788) );
  XNOR2X1 U26695 ( .A(top_core_Key[106]), .B(top_core_EC_round_result_18_), 
        .Y(n789) );
  XNOR2X1 U26696 ( .A(top_core_Key[105]), .B(top_core_EC_round_result_17_), 
        .Y(n790) );
  XNOR2X1 U26697 ( .A(top_core_Key[1]), .B(top_core_EC_round_result_121_), .Y(
        n791) );
  XNOR2X1 U26698 ( .A(top_core_Key[26]), .B(top_core_EC_round_result_98_), .Y(
        n792) );
  XNOR2X1 U26699 ( .A(top_core_Key[25]), .B(top_core_EC_round_result_97_), .Y(
        n793) );
  XNOR2X1 U26700 ( .A(top_core_Key[74]), .B(top_core_EC_round_result_50_), .Y(
        n794) );
  XNOR2X1 U26701 ( .A(top_core_Key[73]), .B(top_core_EC_round_result_49_), .Y(
        n795) );
  XNOR2X1 U26702 ( .A(top_core_Key[34]), .B(top_core_EC_round_result_90_), .Y(
        n796) );
  XNOR2X1 U26703 ( .A(top_core_Key[97]), .B(top_core_EC_round_result_25_), .Y(
        n797) );
  XNOR2X1 U26704 ( .A(top_core_Key[16]), .B(top_core_EC_round_result_104_), 
        .Y(n798) );
  XNOR2X1 U26705 ( .A(top_core_Key[80]), .B(top_core_EC_round_result_40_), .Y(
        n799) );
  XNOR2X1 U26706 ( .A(top_core_Key[17]), .B(top_core_EC_round_result_105_), 
        .Y(n800) );
  XNOR2X1 U26707 ( .A(top_core_Key[45]), .B(top_core_EC_round_result_85_), .Y(
        n801) );
  XNOR2X1 U26708 ( .A(top_core_Key[44]), .B(top_core_EC_round_result_84_), .Y(
        n802) );
  XNOR2X1 U26709 ( .A(top_core_Key[64]), .B(top_core_EC_round_result_56_), .Y(
        n803) );
  XNOR2X1 U26710 ( .A(top_core_Key[81]), .B(top_core_EC_round_result_41_), .Y(
        n804) );
  XNOR2X1 U26711 ( .A(top_core_Key[125]), .B(top_core_EC_round_result_5_), .Y(
        n805) );
  XNOR2X1 U26712 ( .A(top_core_Key[124]), .B(top_core_EC_round_result_4_), .Y(
        n806) );
  XNOR2X1 U26713 ( .A(top_core_Key[0]), .B(top_core_EC_round_result_120_), .Y(
        n807) );
  XNOR2X1 U26714 ( .A(top_core_Key[112]), .B(top_core_EC_round_result_8_), .Y(
        n808) );
  XNOR2X1 U26715 ( .A(top_core_Key[48]), .B(top_core_EC_round_result_72_), .Y(
        n809) );
  XNOR2X1 U26716 ( .A(top_core_Key[49]), .B(top_core_EC_round_result_73_), .Y(
        n810) );
  XNOR2X1 U26717 ( .A(top_core_Key[13]), .B(top_core_EC_round_result_117_), 
        .Y(n811) );
  XNOR2X1 U26718 ( .A(top_core_Key[12]), .B(top_core_EC_round_result_116_), 
        .Y(n812) );
  XNOR2X1 U26719 ( .A(top_core_Key[93]), .B(top_core_EC_round_result_37_), .Y(
        n813) );
  XNOR2X1 U26720 ( .A(top_core_Key[92]), .B(top_core_EC_round_result_36_), .Y(
        n814) );
  XNOR2X1 U26721 ( .A(top_core_Key[96]), .B(top_core_EC_round_result_24_), .Y(
        n815) );
  XNOR2X1 U26722 ( .A(top_core_Key[56]), .B(top_core_EC_round_result_64_), .Y(
        n816) );
  XNOR2X1 U26723 ( .A(top_core_Key[104]), .B(top_core_EC_round_result_16_), 
        .Y(n817) );
  XNOR2X1 U26724 ( .A(top_core_Key[24]), .B(top_core_EC_round_result_96_), .Y(
        n818) );
  XNOR2X1 U26725 ( .A(top_core_Key[72]), .B(top_core_EC_round_result_48_), .Y(
        n819) );
  XNOR2X1 U26726 ( .A(top_core_Key[32]), .B(top_core_EC_round_result_88_), .Y(
        n820) );
  XNOR2X1 U26727 ( .A(top_core_Key[18]), .B(top_core_EC_round_result_106_), 
        .Y(n821) );
  XNOR2X1 U26728 ( .A(top_core_Key[85]), .B(top_core_EC_round_result_45_), .Y(
        n822) );
  XNOR2X1 U26729 ( .A(top_core_Key[84]), .B(top_core_EC_round_result_44_), .Y(
        n823) );
  XNOR2X1 U26730 ( .A(top_core_Key[66]), .B(top_core_EC_round_result_58_), .Y(
        n824) );
  XNOR2X1 U26731 ( .A(top_core_Key[114]), .B(top_core_EC_round_result_10_), 
        .Y(n825) );
  XNOR2X1 U26732 ( .A(top_core_Key[126]), .B(top_core_EC_round_result_6_), .Y(
        n826) );
  XNOR2X1 U26733 ( .A(top_core_Key[4]), .B(top_core_EC_round_result_124_), .Y(
        n827) );
  XNOR2X1 U26734 ( .A(top_core_Key[53]), .B(top_core_EC_round_result_77_), .Y(
        n828) );
  XNOR2X1 U26735 ( .A(top_core_Key[52]), .B(top_core_EC_round_result_76_), .Y(
        n829) );
  XNOR2X1 U26736 ( .A(top_core_Key[5]), .B(top_core_EC_round_result_125_), .Y(
        n830) );
  XNOR2X1 U26737 ( .A(top_core_Key[21]), .B(top_core_EC_round_result_109_), 
        .Y(n831) );
  XNOR2X1 U26738 ( .A(top_core_Key[20]), .B(top_core_EC_round_result_108_), 
        .Y(n832) );
  XNOR2X1 U26739 ( .A(top_core_Key[46]), .B(top_core_EC_round_result_86_), .Y(
        n833) );
  XNOR2X1 U26740 ( .A(top_core_Key[69]), .B(top_core_EC_round_result_61_), .Y(
        n834) );
  XNOR2X1 U26741 ( .A(top_core_Key[117]), .B(top_core_EC_round_result_13_), 
        .Y(n835) );
  XNOR2X1 U26742 ( .A(top_core_Key[14]), .B(top_core_EC_round_result_118_), 
        .Y(n836) );
  XNOR2X1 U26743 ( .A(top_core_Key[94]), .B(top_core_EC_round_result_38_), .Y(
        n837) );
  XNOR2X1 U26744 ( .A(top_core_Key[60]), .B(top_core_EC_round_result_68_), .Y(
        n838) );
  XNOR2X1 U26745 ( .A(top_core_Key[61]), .B(top_core_EC_round_result_69_), .Y(
        n839) );
  XNOR2X1 U26746 ( .A(top_core_Key[108]), .B(top_core_EC_round_result_20_), 
        .Y(n840) );
  XNOR2X1 U26747 ( .A(top_core_Key[109]), .B(top_core_EC_round_result_21_), 
        .Y(n841) );
  XNOR2X1 U26748 ( .A(top_core_Key[28]), .B(top_core_EC_round_result_100_), 
        .Y(n842) );
  XNOR2X1 U26749 ( .A(top_core_Key[29]), .B(top_core_EC_round_result_101_), 
        .Y(n843) );
  XNOR2X1 U26750 ( .A(top_core_Key[76]), .B(top_core_EC_round_result_52_), .Y(
        n844) );
  XNOR2X1 U26751 ( .A(top_core_Key[77]), .B(top_core_EC_round_result_53_), .Y(
        n845) );
  XNOR2X1 U26752 ( .A(top_core_Key[36]), .B(top_core_EC_round_result_92_), .Y(
        n846) );
  XNOR2X1 U26753 ( .A(top_core_Key[86]), .B(top_core_EC_round_result_46_), .Y(
        n847) );
  XNOR2X1 U26754 ( .A(top_core_Key[68]), .B(top_core_EC_round_result_60_), .Y(
        n848) );
  XNOR2X1 U26755 ( .A(top_core_Key[101]), .B(top_core_EC_round_result_29_), 
        .Y(n849) );
  XNOR2X1 U26756 ( .A(top_core_Key[100]), .B(top_core_EC_round_result_28_), 
        .Y(n850) );
  XNOR2X1 U26757 ( .A(top_core_Key[37]), .B(top_core_EC_round_result_93_), .Y(
        n851) );
  XNOR2X1 U26758 ( .A(top_core_Key[116]), .B(top_core_EC_round_result_12_), 
        .Y(n852) );
  XNOR2X1 U26759 ( .A(top_core_Key[54]), .B(top_core_EC_round_result_78_), .Y(
        n853) );
  XNOR2X1 U26760 ( .A(top_core_Key[22]), .B(top_core_EC_round_result_110_), 
        .Y(n854) );
  XNOR2X1 U26761 ( .A(top_core_Key[43]), .B(top_core_EC_round_result_83_), .Y(
        n855) );
  XNOR2X1 U26762 ( .A(top_core_Key[123]), .B(top_core_EC_round_result_3_), .Y(
        n856) );
  XNOR2X1 U26763 ( .A(top_core_Key[70]), .B(top_core_EC_round_result_62_), .Y(
        n857) );
  XNOR2X1 U26764 ( .A(top_core_Key[6]), .B(top_core_EC_round_result_126_), .Y(
        n858) );
  XNOR2X1 U26765 ( .A(top_core_Key[118]), .B(top_core_EC_round_result_14_), 
        .Y(n859) );
  XNOR2X1 U26766 ( .A(top_core_Key[11]), .B(top_core_EC_round_result_115_), 
        .Y(n860) );
  XNOR2X1 U26767 ( .A(top_core_Key[91]), .B(top_core_EC_round_result_35_), .Y(
        n861) );
  XNOR2X1 U26768 ( .A(top_core_Key[62]), .B(top_core_EC_round_result_70_), .Y(
        n862) );
  XNOR2X1 U26769 ( .A(top_core_Key[110]), .B(top_core_EC_round_result_22_), 
        .Y(n863) );
  XNOR2X1 U26770 ( .A(top_core_Key[30]), .B(top_core_EC_round_result_102_), 
        .Y(n864) );
  XNOR2X1 U26771 ( .A(top_core_Key[78]), .B(top_core_EC_round_result_54_), .Y(
        n865) );
  XNOR2X1 U26772 ( .A(top_core_Key[38]), .B(top_core_EC_round_result_94_), .Y(
        n866) );
  XNOR2X1 U26773 ( .A(top_core_Key[102]), .B(top_core_EC_round_result_30_), 
        .Y(n867) );
  XNOR2X1 U26774 ( .A(top_core_Key[83]), .B(top_core_EC_round_result_43_), .Y(
        n868) );
  XNOR2X1 U26775 ( .A(top_core_Key[51]), .B(top_core_EC_round_result_75_), .Y(
        n869) );
  XNOR2X1 U26776 ( .A(top_core_Key[3]), .B(top_core_EC_round_result_123_), .Y(
        n870) );
  XNOR2X1 U26777 ( .A(top_core_Key[99]), .B(top_core_EC_round_result_27_), .Y(
        n871) );
  XNOR2X1 U26778 ( .A(top_core_Key[59]), .B(top_core_EC_round_result_67_), .Y(
        n872) );
  XNOR2X1 U26779 ( .A(top_core_Key[19]), .B(top_core_EC_round_result_107_), 
        .Y(n873) );
  XNOR2X1 U26780 ( .A(top_core_Key[107]), .B(top_core_EC_round_result_19_), 
        .Y(n874) );
  XNOR2X1 U26781 ( .A(top_core_Key[67]), .B(top_core_EC_round_result_59_), .Y(
        n875) );
  XNOR2X1 U26782 ( .A(top_core_Key[27]), .B(top_core_EC_round_result_99_), .Y(
        n876) );
  XNOR2X1 U26783 ( .A(top_core_Key[115]), .B(top_core_EC_round_result_11_), 
        .Y(n877) );
  XNOR2X1 U26784 ( .A(top_core_Key[75]), .B(top_core_EC_round_result_51_), .Y(
        n878) );
  XNOR2X1 U26785 ( .A(top_core_Key[35]), .B(top_core_EC_round_result_91_), .Y(
        n879) );
  XNOR2X1 U26786 ( .A(top_core_Key[127]), .B(top_core_EC_round_result_7_), .Y(
        n880) );
  XNOR2X1 U26787 ( .A(top_core_Key[47]), .B(top_core_EC_round_result_87_), .Y(
        n881) );
  XNOR2X1 U26788 ( .A(top_core_Key[15]), .B(top_core_EC_round_result_119_), 
        .Y(n882) );
  XNOR2X1 U26789 ( .A(top_core_Key[95]), .B(top_core_EC_round_result_39_), .Y(
        n883) );
  XNOR2X1 U26790 ( .A(top_core_Key[63]), .B(top_core_EC_round_result_71_), .Y(
        n884) );
  XNOR2X1 U26791 ( .A(top_core_Key[23]), .B(top_core_EC_round_result_111_), 
        .Y(n885) );
  XNOR2X1 U26792 ( .A(top_core_Key[87]), .B(top_core_EC_round_result_47_), .Y(
        n886) );
  XNOR2X1 U26793 ( .A(top_core_Key[111]), .B(top_core_EC_round_result_23_), 
        .Y(n887) );
  XNOR2X1 U26794 ( .A(top_core_Key[71]), .B(top_core_EC_round_result_63_), .Y(
        n888) );
  XNOR2X1 U26795 ( .A(top_core_Key[7]), .B(top_core_EC_round_result_127_), .Y(
        n889) );
  XNOR2X1 U26796 ( .A(top_core_Key[31]), .B(top_core_EC_round_result_103_), 
        .Y(n890) );
  XNOR2X1 U26797 ( .A(top_core_Key[119]), .B(top_core_EC_round_result_15_), 
        .Y(n891) );
  XNOR2X1 U26798 ( .A(top_core_Key[55]), .B(top_core_EC_round_result_79_), .Y(
        n892) );
  XNOR2X1 U26799 ( .A(top_core_Key[79]), .B(top_core_EC_round_result_55_), .Y(
        n893) );
  XNOR2X1 U26800 ( .A(top_core_Key[39]), .B(top_core_EC_round_result_95_), .Y(
        n894) );
  XNOR2X1 U26801 ( .A(top_core_Key[103]), .B(top_core_EC_round_result_31_), 
        .Y(n895) );
  XOR2X1 U26802 ( .A(n7248), .B(n3973), .Y(top_core_EC_n866) );
  AOI21X1 U26803 ( .A0(n7247), .A1(top_core_EC_rounds_3_), .B0(
        top_core_EC_N577), .Y(n7248) );
  XNOR2X1 U26804 ( .A(top_core_EC_N575), .B(n3985), .Y(top_core_EC_n867) );
  AOI222X1 U26806 ( .A0(top_core_KE_CipherKey0_183_), .A1(n2168), .B0(n2173), 
        .B1(top_core_KE_n969), .C0(top_core_KE_prev_key1_reg_119_), .C1(n2180), 
        .Y(top_core_KE_n968) );
  AOI222X1 U26807 ( .A0(top_core_KE_CipherKey0_182_), .A1(n2168), .B0(n2179), 
        .B1(top_core_KE_n976), .C0(top_core_KE_prev_key1_reg_118_), .C1(n2180), 
        .Y(top_core_KE_n975) );
  AOI222X1 U26808 ( .A0(top_core_KE_CipherKey0_181_), .A1(n2168), .B0(n2178), 
        .B1(top_core_KE_n983), .C0(top_core_KE_prev_key1_reg_117_), .C1(n2180), 
        .Y(top_core_KE_n982) );
  AOI222X1 U26809 ( .A0(top_core_KE_CipherKey0_180_), .A1(n2168), .B0(n2172), 
        .B1(top_core_KE_n990), .C0(top_core_KE_prev_key1_reg_116_), .C1(n2180), 
        .Y(top_core_KE_n989) );
  AOI222X1 U26810 ( .A0(top_core_KE_CipherKey0_179_), .A1(n2168), .B0(n2179), 
        .B1(top_core_KE_n997), .C0(top_core_KE_prev_key1_reg_115_), .C1(n2180), 
        .Y(top_core_KE_n996) );
  AOI222X1 U26811 ( .A0(top_core_KE_CipherKey0_178_), .A1(n2168), .B0(n2179), 
        .B1(top_core_KE_n1004), .C0(top_core_KE_prev_key1_reg_114_), .C1(n2181), .Y(top_core_KE_n1003) );
  AOI222X1 U26812 ( .A0(top_core_KE_CipherKey0_177_), .A1(n2168), .B0(n2179), 
        .B1(top_core_KE_n1011), .C0(top_core_KE_prev_key1_reg_113_), .C1(n2181), .Y(top_core_KE_n1010) );
  AOI222X1 U26813 ( .A0(top_core_KE_CipherKey0_176_), .A1(n2168), .B0(n2179), 
        .B1(top_core_KE_n1018), .C0(top_core_KE_prev_key1_reg_112_), .C1(n2181), .Y(top_core_KE_n1017) );
  AOI222X1 U26814 ( .A0(top_core_KE_CipherKey0_175_), .A1(n2168), .B0(n2179), 
        .B1(top_core_KE_n1025), .C0(top_core_KE_prev_key1_reg_111_), .C1(n2181), .Y(top_core_KE_n1024) );
  AOI222X1 U26815 ( .A0(top_core_KE_CipherKey0_174_), .A1(n2168), .B0(n2179), 
        .B1(top_core_KE_n1032), .C0(top_core_KE_prev_key1_reg_110_), .C1(n2181), .Y(top_core_KE_n1031) );
  AOI222X1 U26816 ( .A0(top_core_KE_CipherKey0_173_), .A1(n2168), .B0(n2179), 
        .B1(top_core_KE_n1039), .C0(top_core_KE_prev_key1_reg_109_), .C1(n2181), .Y(top_core_KE_n1038) );
  AOI222X1 U26817 ( .A0(top_core_KE_CipherKey0_172_), .A1(n2168), .B0(n2179), 
        .B1(top_core_KE_n1046), .C0(top_core_KE_prev_key1_reg_108_), .C1(n2181), .Y(top_core_KE_n1045) );
  AOI222X1 U26818 ( .A0(top_core_KE_CipherKey0_171_), .A1(n2167), .B0(n2179), 
        .B1(top_core_KE_n1053), .C0(top_core_KE_prev_key1_reg_107_), .C1(n2181), .Y(top_core_KE_n1052) );
  AOI222X1 U26819 ( .A0(top_core_KE_CipherKey0_170_), .A1(n2167), .B0(n2179), 
        .B1(top_core_KE_n1060), .C0(top_core_KE_prev_key1_reg_106_), .C1(n2181), .Y(top_core_KE_n1059) );
  AOI222X1 U26820 ( .A0(top_core_KE_CipherKey0_169_), .A1(n2167), .B0(n2179), 
        .B1(top_core_KE_n1067), .C0(top_core_KE_prev_key1_reg_105_), .C1(n2181), .Y(top_core_KE_n1066) );
  AOI222X1 U26821 ( .A0(top_core_KE_CipherKey0_168_), .A1(n2167), .B0(n2179), 
        .B1(top_core_KE_n1074), .C0(top_core_KE_prev_key1_reg_104_), .C1(n2181), .Y(top_core_KE_n1073) );
  AOI222X1 U26822 ( .A0(top_core_KE_CipherKey0_167_), .A1(n2167), .B0(n2179), 
        .B1(top_core_KE_n1081), .C0(top_core_KE_prev_key1_reg_103_), .C1(n2181), .Y(top_core_KE_n1080) );
  AOI222X1 U26823 ( .A0(top_core_KE_CipherKey0_166_), .A1(n2167), .B0(n2178), 
        .B1(top_core_KE_n1088), .C0(top_core_KE_prev_key1_reg_102_), .C1(n2183), .Y(top_core_KE_n1087) );
  AOI222X1 U26824 ( .A0(top_core_KE_CipherKey0_165_), .A1(n2167), .B0(n2178), 
        .B1(top_core_KE_n1095), .C0(top_core_KE_prev_key1_reg_101_), .C1(n2184), .Y(top_core_KE_n1094) );
  AOI222X1 U26825 ( .A0(top_core_KE_CipherKey0_164_), .A1(n2167), .B0(n2178), 
        .B1(top_core_KE_n1102), .C0(top_core_KE_prev_key1_reg_100_), .C1(n2185), .Y(top_core_KE_n1101) );
  AOI222X1 U26826 ( .A0(top_core_KE_CipherKey0_163_), .A1(n2167), .B0(n2178), 
        .B1(top_core_KE_n1109), .C0(top_core_KE_prev_key1_reg_99_), .C1(n2187), 
        .Y(top_core_KE_n1108) );
  AOI222X1 U26827 ( .A0(top_core_KE_CipherKey0_162_), .A1(n2167), .B0(n2178), 
        .B1(top_core_KE_n1116), .C0(top_core_KE_prev_key1_reg_98_), .C1(n2186), 
        .Y(top_core_KE_n1115) );
  AOI222X1 U26828 ( .A0(top_core_KE_CipherKey0_161_), .A1(n2167), .B0(n2178), 
        .B1(top_core_KE_n1123), .C0(top_core_KE_prev_key1_reg_97_), .C1(n2182), 
        .Y(top_core_KE_n1122) );
  AOI222X1 U26829 ( .A0(top_core_KE_CipherKey0_160_), .A1(n2167), .B0(n2178), 
        .B1(top_core_KE_n1130), .C0(top_core_KE_prev_key1_reg_96_), .C1(n2180), 
        .Y(top_core_KE_n1129) );
  AOI222X1 U26830 ( .A0(top_core_KE_CipherKey0_191_), .A1(top_core_KE_n907), 
        .B0(n2177), .B1(top_core_KE_n909), .C0(n2183), .C1(
        top_core_KE_prev_key1_reg_127_), .Y(top_core_KE_n906) );
  AOI222X1 U26831 ( .A0(top_core_KE_CipherKey0_190_), .A1(top_core_KE_n907), 
        .B0(n2174), .B1(top_core_KE_n920), .C0(top_core_KE_prev_key1_reg_126_), 
        .C1(n2180), .Y(top_core_KE_n919) );
  AOI222X1 U26832 ( .A0(top_core_KE_CipherKey0_189_), .A1(top_core_KE_n907), 
        .B0(n2176), .B1(top_core_KE_n927), .C0(top_core_KE_prev_key1_reg_125_), 
        .C1(n2180), .Y(top_core_KE_n926) );
  AOI222X1 U26833 ( .A0(top_core_KE_CipherKey0_188_), .A1(top_core_KE_n907), 
        .B0(n2175), .B1(top_core_KE_n934), .C0(top_core_KE_prev_key1_reg_124_), 
        .C1(n2180), .Y(top_core_KE_n933) );
  AOI222X1 U26834 ( .A0(top_core_KE_CipherKey0_187_), .A1(top_core_KE_n907), 
        .B0(n2171), .B1(top_core_KE_n941), .C0(top_core_KE_prev_key1_reg_123_), 
        .C1(n2180), .Y(top_core_KE_n940) );
  AOI222X1 U26835 ( .A0(top_core_KE_CipherKey0_186_), .A1(top_core_KE_n907), 
        .B0(n2173), .B1(top_core_KE_n948), .C0(top_core_KE_prev_key1_reg_122_), 
        .C1(n2180), .Y(top_core_KE_n947) );
  AOI222X1 U26836 ( .A0(top_core_KE_CipherKey0_185_), .A1(top_core_KE_n907), 
        .B0(n2179), .B1(top_core_KE_n955), .C0(top_core_KE_prev_key1_reg_121_), 
        .C1(n2180), .Y(top_core_KE_n954) );
  AOI222X1 U26837 ( .A0(top_core_KE_CipherKey0_184_), .A1(top_core_KE_n907), 
        .B0(n2178), .B1(top_core_KE_n962), .C0(top_core_KE_prev_key1_reg_120_), 
        .C1(n2180), .Y(top_core_KE_n961) );
  AOI222X1 U26838 ( .A0(top_core_KE_CipherKey0_119_), .A1(n2163), .B0(n2175), 
        .B1(top_core_KE_n1425), .C0(n2184), .C1(top_core_KE_n1426), .Y(
        top_core_KE_n1424) );
  AOI222X1 U26839 ( .A0(top_core_KE_CipherKey0_118_), .A1(n2163), .B0(n2175), 
        .B1(top_core_KE_n1433), .C0(n2184), .C1(top_core_KE_n1434), .Y(
        top_core_KE_n1432) );
  AOI222X1 U26840 ( .A0(top_core_KE_CipherKey0_117_), .A1(n2163), .B0(n2175), 
        .B1(top_core_KE_n1441), .C0(n2184), .C1(top_core_KE_n1442), .Y(
        top_core_KE_n1440) );
  AOI222X1 U26841 ( .A0(top_core_KE_CipherKey0_116_), .A1(n2163), .B0(n2175), 
        .B1(top_core_KE_n1449), .C0(n2184), .C1(top_core_KE_n1450), .Y(
        top_core_KE_n1448) );
  AOI222X1 U26842 ( .A0(top_core_KE_CipherKey0_115_), .A1(n2163), .B0(n2175), 
        .B1(top_core_KE_n1457), .C0(n2184), .C1(top_core_KE_n1458), .Y(
        top_core_KE_n1456) );
  AOI222X1 U26843 ( .A0(top_core_KE_CipherKey0_114_), .A1(n2163), .B0(n2174), 
        .B1(top_core_KE_n1465), .C0(n2184), .C1(top_core_KE_n1466), .Y(
        top_core_KE_n1464) );
  AOI222X1 U26844 ( .A0(top_core_KE_CipherKey0_113_), .A1(n2163), .B0(n2174), 
        .B1(top_core_KE_n1473), .C0(n2184), .C1(top_core_KE_n1474), .Y(
        top_core_KE_n1472) );
  AOI222X1 U26845 ( .A0(top_core_KE_CipherKey0_112_), .A1(n2163), .B0(n2174), 
        .B1(top_core_KE_n1481), .C0(n2184), .C1(top_core_KE_n1482), .Y(
        top_core_KE_n1480) );
  AOI222X1 U26846 ( .A0(top_core_KE_CipherKey0_111_), .A1(n2162), .B0(n2174), 
        .B1(top_core_KE_n1489), .C0(n2184), .C1(top_core_KE_n1490), .Y(
        top_core_KE_n1488) );
  AOI222X1 U26847 ( .A0(top_core_KE_CipherKey0_110_), .A1(n2162), .B0(n2174), 
        .B1(top_core_KE_n1497), .C0(n2184), .C1(top_core_KE_n1498), .Y(
        top_core_KE_n1496) );
  AOI222X1 U26848 ( .A0(top_core_KE_CipherKey0_109_), .A1(n2162), .B0(n2174), 
        .B1(top_core_KE_n1505), .C0(n2184), .C1(top_core_KE_n1506), .Y(
        top_core_KE_n1504) );
  AOI222X1 U26849 ( .A0(top_core_KE_CipherKey0_108_), .A1(n2162), .B0(n2174), 
        .B1(top_core_KE_n1513), .C0(n2184), .C1(top_core_KE_n1514), .Y(
        top_core_KE_n1512) );
  AOI222X1 U26850 ( .A0(top_core_KE_CipherKey0_107_), .A1(n2162), .B0(n2174), 
        .B1(top_core_KE_n1521), .C0(n2184), .C1(top_core_KE_n1522), .Y(
        top_core_KE_n1520) );
  AOI222X1 U26851 ( .A0(top_core_KE_CipherKey0_106_), .A1(n2162), .B0(n2174), 
        .B1(top_core_KE_n1529), .C0(n2185), .C1(top_core_KE_n1530), .Y(
        top_core_KE_n1528) );
  AOI222X1 U26852 ( .A0(top_core_KE_CipherKey0_105_), .A1(n2162), .B0(n2174), 
        .B1(top_core_KE_n1537), .C0(n2185), .C1(top_core_KE_n1538), .Y(
        top_core_KE_n1536) );
  AOI222X1 U26853 ( .A0(top_core_KE_CipherKey0_104_), .A1(n2162), .B0(n2174), 
        .B1(top_core_KE_n1545), .C0(n2185), .C1(top_core_KE_n1546), .Y(
        top_core_KE_n1544) );
  AOI222X1 U26854 ( .A0(top_core_KE_CipherKey0_103_), .A1(n2162), .B0(n2174), 
        .B1(top_core_KE_n1553), .C0(n2185), .C1(top_core_KE_n1554), .Y(
        top_core_KE_n1552) );
  AOI222X1 U26855 ( .A0(top_core_KE_CipherKey0_102_), .A1(n2162), .B0(n2174), 
        .B1(top_core_KE_n1561), .C0(n2185), .C1(top_core_KE_n1562), .Y(
        top_core_KE_n1560) );
  AOI222X1 U26856 ( .A0(top_core_KE_CipherKey0_101_), .A1(n2162), .B0(n2173), 
        .B1(top_core_KE_n1569), .C0(n2185), .C1(top_core_KE_n1570), .Y(
        top_core_KE_n1568) );
  AOI222X1 U26857 ( .A0(top_core_KE_CipherKey0_100_), .A1(n2162), .B0(n2173), 
        .B1(top_core_KE_n1577), .C0(n2185), .C1(top_core_KE_n1578), .Y(
        top_core_KE_n1576) );
  AOI222X1 U26858 ( .A0(top_core_KE_CipherKey0_99_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1585), .C0(n2185), .C1(top_core_KE_n1586), .Y(
        top_core_KE_n1584) );
  AOI222X1 U26859 ( .A0(top_core_KE_CipherKey0_98_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1593), .C0(n2185), .C1(top_core_KE_n1594), .Y(
        top_core_KE_n1592) );
  AOI222X1 U26860 ( .A0(top_core_KE_CipherKey0_97_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1601), .C0(n2185), .C1(top_core_KE_n1602), .Y(
        top_core_KE_n1600) );
  AOI222X1 U26861 ( .A0(top_core_KE_CipherKey0_96_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1609), .C0(n2185), .C1(top_core_KE_n1610), .Y(
        top_core_KE_n1608) );
  AOI222X1 U26862 ( .A0(top_core_KE_CipherKey0_159_), .A1(n2166), .B0(n2178), 
        .B1(top_core_KE_n1137), .C0(n1341), .C1(n2181), .Y(top_core_KE_n1136)
         );
  AOI222X1 U26863 ( .A0(top_core_KE_CipherKey0_158_), .A1(n2166), .B0(n2178), 
        .B1(top_core_KE_n1144), .C0(n1369), .C1(n2183), .Y(top_core_KE_n1143)
         );
  AOI222X1 U26864 ( .A0(top_core_KE_CipherKey0_157_), .A1(n2166), .B0(n2178), 
        .B1(top_core_KE_n1151), .C0(n1637), .C1(n2184), .Y(top_core_KE_n1150)
         );
  AOI222X1 U26865 ( .A0(top_core_KE_CipherKey0_156_), .A1(n2166), .B0(n2178), 
        .B1(top_core_KE_n1158), .C0(n1365), .C1(n2185), .Y(top_core_KE_n1157)
         );
  AOI222X1 U26866 ( .A0(top_core_KE_CipherKey0_155_), .A1(n2166), .B0(n2178), 
        .B1(top_core_KE_n1165), .C0(n1361), .C1(n2187), .Y(top_core_KE_n1164)
         );
  AOI222X1 U26867 ( .A0(top_core_KE_CipherKey0_154_), .A1(n2166), .B0(n2178), 
        .B1(top_core_KE_n1172), .C0(n1647), .C1(n2182), .Y(top_core_KE_n1171)
         );
  AOI222X1 U26868 ( .A0(top_core_KE_CipherKey0_153_), .A1(n2166), .B0(n2177), 
        .B1(top_core_KE_n1179), .C0(n1652), .C1(n2182), .Y(top_core_KE_n1178)
         );
  AOI222X1 U26869 ( .A0(top_core_KE_CipherKey0_152_), .A1(n2166), .B0(n2177), 
        .B1(top_core_KE_n1186), .C0(n1659), .C1(n2182), .Y(top_core_KE_n1185)
         );
  AOI222X1 U26870 ( .A0(top_core_KE_CipherKey0_151_), .A1(n2166), .B0(n2177), 
        .B1(top_core_KE_n1193), .C0(n1340), .C1(n2182), .Y(top_core_KE_n1192)
         );
  AOI222X1 U26871 ( .A0(top_core_KE_CipherKey0_150_), .A1(n2166), .B0(n2177), 
        .B1(top_core_KE_n1200), .C0(n1356), .C1(n2182), .Y(top_core_KE_n1199)
         );
  AOI222X1 U26872 ( .A0(top_core_KE_CipherKey0_149_), .A1(n2166), .B0(n2177), 
        .B1(top_core_KE_n1207), .C0(n1667), .C1(n2182), .Y(top_core_KE_n1206)
         );
  AOI222X1 U26873 ( .A0(top_core_KE_CipherKey0_148_), .A1(n2166), .B0(n2177), 
        .B1(top_core_KE_n1214), .C0(n1367), .C1(n2182), .Y(top_core_KE_n1213)
         );
  AOI222X1 U26874 ( .A0(top_core_KE_CipherKey0_147_), .A1(n2165), .B0(n2177), 
        .B1(top_core_KE_n1221), .C0(n1363), .C1(n2182), .Y(top_core_KE_n1220)
         );
  AOI222X1 U26875 ( .A0(top_core_KE_CipherKey0_146_), .A1(n2165), .B0(n2177), 
        .B1(top_core_KE_n1228), .C0(n1674), .C1(n2182), .Y(top_core_KE_n1227)
         );
  AOI222X1 U26876 ( .A0(top_core_KE_CipherKey0_145_), .A1(n2165), .B0(n2177), 
        .B1(top_core_KE_n1235), .C0(n1681), .C1(n2182), .Y(top_core_KE_n1234)
         );
  AOI222X1 U26877 ( .A0(top_core_KE_CipherKey0_144_), .A1(n2165), .B0(n2177), 
        .B1(top_core_KE_n1242), .C0(n1688), .C1(n2182), .Y(top_core_KE_n1241)
         );
  AOI222X1 U26878 ( .A0(top_core_KE_CipherKey0_143_), .A1(n2165), .B0(n2177), 
        .B1(top_core_KE_n1249), .C0(n1337), .C1(n2182), .Y(top_core_KE_n1248)
         );
  AOI222X1 U26879 ( .A0(top_core_KE_CipherKey0_142_), .A1(n2165), .B0(n2177), 
        .B1(top_core_KE_n1256), .C0(n1355), .C1(top_core_KE_n910), .Y(
        top_core_KE_n1255) );
  AOI222X1 U26880 ( .A0(top_core_KE_CipherKey0_141_), .A1(n2165), .B0(n2177), 
        .B1(top_core_KE_n1263), .C0(n1696), .C1(top_core_KE_n910), .Y(
        top_core_KE_n1262) );
  AOI222X1 U26881 ( .A0(top_core_KE_CipherKey0_140_), .A1(n2165), .B0(n2176), 
        .B1(top_core_KE_n1270), .C0(n1351), .C1(top_core_KE_n910), .Y(
        top_core_KE_n1269) );
  AOI222X1 U26882 ( .A0(top_core_KE_CipherKey0_139_), .A1(n2165), .B0(n2176), 
        .B1(top_core_KE_n1277), .C0(n1347), .C1(top_core_KE_n910), .Y(
        top_core_KE_n1276) );
  AOI222X1 U26883 ( .A0(top_core_KE_CipherKey0_138_), .A1(n2165), .B0(n2176), 
        .B1(top_core_KE_n1284), .C0(n1703), .C1(top_core_KE_n910), .Y(
        top_core_KE_n1283) );
  AOI222X1 U26884 ( .A0(top_core_KE_CipherKey0_137_), .A1(n2165), .B0(n2176), 
        .B1(top_core_KE_n1291), .C0(n1710), .C1(top_core_KE_n910), .Y(
        top_core_KE_n1290) );
  AOI222X1 U26885 ( .A0(top_core_KE_CipherKey0_136_), .A1(n2165), .B0(n2176), 
        .B1(top_core_KE_n1298), .C0(n1717), .C1(n2182), .Y(top_core_KE_n1297)
         );
  AOI222X1 U26886 ( .A0(top_core_KE_CipherKey0_135_), .A1(n2164), .B0(n2176), 
        .B1(top_core_KE_n1305), .C0(n1336), .C1(n2180), .Y(top_core_KE_n1304)
         );
  AOI222X1 U26887 ( .A0(top_core_KE_CipherKey0_134_), .A1(n2164), .B0(n2176), 
        .B1(top_core_KE_n1312), .C0(n1342), .C1(n2181), .Y(top_core_KE_n1311)
         );
  AOI222X1 U26888 ( .A0(top_core_KE_CipherKey0_133_), .A1(n2164), .B0(n2176), 
        .B1(top_core_KE_n1319), .C0(n1725), .C1(n2181), .Y(top_core_KE_n1318)
         );
  AOI222X1 U26889 ( .A0(top_core_KE_CipherKey0_132_), .A1(n2164), .B0(n2176), 
        .B1(top_core_KE_n1326), .C0(n1353), .C1(n2182), .Y(top_core_KE_n1325)
         );
  AOI222X1 U26890 ( .A0(top_core_KE_CipherKey0_131_), .A1(n2164), .B0(n2176), 
        .B1(top_core_KE_n1333), .C0(n1349), .C1(n2180), .Y(top_core_KE_n1332)
         );
  AOI222X1 U26891 ( .A0(top_core_KE_CipherKey0_130_), .A1(n2164), .B0(n2176), 
        .B1(top_core_KE_n1340), .C0(n1732), .C1(n2183), .Y(top_core_KE_n1339)
         );
  AOI222X1 U26892 ( .A0(top_core_KE_CipherKey0_129_), .A1(n2164), .B0(n2176), 
        .B1(top_core_KE_n1347), .C0(n1739), .C1(n2183), .Y(top_core_KE_n1346)
         );
  AOI222X1 U26893 ( .A0(top_core_KE_CipherKey0_128_), .A1(n2164), .B0(n2176), 
        .B1(top_core_KE_n1354), .C0(n1746), .C1(n2183), .Y(top_core_KE_n1353)
         );
  AOI222X1 U26894 ( .A0(top_core_KE_CipherKey0_127_), .A1(n2164), .B0(n2175), 
        .B1(top_core_KE_n1361), .C0(n2183), .C1(top_core_KE_n1362), .Y(
        top_core_KE_n1360) );
  AOI222X1 U26895 ( .A0(top_core_KE_CipherKey0_126_), .A1(n2164), .B0(n2175), 
        .B1(top_core_KE_n1369), .C0(n2183), .C1(top_core_KE_n1370), .Y(
        top_core_KE_n1368) );
  AOI222X1 U26896 ( .A0(top_core_KE_CipherKey0_125_), .A1(n2164), .B0(n2175), 
        .B1(top_core_KE_n1377), .C0(n2183), .C1(top_core_KE_n1378), .Y(
        top_core_KE_n1376) );
  AOI222X1 U26897 ( .A0(top_core_KE_CipherKey0_124_), .A1(n2164), .B0(n2175), 
        .B1(top_core_KE_n1385), .C0(n2183), .C1(top_core_KE_n1386), .Y(
        top_core_KE_n1384) );
  AOI222X1 U26898 ( .A0(top_core_KE_CipherKey0_123_), .A1(n2163), .B0(n2175), 
        .B1(top_core_KE_n1393), .C0(n2183), .C1(top_core_KE_n1394), .Y(
        top_core_KE_n1392) );
  AOI222X1 U26899 ( .A0(top_core_KE_CipherKey0_122_), .A1(n2163), .B0(n2175), 
        .B1(top_core_KE_n1401), .C0(n2183), .C1(top_core_KE_n1402), .Y(
        top_core_KE_n1400) );
  AOI222X1 U26900 ( .A0(top_core_KE_CipherKey0_121_), .A1(n2163), .B0(n2175), 
        .B1(top_core_KE_n1409), .C0(n2183), .C1(top_core_KE_n1410), .Y(
        top_core_KE_n1408) );
  AOI222X1 U26901 ( .A0(top_core_KE_CipherKey0_120_), .A1(n2163), .B0(n2175), 
        .B1(top_core_KE_n1417), .C0(n2183), .C1(top_core_KE_n1418), .Y(
        top_core_KE_n1416) );
  AOI222X1 U26902 ( .A0(top_core_KE_CipherKey0_95_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1617), .C0(n2185), .C1(top_core_KE_n1618), .Y(
        top_core_KE_n1616) );
  AOI222X1 U26903 ( .A0(top_core_KE_CipherKey0_94_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1625), .C0(n2185), .C1(top_core_KE_n1626), .Y(
        top_core_KE_n1624) );
  AOI222X1 U26904 ( .A0(top_core_KE_CipherKey0_93_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1633), .C0(n2186), .C1(top_core_KE_n1634), .Y(
        top_core_KE_n1632) );
  AOI222X1 U26905 ( .A0(top_core_KE_CipherKey0_92_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1641), .C0(n2186), .C1(top_core_KE_n1642), .Y(
        top_core_KE_n1640) );
  AOI222X1 U26906 ( .A0(top_core_KE_CipherKey0_91_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1649), .C0(n2186), .C1(top_core_KE_n1650), .Y(
        top_core_KE_n1648) );
  AOI222X1 U26907 ( .A0(top_core_KE_CipherKey0_90_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1657), .C0(n2186), .C1(top_core_KE_n1658), .Y(
        top_core_KE_n1656) );
  AOI222X1 U26908 ( .A0(top_core_KE_CipherKey0_89_), .A1(n2161), .B0(n2173), 
        .B1(top_core_KE_n1665), .C0(n2186), .C1(top_core_KE_n1666), .Y(
        top_core_KE_n1664) );
  AOI222X1 U26909 ( .A0(top_core_KE_CipherKey0_88_), .A1(n2161), .B0(n2172), 
        .B1(top_core_KE_n1673), .C0(n2186), .C1(top_core_KE_n1674), .Y(
        top_core_KE_n1672) );
  AOI222X1 U26910 ( .A0(top_core_KE_CipherKey0_87_), .A1(n2163), .B0(n2172), 
        .B1(top_core_KE_n1681), .C0(n2186), .C1(top_core_KE_n1682), .Y(
        top_core_KE_n1680) );
  AOI222X1 U26911 ( .A0(top_core_KE_CipherKey0_86_), .A1(n2168), .B0(n2172), 
        .B1(top_core_KE_n1689), .C0(n2186), .C1(top_core_KE_n1690), .Y(
        top_core_KE_n1688) );
  AOI222X1 U26912 ( .A0(top_core_KE_CipherKey0_85_), .A1(n2167), .B0(n2172), 
        .B1(top_core_KE_n1697), .C0(n2186), .C1(top_core_KE_n1698), .Y(
        top_core_KE_n1696) );
  AOI222X1 U26913 ( .A0(top_core_KE_CipherKey0_84_), .A1(n2165), .B0(n2172), 
        .B1(top_core_KE_n1705), .C0(n2186), .C1(top_core_KE_n1706), .Y(
        top_core_KE_n1704) );
  AOI222X1 U26914 ( .A0(top_core_KE_CipherKey0_83_), .A1(n2161), .B0(n2172), 
        .B1(top_core_KE_n1713), .C0(n2186), .C1(top_core_KE_n1714), .Y(
        top_core_KE_n1712) );
  AOI222X1 U26915 ( .A0(top_core_KE_CipherKey0_82_), .A1(n2162), .B0(n2172), 
        .B1(top_core_KE_n1721), .C0(n2186), .C1(top_core_KE_n1722), .Y(
        top_core_KE_n1720) );
  AOI222X1 U26916 ( .A0(top_core_KE_CipherKey0_81_), .A1(n2166), .B0(n2172), 
        .B1(top_core_KE_n1729), .C0(n2186), .C1(top_core_KE_n1730), .Y(
        top_core_KE_n1728) );
  AOI222X1 U26917 ( .A0(top_core_KE_CipherKey0_80_), .A1(n2164), .B0(n2172), 
        .B1(top_core_KE_n1737), .C0(n2187), .C1(top_core_KE_n1738), .Y(
        top_core_KE_n1736) );
  AOI222X1 U26918 ( .A0(top_core_KE_CipherKey0_79_), .A1(n2163), .B0(n2172), 
        .B1(top_core_KE_n1745), .C0(n2187), .C1(top_core_KE_n1746), .Y(
        top_core_KE_n1744) );
  AOI222X1 U26919 ( .A0(top_core_KE_CipherKey0_78_), .A1(n2168), .B0(n2172), 
        .B1(top_core_KE_n1753), .C0(n2187), .C1(top_core_KE_n1754), .Y(
        top_core_KE_n1752) );
  AOI222X1 U26920 ( .A0(top_core_KE_CipherKey0_77_), .A1(n2167), .B0(n2172), 
        .B1(top_core_KE_n1761), .C0(n2187), .C1(top_core_KE_n1762), .Y(
        top_core_KE_n1760) );
  AOI222X1 U26921 ( .A0(top_core_KE_CipherKey0_76_), .A1(n2165), .B0(n2172), 
        .B1(top_core_KE_n1769), .C0(n2187), .C1(top_core_KE_n1770), .Y(
        top_core_KE_n1768) );
  AOI222X1 U26922 ( .A0(top_core_KE_CipherKey0_75_), .A1(top_core_KE_n907), 
        .B0(n2171), .B1(top_core_KE_n1777), .C0(n2187), .C1(top_core_KE_n1778), 
        .Y(top_core_KE_n1776) );
  AOI222X1 U26923 ( .A0(top_core_KE_CipherKey0_74_), .A1(n2162), .B0(n2171), 
        .B1(top_core_KE_n1785), .C0(n2187), .C1(top_core_KE_n1786), .Y(
        top_core_KE_n1784) );
  AOI222X1 U26924 ( .A0(top_core_KE_CipherKey0_73_), .A1(n2166), .B0(n2171), 
        .B1(top_core_KE_n1793), .C0(n2187), .C1(top_core_KE_n1794), .Y(
        top_core_KE_n1792) );
  AOI222X1 U26925 ( .A0(top_core_KE_CipherKey0_72_), .A1(n2164), .B0(n2171), 
        .B1(top_core_KE_n1801), .C0(n2187), .C1(top_core_KE_n1802), .Y(
        top_core_KE_n1800) );
  AOI222X1 U26926 ( .A0(top_core_KE_CipherKey0_71_), .A1(n2163), .B0(n2171), 
        .B1(top_core_KE_n1809), .C0(n2187), .C1(top_core_KE_n1810), .Y(
        top_core_KE_n1808) );
  AOI222X1 U26927 ( .A0(top_core_KE_CipherKey0_70_), .A1(n2168), .B0(n2171), 
        .B1(top_core_KE_n1817), .C0(n2187), .C1(top_core_KE_n1818), .Y(
        top_core_KE_n1816) );
  AOI222X1 U26928 ( .A0(top_core_KE_CipherKey0_69_), .A1(n2167), .B0(n2171), 
        .B1(top_core_KE_n1825), .C0(n2187), .C1(top_core_KE_n1826), .Y(
        top_core_KE_n1824) );
  AOI222X1 U26929 ( .A0(top_core_KE_CipherKey0_68_), .A1(n2165), .B0(n2171), 
        .B1(top_core_KE_n1833), .C0(n2187), .C1(top_core_KE_n1834), .Y(
        top_core_KE_n1832) );
  AOI222X1 U26930 ( .A0(top_core_KE_CipherKey0_67_), .A1(n2161), .B0(n2171), 
        .B1(top_core_KE_n1841), .C0(top_core_KE_n910), .C1(top_core_KE_n1842), 
        .Y(top_core_KE_n1840) );
  AOI222X1 U26931 ( .A0(top_core_KE_CipherKey0_66_), .A1(n2164), .B0(n2171), 
        .B1(top_core_KE_n1849), .C0(top_core_KE_n910), .C1(top_core_KE_n1850), 
        .Y(top_core_KE_n1848) );
  AOI222X1 U26932 ( .A0(top_core_KE_CipherKey0_65_), .A1(n2162), .B0(n2171), 
        .B1(top_core_KE_n1857), .C0(top_core_KE_n910), .C1(top_core_KE_n1858), 
        .Y(top_core_KE_n1856) );
  AOI222X1 U26933 ( .A0(top_core_KE_CipherKey0_64_), .A1(n2166), .B0(n2171), 
        .B1(top_core_KE_n1868), .C0(n2183), .C1(top_core_KE_n1869), .Y(
        top_core_KE_n1867) );
  AND2X2 U26934 ( .A(top_core_io_n1179), .B(top_core_io_NK_0_), .Y(
        top_core_io_N126) );
  AND2X2 U26935 ( .A(top_core_io_n1180), .B(top_core_io_NK_0_), .Y(
        top_core_io_N125) );
  INVX1 U26936 ( .A(top_core_KE_CipherKey0_126_), .Y(n7117) );
  INVX1 U26937 ( .A(top_core_KE_CipherKey0_125_), .Y(n7116) );
  INVX1 U26938 ( .A(top_core_KE_CipherKey0_124_), .Y(n7115) );
  INVX1 U26939 ( .A(top_core_KE_CipherKey0_123_), .Y(n7114) );
  INVX1 U26940 ( .A(top_core_KE_CipherKey0_122_), .Y(n7113) );
  INVX1 U26941 ( .A(top_core_KE_CipherKey0_121_), .Y(n7112) );
  INVX1 U26942 ( .A(top_core_KE_CipherKey0_120_), .Y(n7111) );
  INVX1 U26943 ( .A(top_core_KE_CipherKey0_111_), .Y(n7110) );
  INVX1 U26944 ( .A(top_core_KE_CipherKey0_110_), .Y(n7109) );
  INVX1 U26945 ( .A(top_core_KE_CipherKey0_109_), .Y(n7108) );
  INVX1 U26946 ( .A(top_core_KE_CipherKey0_108_), .Y(n7107) );
  INVX1 U26947 ( .A(top_core_KE_CipherKey0_107_), .Y(n7106) );
  INVX1 U26948 ( .A(top_core_KE_CipherKey0_106_), .Y(n7105) );
  INVX1 U26949 ( .A(top_core_KE_CipherKey0_105_), .Y(n7104) );
  INVX1 U26950 ( .A(top_core_KE_CipherKey0_104_), .Y(n7103) );
  INVX1 U26951 ( .A(top_core_KE_CipherKey0_103_), .Y(n7102) );
  INVX1 U26952 ( .A(top_core_KE_CipherKey0_102_), .Y(n7101) );
  INVX1 U26953 ( .A(top_core_KE_CipherKey0_101_), .Y(n7100) );
  INVX1 U26954 ( .A(top_core_KE_CipherKey0_100_), .Y(n7099) );
  INVX1 U26955 ( .A(top_core_KE_CipherKey0_99_), .Y(n7098) );
  INVX1 U26956 ( .A(top_core_KE_CipherKey0_98_), .Y(n7097) );
  INVX1 U26957 ( .A(top_core_KE_CipherKey0_97_), .Y(n7096) );
  INVX1 U26958 ( .A(top_core_KE_CipherKey0_96_), .Y(n7095) );
  INVX1 U26959 ( .A(top_core_KE_CipherKey0_95_), .Y(n7094) );
  INVX1 U26960 ( .A(top_core_KE_CipherKey0_94_), .Y(n7093) );
  INVX1 U26961 ( .A(top_core_KE_CipherKey0_93_), .Y(n7092) );
  INVX1 U26962 ( .A(top_core_KE_CipherKey0_92_), .Y(n7091) );
  INVX1 U26963 ( .A(top_core_KE_CipherKey0_91_), .Y(n7090) );
  INVX1 U26964 ( .A(top_core_KE_CipherKey0_90_), .Y(n7089) );
  INVX1 U26965 ( .A(top_core_KE_CipherKey0_89_), .Y(n7088) );
  INVX1 U26966 ( .A(top_core_KE_CipherKey0_88_), .Y(n7087) );
  INVX1 U26967 ( .A(top_core_KE_CipherKey0_191_), .Y(n7181) );
  INVX1 U26968 ( .A(top_core_KE_CipherKey0_190_), .Y(n7180) );
  INVX1 U26969 ( .A(top_core_KE_CipherKey0_189_), .Y(n7179) );
  INVX1 U26970 ( .A(top_core_KE_CipherKey0_188_), .Y(n7178) );
  INVX1 U26971 ( .A(top_core_KE_CipherKey0_187_), .Y(n7177) );
  INVX1 U26972 ( .A(top_core_KE_CipherKey0_186_), .Y(n7176) );
  INVX1 U26973 ( .A(top_core_KE_CipherKey0_185_), .Y(n7175) );
  INVX1 U26974 ( .A(top_core_KE_CipherKey0_184_), .Y(n7174) );
  INVX1 U26975 ( .A(top_core_KE_CipherKey0_183_), .Y(n7173) );
  INVX1 U26976 ( .A(top_core_KE_CipherKey0_182_), .Y(n7172) );
  INVX1 U26977 ( .A(top_core_KE_CipherKey0_181_), .Y(n7171) );
  INVX1 U26978 ( .A(top_core_KE_CipherKey0_180_), .Y(n7170) );
  INVX1 U26979 ( .A(top_core_KE_CipherKey0_179_), .Y(n7169) );
  INVX1 U26980 ( .A(top_core_KE_CipherKey0_178_), .Y(n7168) );
  INVX1 U26981 ( .A(top_core_KE_CipherKey0_177_), .Y(n7167) );
  INVX1 U26982 ( .A(top_core_KE_CipherKey0_176_), .Y(n7166) );
  INVX1 U26983 ( .A(top_core_KE_CipherKey0_175_), .Y(n7165) );
  INVX1 U26984 ( .A(top_core_KE_CipherKey0_174_), .Y(n7164) );
  INVX1 U26985 ( .A(top_core_KE_CipherKey0_173_), .Y(n7163) );
  INVX1 U26986 ( .A(top_core_KE_CipherKey0_172_), .Y(n7162) );
  INVX1 U26987 ( .A(top_core_KE_CipherKey0_171_), .Y(n7161) );
  INVX1 U26988 ( .A(top_core_KE_CipherKey0_170_), .Y(n7160) );
  INVX1 U26989 ( .A(top_core_KE_CipherKey0_169_), .Y(n7159) );
  INVX1 U26990 ( .A(top_core_KE_CipherKey0_168_), .Y(n7158) );
  INVX1 U26991 ( .A(top_core_KE_CipherKey0_167_), .Y(n7157) );
  INVX1 U26992 ( .A(top_core_KE_CipherKey0_166_), .Y(n7156) );
  INVX1 U26993 ( .A(top_core_KE_CipherKey0_165_), .Y(n7155) );
  INVX1 U26994 ( .A(top_core_KE_CipherKey0_164_), .Y(n7154) );
  INVX1 U26995 ( .A(top_core_KE_CipherKey0_163_), .Y(n7153) );
  INVX1 U26996 ( .A(top_core_KE_CipherKey0_162_), .Y(n7152) );
  INVX1 U26997 ( .A(top_core_KE_CipherKey0_161_), .Y(n7151) );
  INVX1 U26998 ( .A(top_core_KE_CipherKey0_160_), .Y(n7150) );
  INVX1 U26999 ( .A(top_core_KE_CipherKey0_159_), .Y(n7149) );
  INVX1 U27000 ( .A(top_core_KE_CipherKey0_158_), .Y(n7148) );
  INVX1 U27001 ( .A(top_core_KE_CipherKey0_157_), .Y(n7147) );
  INVX1 U27002 ( .A(top_core_KE_CipherKey0_156_), .Y(n7146) );
  INVX1 U27003 ( .A(top_core_KE_CipherKey0_155_), .Y(n7145) );
  INVX1 U27004 ( .A(top_core_KE_CipherKey0_154_), .Y(n7144) );
  INVX1 U27005 ( .A(top_core_KE_CipherKey0_153_), .Y(n7143) );
  INVX1 U27006 ( .A(top_core_KE_CipherKey0_152_), .Y(n7142) );
  INVX1 U27007 ( .A(top_core_KE_CipherKey0_151_), .Y(n7141) );
  INVX1 U27008 ( .A(top_core_KE_CipherKey0_150_), .Y(n7140) );
  INVX1 U27009 ( .A(top_core_KE_CipherKey0_149_), .Y(n7139) );
  INVX1 U27010 ( .A(top_core_KE_CipherKey0_148_), .Y(n7138) );
  INVX1 U27011 ( .A(top_core_KE_CipherKey0_147_), .Y(n7137) );
  INVX1 U27012 ( .A(top_core_KE_CipherKey0_146_), .Y(n7136) );
  INVX1 U27013 ( .A(top_core_KE_CipherKey0_145_), .Y(n7135) );
  INVX1 U27014 ( .A(top_core_KE_CipherKey0_144_), .Y(n7134) );
  INVX1 U27015 ( .A(top_core_KE_CipherKey0_143_), .Y(n7133) );
  INVX1 U27016 ( .A(top_core_KE_CipherKey0_142_), .Y(n7132) );
  INVX1 U27017 ( .A(top_core_KE_CipherKey0_141_), .Y(n7131) );
  INVX1 U27018 ( .A(top_core_KE_CipherKey0_140_), .Y(n7130) );
  INVX1 U27019 ( .A(top_core_KE_CipherKey0_139_), .Y(n7129) );
  INVX1 U27020 ( .A(top_core_KE_CipherKey0_138_), .Y(n7128) );
  INVX1 U27021 ( .A(top_core_KE_CipherKey0_137_), .Y(n7127) );
  INVX1 U27022 ( .A(top_core_KE_CipherKey0_136_), .Y(n7126) );
  INVX1 U27023 ( .A(top_core_KE_CipherKey0_135_), .Y(n7125) );
  INVX1 U27024 ( .A(top_core_KE_CipherKey0_134_), .Y(n7124) );
  INVX1 U27025 ( .A(top_core_KE_CipherKey0_133_), .Y(n7123) );
  INVX1 U27026 ( .A(top_core_KE_CipherKey0_132_), .Y(n7122) );
  INVX1 U27027 ( .A(top_core_KE_CipherKey0_131_), .Y(n7121) );
  INVX1 U27028 ( .A(top_core_KE_CipherKey0_130_), .Y(n7120) );
  INVX1 U27029 ( .A(top_core_KE_CipherKey0_129_), .Y(n7119) );
  INVX1 U27030 ( .A(top_core_KE_CipherKey0_128_), .Y(n7118) );
  INVX1 U27031 ( .A(top_core_KE_CipherKey0_62_), .Y(n7086) );
  INVX1 U27032 ( .A(top_core_KE_CipherKey0_61_), .Y(n7085) );
  INVX1 U27033 ( .A(top_core_KE_CipherKey0_60_), .Y(n7084) );
  INVX1 U27034 ( .A(top_core_KE_CipherKey0_59_), .Y(n7083) );
  INVX1 U27035 ( .A(top_core_KE_CipherKey0_58_), .Y(n7082) );
  INVX1 U27036 ( .A(top_core_KE_CipherKey0_57_), .Y(n7081) );
  INVX1 U27037 ( .A(top_core_KE_CipherKey0_56_), .Y(n7080) );
  INVX1 U27038 ( .A(top_core_KE_CipherKey0_55_), .Y(n7079) );
  INVX1 U27039 ( .A(top_core_KE_CipherKey0_54_), .Y(n7078) );
  INVX1 U27040 ( .A(top_core_KE_CipherKey0_53_), .Y(n7077) );
  INVX1 U27041 ( .A(top_core_KE_CipherKey0_52_), .Y(n7076) );
  INVX1 U27042 ( .A(top_core_KE_CipherKey0_51_), .Y(n7075) );
  INVX1 U27043 ( .A(top_core_KE_CipherKey0_50_), .Y(n7074) );
  INVX1 U27044 ( .A(top_core_KE_CipherKey0_49_), .Y(n7073) );
  INVX1 U27045 ( .A(top_core_KE_CipherKey0_48_), .Y(n7072) );
  INVX1 U27046 ( .A(top_core_KE_CipherKey0_47_), .Y(n7071) );
  INVX1 U27047 ( .A(top_core_KE_CipherKey0_46_), .Y(n7070) );
  INVX1 U27048 ( .A(top_core_KE_CipherKey0_45_), .Y(n7069) );
  INVX1 U27049 ( .A(top_core_KE_CipherKey0_44_), .Y(n7068) );
  INVX1 U27050 ( .A(top_core_KE_CipherKey0_43_), .Y(n7067) );
  INVX1 U27051 ( .A(top_core_KE_CipherKey0_42_), .Y(n7066) );
  INVX1 U27052 ( .A(top_core_KE_CipherKey0_41_), .Y(n7065) );
  INVX1 U27053 ( .A(top_core_KE_CipherKey0_40_), .Y(n7064) );
  INVX1 U27054 ( .A(top_core_KE_CipherKey0_39_), .Y(n7063) );
  INVX1 U27055 ( .A(top_core_KE_CipherKey0_38_), .Y(n7062) );
  INVX1 U27056 ( .A(top_core_KE_CipherKey0_37_), .Y(n7061) );
  INVX1 U27057 ( .A(top_core_KE_CipherKey0_36_), .Y(n7060) );
  INVX1 U27058 ( .A(top_core_KE_CipherKey0_35_), .Y(n7059) );
  INVX1 U27059 ( .A(top_core_KE_CipherKey0_34_), .Y(n7058) );
  INVX1 U27060 ( .A(top_core_KE_CipherKey0_33_), .Y(n7057) );
  INVX1 U27061 ( .A(top_core_KE_CipherKey0_32_), .Y(n7056) );
  INVX1 U27062 ( .A(top_core_KE_CipherKey0_31_), .Y(n7055) );
  INVX1 U27063 ( .A(top_core_KE_CipherKey0_30_), .Y(n7054) );
  INVX1 U27064 ( .A(top_core_KE_CipherKey0_29_), .Y(n7053) );
  INVX1 U27065 ( .A(top_core_KE_CipherKey0_28_), .Y(n7052) );
  INVX1 U27066 ( .A(top_core_KE_CipherKey0_27_), .Y(n7051) );
  INVX1 U27067 ( .A(top_core_KE_CipherKey0_26_), .Y(n7050) );
  INVX1 U27068 ( .A(top_core_KE_CipherKey0_25_), .Y(n7049) );
  INVX1 U27069 ( .A(top_core_KE_CipherKey0_24_), .Y(n7048) );
  INVX1 U27070 ( .A(top_core_KE_CipherKey0_23_), .Y(n7047) );
  INVX1 U27071 ( .A(top_core_KE_CipherKey0_22_), .Y(n7046) );
  INVX1 U27072 ( .A(top_core_KE_CipherKey0_21_), .Y(n7045) );
  INVX1 U27073 ( .A(top_core_KE_CipherKey0_20_), .Y(n7044) );
  INVX1 U27074 ( .A(top_core_KE_CipherKey0_19_), .Y(n7043) );
  INVX1 U27075 ( .A(top_core_KE_CipherKey0_18_), .Y(n7042) );
  INVX1 U27076 ( .A(top_core_KE_CipherKey0_17_), .Y(n7041) );
  INVX1 U27077 ( .A(top_core_KE_CipherKey0_16_), .Y(n7040) );
  INVX1 U27078 ( .A(top_core_KE_CipherKey0_15_), .Y(n7039) );
  INVX1 U27079 ( .A(top_core_KE_CipherKey0_14_), .Y(n7038) );
  INVX1 U27080 ( .A(top_core_KE_CipherKey0_13_), .Y(n7037) );
  INVX1 U27081 ( .A(top_core_KE_CipherKey0_12_), .Y(n7036) );
  INVX1 U27082 ( .A(top_core_KE_CipherKey0_11_), .Y(n7035) );
  INVX1 U27083 ( .A(top_core_KE_CipherKey0_10_), .Y(n7034) );
  INVX1 U27084 ( .A(top_core_KE_CipherKey0_9_), .Y(n7033) );
  INVX1 U27085 ( .A(top_core_KE_CipherKey0_8_), .Y(n7032) );
  INVX1 U27086 ( .A(top_core_KE_CipherKey0_7_), .Y(n7031) );
  INVX1 U27087 ( .A(top_core_KE_CipherKey0_6_), .Y(n7030) );
  INVX1 U27088 ( .A(top_core_KE_CipherKey0_5_), .Y(n7029) );
  INVX1 U27089 ( .A(top_core_KE_CipherKey0_4_), .Y(n7028) );
  INVX1 U27090 ( .A(top_core_KE_CipherKey0_3_), .Y(n7027) );
  INVX1 U27091 ( .A(top_core_KE_CipherKey0_2_), .Y(n7026) );
  INVX1 U27092 ( .A(top_core_KE_CipherKey0_1_), .Y(n7025) );
  INVX1 U27093 ( .A(top_core_KE_CipherKey0_0_), .Y(n7024) );
  INVX1 U27094 ( .A(top_core_KE_CipherKey0_255_), .Y(n7245) );
  INVX1 U27095 ( .A(top_core_KE_CipherKey0_254_), .Y(n7244) );
  INVX1 U27096 ( .A(top_core_KE_CipherKey0_253_), .Y(n7243) );
  INVX1 U27097 ( .A(top_core_KE_CipherKey0_252_), .Y(n7242) );
  INVX1 U27098 ( .A(top_core_KE_CipherKey0_251_), .Y(n7241) );
  INVX1 U27099 ( .A(top_core_KE_CipherKey0_250_), .Y(n7240) );
  INVX1 U27100 ( .A(top_core_KE_CipherKey0_249_), .Y(n7239) );
  INVX1 U27101 ( .A(top_core_KE_CipherKey0_248_), .Y(n7238) );
  INVX1 U27102 ( .A(top_core_KE_CipherKey0_247_), .Y(n7237) );
  INVX1 U27103 ( .A(top_core_KE_CipherKey0_246_), .Y(n7236) );
  INVX1 U27104 ( .A(top_core_KE_CipherKey0_245_), .Y(n7235) );
  INVX1 U27105 ( .A(top_core_KE_CipherKey0_244_), .Y(n7234) );
  INVX1 U27106 ( .A(top_core_KE_CipherKey0_243_), .Y(n7233) );
  INVX1 U27107 ( .A(top_core_KE_CipherKey0_242_), .Y(n7232) );
  INVX1 U27108 ( .A(top_core_KE_CipherKey0_241_), .Y(n7231) );
  INVX1 U27109 ( .A(top_core_KE_CipherKey0_240_), .Y(n7230) );
  INVX1 U27110 ( .A(top_core_KE_CipherKey0_239_), .Y(n7229) );
  INVX1 U27111 ( .A(top_core_KE_CipherKey0_238_), .Y(n7228) );
  INVX1 U27112 ( .A(top_core_KE_CipherKey0_237_), .Y(n7227) );
  INVX1 U27113 ( .A(top_core_KE_CipherKey0_236_), .Y(n7226) );
  INVX1 U27114 ( .A(top_core_KE_CipherKey0_235_), .Y(n7225) );
  INVX1 U27115 ( .A(top_core_KE_CipherKey0_234_), .Y(n7224) );
  INVX1 U27116 ( .A(top_core_KE_CipherKey0_233_), .Y(n7223) );
  INVX1 U27117 ( .A(top_core_KE_CipherKey0_232_), .Y(n7222) );
  INVX1 U27118 ( .A(top_core_KE_CipherKey0_231_), .Y(n7221) );
  INVX1 U27119 ( .A(top_core_KE_CipherKey0_230_), .Y(n7220) );
  INVX1 U27120 ( .A(top_core_KE_CipherKey0_229_), .Y(n7219) );
  INVX1 U27121 ( .A(top_core_KE_CipherKey0_228_), .Y(n7218) );
  INVX1 U27122 ( .A(top_core_KE_CipherKey0_227_), .Y(n7217) );
  INVX1 U27123 ( .A(top_core_KE_CipherKey0_226_), .Y(n7216) );
  INVX1 U27124 ( .A(top_core_KE_CipherKey0_225_), .Y(n7215) );
  INVX1 U27125 ( .A(top_core_KE_CipherKey0_224_), .Y(n7214) );
  INVX1 U27126 ( .A(top_core_KE_CipherKey0_223_), .Y(n7213) );
  INVX1 U27127 ( .A(top_core_KE_CipherKey0_222_), .Y(n7212) );
  INVX1 U27128 ( .A(top_core_KE_CipherKey0_221_), .Y(n7211) );
  INVX1 U27129 ( .A(top_core_KE_CipherKey0_220_), .Y(n7210) );
  INVX1 U27130 ( .A(top_core_KE_CipherKey0_219_), .Y(n7209) );
  INVX1 U27131 ( .A(top_core_KE_CipherKey0_218_), .Y(n7208) );
  INVX1 U27132 ( .A(top_core_KE_CipherKey0_217_), .Y(n7207) );
  INVX1 U27133 ( .A(top_core_KE_CipherKey0_216_), .Y(n7206) );
  INVX1 U27134 ( .A(top_core_KE_CipherKey0_215_), .Y(n7205) );
  INVX1 U27135 ( .A(top_core_KE_CipherKey0_214_), .Y(n7204) );
  INVX1 U27136 ( .A(top_core_KE_CipherKey0_213_), .Y(n7203) );
  INVX1 U27137 ( .A(top_core_KE_CipherKey0_212_), .Y(n7202) );
  INVX1 U27138 ( .A(top_core_KE_CipherKey0_211_), .Y(n7201) );
  INVX1 U27139 ( .A(top_core_KE_CipherKey0_210_), .Y(n7200) );
  INVX1 U27140 ( .A(top_core_KE_CipherKey0_209_), .Y(n7199) );
  INVX1 U27141 ( .A(top_core_KE_CipherKey0_208_), .Y(n7198) );
  INVX1 U27142 ( .A(top_core_KE_CipherKey0_207_), .Y(n7197) );
  INVX1 U27143 ( .A(top_core_KE_CipherKey0_206_), .Y(n7196) );
  INVX1 U27144 ( .A(top_core_KE_CipherKey0_205_), .Y(n7195) );
  INVX1 U27145 ( .A(top_core_KE_CipherKey0_204_), .Y(n7194) );
  INVX1 U27146 ( .A(top_core_KE_CipherKey0_203_), .Y(n7193) );
  INVX1 U27147 ( .A(top_core_KE_CipherKey0_202_), .Y(n7192) );
  INVX1 U27148 ( .A(top_core_KE_CipherKey0_201_), .Y(n7191) );
  INVX1 U27149 ( .A(top_core_KE_CipherKey0_200_), .Y(n7190) );
  INVX1 U27150 ( .A(top_core_KE_CipherKey0_199_), .Y(n7189) );
  INVX1 U27151 ( .A(top_core_KE_CipherKey0_198_), .Y(n7188) );
  INVX1 U27152 ( .A(top_core_KE_CipherKey0_197_), .Y(n7187) );
  INVX1 U27153 ( .A(top_core_KE_CipherKey0_196_), .Y(n7186) );
  INVX1 U27154 ( .A(top_core_KE_CipherKey0_195_), .Y(n7185) );
  INVX1 U27155 ( .A(top_core_KE_CipherKey0_194_), .Y(n7184) );
  INVX1 U27156 ( .A(top_core_KE_CipherKey0_193_), .Y(n7183) );
  INVX1 U27157 ( .A(top_core_KE_CipherKey0_192_), .Y(n7182) );
  INVX1 U27158 ( .A(top_core_KE_prev_key1_reg_29_), .Y(n1759) );
  INVX1 U27159 ( .A(top_core_KE_prev_key1_reg_90_), .Y(n1650) );
  INVX1 U27160 ( .A(top_core_KE_prev_key1_reg_93_), .Y(n1642) );
  INVX1 U27161 ( .A(top_core_c_ready), .Y(n3644) );
  INVX1 U27162 ( .A(top_core_Addr[0]), .Y(n4034) );
  OR2X2 U27163 ( .A(n3541), .B(top_core_Core_Full), .Y(n896) );
  INVX1 U27164 ( .A(top_core_KE_prev_key1_reg_85_), .Y(n1665) );
  INVX1 U27165 ( .A(top_core_KE_prev_key1_reg_69_), .Y(n1723) );
  INVX1 U27166 ( .A(top_core_KE_prev_key1_reg_77_), .Y(n1694) );
  INVX1 U27167 ( .A(top_core_EC_operation), .Y(n2366) );
  DFFSRX2 top_core_io_inter_ok_reg ( .D(top_core_io_n1183), .CK(n_CLK), .SN(
        1'b1), .RN(n_RSTB), .Q(top_core_io_inter_ok), .QN(n4257) );
  XOR2XL U2 ( .A(n3989), .B(n7246), .Y(top_core_EC_n863) );
  OR2X1 U3 ( .A(n7246), .B(top_core_EC_rounds_2_), .Y(n7247) );
  OAI2BB2X1 U16777 ( .B0(n4195), .B1(n2), .A0N(n2), .A1N(n7246), .Y(
        top_core_EC_n1296) );
  OAI2BB1XL U18929 ( .A0N(n7246), .A1N(top_core_EC_rounds_2_), .B0(n7247), .Y(
        top_core_EC_N575) );
  NAND4BBX1 U18983 ( .AN(n18879), .BN(n4035), .C(top_core_EC_n1033), .D(
        top_core_EC_n1034), .Y(top_core_EC_n944) );
  XOR2X1 U23793 ( .A(top_core_EC_rounds_3_), .B(n3963), .Y(n18879) );
  PIW gen_data_pin_0__PDIN ( .PAD(DIN[0]), .C(n_DIN[0]) );
  PO16W gen_data_pin_0__PDOUT ( .I(n_DOUT[0]), .PAD(DOUT[0]) );
  PIW gen_data_pin_1__PDIN ( .PAD(DIN[1]), .C(n_DIN[1]) );
  PO16W gen_data_pin_1__PDOUT ( .I(n_DOUT[1]), .PAD(DOUT[1]) );
  PIW gen_data_pin_2__PDIN ( .PAD(DIN[2]), .C(n_DIN[2]) );
  PO16W gen_data_pin_2__PDOUT ( .I(n_DOUT[2]), .PAD(DOUT[2]) );
  PIW gen_data_pin_3__PDIN ( .PAD(DIN[3]), .C(n_DIN[3]) );
  PO16W gen_data_pin_3__PDOUT ( .I(n_DOUT[3]), .PAD(DOUT[3]) );
  PIW gen_data_pin_4__PDIN ( .PAD(DIN[4]), .C(n_DIN[4]) );
  PO16W gen_data_pin_4__PDOUT ( .I(n_DOUT[4]), .PAD(DOUT[4]) );
  PIW gen_data_pin_5__PDIN ( .PAD(DIN[5]), .C(n_DIN[5]) );
  PO16W gen_data_pin_5__PDOUT ( .I(n_DOUT[5]), .PAD(DOUT[5]) );
  PIW gen_data_pin_6__PDIN ( .PAD(DIN[6]), .C(n_DIN[6]) );
  PO16W gen_data_pin_6__PDOUT ( .I(n_DOUT[6]), .PAD(DOUT[6]) );
  PIW gen_data_pin_7__PDIN ( .PAD(DIN[7]), .C(n_DIN[7]) );
  PO16W gen_data_pin_7__PDOUT ( .I(n_DOUT[7]), .PAD(DOUT[7]) );
  PIW gen_addr_pin_0__PDIN ( .PAD(ADDR[0]), .C(n_ADDR[0]) );
  PIW gen_addr_pin_1__PDIN ( .PAD(ADDR[1]), .C(n_ADDR[1]) );
  PIW gen_addr_pin_2__PDIN ( .PAD(ADDR[2]), .C(n_ADDR[2]) );
  PIW gen_addr_pin_3__PDIN ( .PAD(ADDR[3]), .C(n_ADDR[3]) );
  PIW gen_addr_pin_4__PDIN ( .PAD(ADDR[4]), .C(n_ADDR[4]) );
  PIW gen_addr_pin_5__PDIN ( .PAD(ADDR[5]), .C(n_ADDR[5]) );
  PIW gen_addr_pin_6__PDIN ( .PAD(ADDR[6]), .C(n_ADDR[6]) );
endmodule

