module aes_tbox_r(a,d);
input	[7:0]	a;
output	[23:0]	d;
reg	[23:0]	d;

always @(a)
	case(a)
  8'h00: d = 24'b111101101010010001010010;
  8'h01: d = 24'b000110110001001000001001;
  8'h02: d = 24'b101111101101010001101010;
  8'h03: d = 24'b011001001011000111010101;
  8'h04: d = 24'b010100000110000000110000;
  8'h05: d = 24'b010110100110110000110110;
  8'h06: d = 24'b111101000101000110100101;
  8'h07: d = 24'b010010000111000000111000;
  8'h08: d = 24'b110110100110010110111111;
  8'h09: d = 24'b110000001000000001000000;
  8'h0a: d = 24'b111111100101110110100011;
  8'h0b: d = 24'b101110010010011110011110;
  8'h0c: d = 24'b100110000001100110000001;
  8'h0d: d = 24'b000011101111110111110011;
  8'h0e: d = 24'b011000101011010111010111;
  8'h0f: d = 24'b000101101110110111111011;
  8'h10: d = 24'b100001001111100001111100;
  8'h11: d = 24'b001111101101110111100011;
  8'h12: d = 24'b010010110111001000111001;
  8'h13: d = 24'b100111010001111110000010;
  8'h14: d = 24'b101101100010110110011011;
  8'h15: d = 24'b011100010101111000101111;
  8'h16: d = 24'b000110101110010111111111;
  8'h17: d = 24'b100100100001010110000111;
  8'h18: d = 24'b010111000110100000110100;
  8'h19: d = 24'b100010010000011110001110;
  8'h1a: d = 24'b110001011000011001000011;
  8'h1b: d = 24'b110011001000100001000100;
  8'h1c: d = 24'b010101111001001111000100;
  8'h1d: d = 24'b011110011010011111011110;
  8'h1e: d = 24'b001000001100100111101001;
  8'h1f: d = 24'b010001101000110111001011;
  8'h20: d = 24'b111111001010100001010100;
  8'h21: d = 24'b100011011111011001111011;
  8'h22: d = 24'b101001110011001110010100;
  8'h23: d = 24'b010101100110010000110010;
  8'h24: d = 24'b111100010101011110100110;
  8'h25: d = 24'b010111011001111111000010;
  8'h26: d = 24'b011001010100011000100011;
  8'h27: d = 24'b010001110111101000111101;
  8'h28: d = 24'b001010011100011111101110;
  8'h29: d = 24'b110101001001100001001100;
  8'h2a: d = 24'b101001000011000110010101;
  8'h2b: d = 24'b000111010001011000001011;
  8'h2c: d = 24'b110001101000010001000010;
  8'h2d: d = 24'b000101011110111111111010;
  8'h2e: d = 24'b010111101001110111000011;
  8'h2f: d = 24'b110100101001110001001110;
  8'h30: d = 24'b000110000001000000001000;
  8'h31: d = 24'b011100100101110000101110;
  8'h32: d = 24'b111110000101100110100001;
  8'h33: d = 24'b101010101100110001100110;
  8'h34: d = 24'b011110000101000000101000;
  8'h35: d = 24'b011100001010100111011001;
  8'h36: d = 24'b011011000100100000100100;
  8'h37: d = 24'b110011010111111110110010;
  8'h38: d = 24'b100110101110110001110110;
  8'h39: d = 24'b111011011011011001011011;
  8'h3a: d = 24'b111111010101111110100010;
  8'h3b: d = 24'b110110111001001001001001;
  8'h3c: d = 24'b101101111101101001101101;
  8'h3d: d = 24'b100001100000110110001011;
  8'h3e: d = 24'b011010001011100111010001;
  8'h3f: d = 24'b011011110100101000100101;
  8'h40: d = 24'b100101101110010001110010;
  8'h41: d = 24'b000100111110101111111000;
  8'h42: d = 24'b000000011111011111110110;
  8'h43: d = 24'b101011001100100001100100;
  8'h44: d = 24'b100100010001011110000110;
  8'h45: d = 24'b101110001101000001101000;
  8'h46: d = 24'b101100110010101110011000;
  8'h47: d = 24'b001110100010110000010110;
  8'h48: d = 24'b011001111011001111010100;
  8'h49: d = 24'b111101110101001110100100;
  8'h4a: d = 24'b111001001011100001011100;
  8'h4b: d = 24'b010011111000001111001100;
  8'h4c: d = 24'b111001111011101001011101;
  8'h4d: d = 24'b101011111100101001100101;
  8'h4e: d = 24'b110000010111011110110110;
  8'h4f: d = 24'b101011010011111110010010;
  8'h50: d = 24'b101101001101100001101100;
  8'h51: d = 24'b100100001110000001110000;
  8'h52: d = 24'b110110001001000001001000;
  8'h53: d = 24'b111100001010000001010000;
  8'h54: d = 24'b000111001110000111111101;
  8'h55: d = 24'b001011001100000111101101;
  8'h56: d = 24'b110100000110100110111001;
  8'h57: d = 24'b011101011010111111011010;
  8'h58: d = 24'b111000101011110001011110;
  8'h59: d = 24'b001111110010101000010101;
  8'h5a: d = 24'b110010101000110001000110;
  8'h5b: d = 24'b111110011010111001010111;
  8'h5c: d = 24'b111100100101010110100111;
  8'h5d: d = 24'b100011000000000110001101;
  8'h5e: d = 24'b101111000010000110011101;
  8'h5f: d = 24'b100101110001001110000100;
  8'h60: d = 24'b101010110011101110010000;
  8'h61: d = 24'b011100111010101111011000;
  8'h62: d = 24'b111001100100110110101011;
  8'h63: d = 24'b000000000000000000000000;
  8'h64: d = 24'b100011110000001110001100;
  8'h65: d = 24'b110111110110001110111100;
  8'h66: d = 24'b011011101011110111010011;
  8'h67: d = 24'b000111100001010000001010;
  8'h68: d = 24'b000000101111010111110111;
  8'h69: d = 24'b001101111101001111100100;
  8'h6a: d = 24'b111010001011000001011000;
  8'h6b: d = 24'b000011110000101000000101;
  8'h6c: d = 24'b110100110110101110111000;
  8'h6d: d = 24'b110011100111110110110011;
  8'h6e: d = 24'b110011111000101001000101;
  8'h6f: d = 24'b000010100000110000000110;
  8'h70: d = 24'b011010111011101111010000;
  8'h71: d = 24'b011101000101100000101100;
  8'h72: d = 24'b001000100011110000011110;
  8'h73: d = 24'b100010100000010110001111;
  8'h74: d = 24'b010001011000111111001010;
  8'h75: d = 24'b010000010111111000111111;
  8'h76: d = 24'b000100010001111000001111;
  8'h77: d = 24'b000001100000010000000010;
  8'h78: d = 24'b010110001001100111000001;
  8'h79: d = 24'b111010100100010110101111;
  8'h7a: d = 24'b110111000110000110111101;
  8'h7b: d = 24'b000001010000011000000011;
  8'h7c: d = 24'b000000110000001000000001;
  8'h7d: d = 24'b001101010010011000010011;
  8'h7e: d = 24'b100001010000111110001010;
  8'h7f: d = 24'b101111011101011001101011;
  8'h80: d = 24'b010011100111010000111010;
  8'h81: d = 24'b101010000011100110010001;
  8'h82: d = 24'b001100110010001000010001;
  8'h83: d = 24'b110000111000001001000001;
  8'h84: d = 24'b110100011001111001001111;
  8'h85: d = 24'b101010011100111001100111;
  8'h86: d = 24'b011111111010001111011100;
  8'h87: d = 24'b001001011100111111101010;
  8'h88: d = 24'b101000100011010110010111;
  8'h89: d = 24'b000011011111111111110010;
  8'h8a: d = 24'b010010101000010111001111;
  8'h8b: d = 24'b010010011000011111001110;
  8'h8c: d = 24'b000010111111101111110000;
  8'h8d: d = 24'b110001110111001110110100;
  8'h8e: d = 24'b001100011101011111100110;
  8'h8f: d = 24'b100101011110011001110011;
  8'h90: d = 24'b101000010011011110010110;
  8'h91: d = 24'b111011110100001110101100;
  8'h92: d = 24'b100111001110100001110100;
  8'h93: d = 24'b011001100100010000100010;
  8'h94: d = 24'b001100101101010111100111;
  8'h95: d = 24'b111011000100000110101101;
  8'h96: d = 24'b010111110110101000110101;
  8'h97: d = 24'b100101000001000110000101;
  8'h98: d = 24'b001111011101111111100010;
  8'h99: d = 24'b000100001110100111111001;
  8'h9a: d = 24'b010110010110111000110111;
  8'h9b: d = 24'b001000111100101111101000;
  8'h9c: d = 24'b001001000011100000011100;
  8'h9d: d = 24'b100111111110101001110101;
  8'h9e: d = 24'b011110101010010111011111;
  8'h9f: d = 24'b101100101101110001101110;
  8'ha0: d = 24'b110010011000111001000111;
  8'ha1: d = 24'b000010001111100111110001;
  8'ha2: d = 24'b001011100011010000011010;
  8'ha3: d = 24'b100100111110001001110001;
  8'ha4: d = 24'b001001110011101000011101;
  8'ha5: d = 24'b011110110101001000101001;
  8'ha6: d = 24'b010101001001000111000101;
  8'ha7: d = 24'b100000000000100110001001;
  8'ha8: d = 24'b101100011101111001101111;
  8'ha9: d = 24'b110000100111010110110111;
  8'haa: d = 24'b101001101100010001100010;
  8'hab: d = 24'b000100100001110000001110;
  8'hac: d = 24'b111001010100111110101010;
  8'had: d = 24'b001010000011000000011000;
  8'hae: d = 24'b110110010110011110111110;
  8'haf: d = 24'b001011010011011000011011;
  8'hb0: d = 24'b000111111110001111111100;
  8'hb1: d = 24'b111110101010110001010110;
  8'hb2: d = 24'b010000100111110000111110;
  8'hb3: d = 24'b110111011001011001001011;
  8'hb4: d = 24'b010100011001011111000110;
  8'hb5: d = 24'b011011011011111111010010;
  8'hb6: d = 24'b100010111111001001111001;
  8'hb7: d = 24'b011000000100000000100000;
  8'hb8: d = 24'b101101010010111110011010;
  8'hb9: d = 24'b011101101010110111011011;
  8'hba: d = 24'b010110111001101111000000;
  8'hbb: d = 24'b000110011110011111111110;
  8'hbc: d = 24'b100010001111000001111000;
  8'hbd: d = 24'b010011001000000111001101;
  8'hbe: d = 24'b111011101011010001011010;
  8'hbf: d = 24'b000001111111001111110100;
  8'hc0: d = 24'b001000010011111000011111;
  8'hc1: d = 24'b011111001010000111011101;
  8'hc2: d = 24'b111000110100101110101000;
  8'hc3: d = 24'b010101010110011000110011;
  8'hc4: d = 24'b100000110000101110001000;
  8'hc5: d = 24'b000010010000111000000111;
  8'hc6: d = 24'b010100101001010111000111;
  8'hc7: d = 24'b010100110110001000110001;
  8'hc8: d = 24'b110010000111100110110001;
  8'hc9: d = 24'b001101100010010000010010;
  8'hca: d = 24'b001100000010000000010000;
  8'hcb: d = 24'b111010111011001001011001;
  8'hcc: d = 24'b011010010100111000100111;
  8'hcd: d = 24'b100110110001101110000000;
  8'hce: d = 24'b001011111100001111101100;
  8'hcf: d = 24'b111000011011111001011111;
  8'hd0: d = 24'b101000001100000001100000;
  8'hd1: d = 24'b111100111010001001010001;
  8'hd2: d = 24'b100000011111111001111111;
  8'hd3: d = 24'b111000000100100110101001;
  8'hd4: d = 24'b001010110011001000011001;
  8'hd5: d = 24'b110001000111000110110101;
  8'hd6: d = 24'b110111101001010001001010;
  8'hd7: d = 24'b000101110001101000001101;
  8'hd8: d = 24'b011101110101101000101101;
  8'hd9: d = 24'b001101001101000111100101;
  8'hda: d = 24'b100011101111010001111010;
  8'hdb: d = 24'b101110100010010110011111;
  8'hdc: d = 24'b101011100011110110010011;
  8'hdd: d = 24'b010000001000100111001001;
  8'hde: d = 24'b101111110010001110011100;
  8'hdf: d = 24'b001010101100010111101111;
  8'he0: d = 24'b111110110101101110100000;
  8'he1: d = 24'b001110111101101111100000;
  8'he2: d = 24'b010011010111011000111011;
  8'he3: d = 24'b110101111001101001001101;
  8'he4: d = 24'b111010010100011110101110;
  8'he5: d = 24'b011111100101010000101010;
  8'he6: d = 24'b000001001111000111110101;
  8'he7: d = 24'b110010110111101110110000;
  8'he8: d = 24'b010000111000101111001000;
  8'he9: d = 24'b001001101100110111101011;
  8'hea: d = 24'b110101100110110110111011;
  8'heb: d = 24'b010001000111100000111100;
  8'hec: d = 24'b100111100001110110000011;
  8'hed: d = 24'b111101011010011001010011;
  8'hee: d = 24'b101100000010100110011001;
  8'hef: d = 24'b101000111100001001100001;
  8'hf0: d = 24'b001110010010111000010111;
  8'hf1: d = 24'b011111010101011000101011;
  8'hf2: d = 24'b000011000000100000000100;
  8'hf3: d = 24'b100000101111110001111110;
  8'hf4: d = 24'b110101010110111110111010;
  8'hf5: d = 24'b100110011110111001110111;
  8'hf6: d = 24'b011000011011011111010110;
  8'hf7: d = 24'b011010100100110000100110;
  8'hf8: d = 24'b001110001101100111100001;
  8'hf9: d = 24'b101110111101001001101001;
  8'hfa: d = 24'b001111000010100000010100;
  8'hfb: d = 24'b101001011100011001100011;
  8'hfc: d = 24'b111111111010101001010101;
  8'hfd: d = 24'b011000110100001000100001;
  8'hfe: d = 24'b000101000001100000001100;
  8'hff: d = 24'b100001111111101001111101;
	endcase

endmodule
